/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 1 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 2 register stage(s) in total */

module CRAFT_GHPCLL_ANF_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [63:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [1023:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1152 ;
    wire signal_1154 ;
    wire signal_1156 ;
    wire signal_1158 ;
    wire signal_1160 ;
    wire signal_1162 ;
    wire signal_1164 ;
    wire signal_1166 ;
    wire signal_1168 ;
    wire signal_1170 ;
    wire signal_1172 ;
    wire signal_1174 ;
    wire signal_1176 ;
    wire signal_1178 ;
    wire signal_1180 ;
    wire signal_1182 ;
    wire signal_1184 ;
    wire signal_1186 ;
    wire signal_1188 ;
    wire signal_1190 ;
    wire signal_1192 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1198 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1204 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1210 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1216 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1222 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1234 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1246 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1252 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1258 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1264 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1270 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1277 ;
    wire signal_1280 ;
    wire signal_1283 ;
    wire signal_1286 ;
    wire signal_1289 ;
    wire signal_1292 ;
    wire signal_1295 ;
    wire signal_1298 ;
    wire signal_1301 ;
    wire signal_1304 ;
    wire signal_1307 ;
    wire signal_1310 ;
    wire signal_1313 ;
    wire signal_1316 ;
    wire signal_1319 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1445 ;
    wire signal_1448 ;
    wire signal_1451 ;
    wire signal_1454 ;
    wire signal_1457 ;
    wire signal_1460 ;
    wire signal_1463 ;
    wire signal_1466 ;
    wire signal_1469 ;
    wire signal_1472 ;
    wire signal_1475 ;
    wire signal_1478 ;
    wire signal_1481 ;
    wire signal_1484 ;
    wire signal_1487 ;
    wire signal_1490 ;
    wire signal_1493 ;
    wire signal_1496 ;
    wire signal_1499 ;
    wire signal_1502 ;
    wire signal_1505 ;
    wire signal_1508 ;
    wire signal_1511 ;
    wire signal_1514 ;
    wire signal_1517 ;
    wire signal_1520 ;
    wire signal_1523 ;
    wire signal_1526 ;
    wire signal_1529 ;
    wire signal_1532 ;
    wire signal_1535 ;
    wire signal_1538 ;
    wire signal_1541 ;
    wire signal_1544 ;
    wire signal_1547 ;
    wire signal_1550 ;
    wire signal_1553 ;
    wire signal_1556 ;
    wire signal_1559 ;
    wire signal_1562 ;
    wire signal_1565 ;
    wire signal_1568 ;
    wire signal_1571 ;
    wire signal_1574 ;
    wire signal_1577 ;
    wire signal_1580 ;
    wire signal_1583 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;

    /* cells in depth 0 */
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_177 ( .a ({signal_1532, signal_894}), .b ({1'b0, signal_266}), .c ({signal_1603, signal_333}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_180 ( .a ({signal_1535, signal_893}), .b ({1'b0, signal_1014}), .c ({signal_1605, signal_335}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_183 ( .a ({signal_1538, signal_892}), .b ({1'b0, signal_1013}), .c ({signal_1607, signal_337}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_186 ( .a ({signal_1541, signal_891}), .b ({1'b0, 1'b0}), .c ({signal_1609, signal_339}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_189 ( .a ({signal_1544, signal_890}), .b ({1'b0, signal_265}), .c ({signal_1611, signal_341}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_192 ( .a ({signal_1547, signal_889}), .b ({1'b0, signal_1011}), .c ({signal_1613, signal_343}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_195 ( .a ({signal_1550, signal_888}), .b ({1'b0, signal_1010}), .c ({signal_1615, signal_345}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_198 ( .a ({signal_1553, signal_887}), .b ({1'b0, signal_1009}), .c ({signal_1617, signal_347}) ) ;
    INV_X1 cell_712 ( .A (signal_1000), .ZN (signal_692) ) ;
    INV_X1 cell_713 ( .A (signal_692), .ZN (signal_693) ) ;
    INV_X1 cell_714 ( .A (signal_692), .ZN (signal_694) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_715 ( .s (signal_1000), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1277, signal_934}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_716 ( .s (signal_693), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1445, signal_933}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_717 ( .s (signal_1000), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1280, signal_932}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_718 ( .s (signal_693), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1448, signal_931}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_719 ( .s (signal_693), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1451, signal_930}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_720 ( .s (signal_693), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1454, signal_929}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_721 ( .s (signal_693), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1457, signal_928}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_722 ( .s (signal_693), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1460, signal_927}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_723 ( .s (signal_693), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1463, signal_926}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_724 ( .s (signal_693), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1466, signal_925}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_725 ( .s (signal_693), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1469, signal_924}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_726 ( .s (signal_693), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1472, signal_923}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_727 ( .s (signal_693), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1475, signal_922}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_728 ( .s (signal_693), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1478, signal_921}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_729 ( .s (signal_693), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1481, signal_920}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_730 ( .s (signal_693), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1484, signal_919}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_731 ( .s (signal_693), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1487, signal_918}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_732 ( .s (signal_693), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1490, signal_917}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_733 ( .s (signal_693), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1493, signal_916}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_734 ( .s (signal_693), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1496, signal_915}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_735 ( .s (signal_693), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1499, signal_914}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_736 ( .s (signal_693), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1502, signal_913}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_737 ( .s (signal_1000), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1283, signal_912}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_738 ( .s (signal_1000), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1286, signal_911}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_739 ( .s (signal_1000), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1289, signal_910}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_740 ( .s (signal_1000), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1292, signal_909}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_741 ( .s (signal_1000), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1295, signal_908}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_742 ( .s (signal_1000), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1298, signal_907}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_743 ( .s (signal_694), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1505, signal_906}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_744 ( .s (signal_694), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1508, signal_905}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_745 ( .s (signal_694), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1511, signal_904}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_746 ( .s (signal_694), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1514, signal_903}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_747 ( .s (signal_694), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1517, signal_902}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_748 ( .s (signal_1000), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1301, signal_901}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_749 ( .s (signal_694), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1520, signal_900}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_750 ( .s (signal_694), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1523, signal_899}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_751 ( .s (signal_1000), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1304, signal_898}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_752 ( .s (signal_694), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1526, signal_897}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_753 ( .s (signal_694), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1529, signal_896}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_754 ( .s (signal_1000), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1307, signal_895}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_755 ( .s (signal_694), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1532, signal_894}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_756 ( .s (signal_694), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1535, signal_893}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_757 ( .s (signal_694), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1538, signal_892}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_758 ( .s (signal_694), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1541, signal_891}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_759 ( .s (signal_694), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1544, signal_890}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_760 ( .s (signal_694), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1547, signal_889}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_761 ( .s (signal_694), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1550, signal_888}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_762 ( .s (signal_694), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1553, signal_887}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_763 ( .s (signal_694), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1556, signal_886}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_764 ( .s (signal_694), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1559, signal_885}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_765 ( .s (signal_694), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1562, signal_884}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_766 ( .s (signal_694), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1565, signal_883}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_767 ( .s (signal_694), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1568, signal_882}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_768 ( .s (signal_1000), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1310, signal_881}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_769 ( .s (signal_1000), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1313, signal_880}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_770 ( .s (signal_694), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1571, signal_879}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_771 ( .s (signal_1000), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1316, signal_878}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_772 ( .s (signal_694), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1574, signal_877}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_773 ( .s (signal_694), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1577, signal_876}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_774 ( .s (signal_1000), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1319, signal_875}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_775 ( .s (signal_694), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1580, signal_874}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_776 ( .s (signal_694), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1583, signal_873}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_777 ( .s (signal_1000), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1322, signal_872}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_778 ( .s (signal_694), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1586, signal_871}) ) ;
    MUX2_X1 cell_779 ( .S (rst), .A (signal_1007), .B (1'b1), .Z (signal_266) ) ;
    MUX2_X1 cell_780 ( .S (rst), .A (signal_1006), .B (1'b0), .Z (signal_1014) ) ;
    MUX2_X1 cell_781 ( .S (rst), .A (signal_1005), .B (1'b0), .Z (signal_1013) ) ;
    MUX2_X1 cell_782 ( .S (rst), .A (signal_1004), .B (1'b1), .Z (signal_265) ) ;
    MUX2_X1 cell_783 ( .S (rst), .A (signal_1003), .B (1'b0), .Z (signal_1011) ) ;
    MUX2_X1 cell_784 ( .S (rst), .A (signal_1002), .B (1'b0), .Z (signal_1010) ) ;
    MUX2_X1 cell_785 ( .S (rst), .A (signal_1001), .B (1'b0), .Z (signal_1009) ) ;
    XOR2_X1 cell_786 ( .A (signal_265), .B (signal_1011), .Z (signal_1008) ) ;
    XOR2_X1 cell_787 ( .A (signal_1014), .B (signal_266), .Z (signal_1012) ) ;
    AND2_X1 cell_802 ( .A1 (signal_1009), .A2 (signal_702), .ZN (signal_267) ) ;
    NOR2_X1 cell_803 ( .A1 (signal_703), .A2 (signal_704), .ZN (signal_702) ) ;
    NAND2_X1 cell_804 ( .A1 (signal_705), .A2 (signal_706), .ZN (signal_704) ) ;
    NOR2_X1 cell_805 ( .A1 (signal_1011), .A2 (signal_1010), .ZN (signal_706) ) ;
    NOR2_X1 cell_806 ( .A1 (signal_1014), .A2 (signal_265), .ZN (signal_705) ) ;
    NAND2_X1 cell_807 ( .A1 (signal_266), .A2 (signal_1013), .ZN (signal_703) ) ;
    MUX2_X1 cell_808 ( .S (rst), .A (signal_1016), .B (1'b0), .Z (signal_1000) ) ;
    MUX2_X1 cell_809 ( .S (rst), .A (signal_1015), .B (1'b0), .Z (signal_999) ) ;
    XNOR2_X1 cell_810 ( .A (signal_707), .B (signal_999), .ZN (signal_1017) ) ;
    XNOR2_X1 cell_811 ( .A (signal_1000), .B (1'b0), .ZN (signal_707) ) ;
    INV_X1 cell_812 ( .A (signal_1000), .ZN (signal_1018) ) ;

    /* cells in depth 1 */
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_0 ( .s (signal_2707), .b ({signal_1146, signal_774}), .a ({signal_2709, signal_2708}), .c ({signal_1148, signal_870}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1 ( .s (signal_2707), .b ({signal_1145, signal_773}), .a ({signal_2711, signal_2710}), .c ({signal_1150, signal_869}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2 ( .s (signal_2707), .b ({signal_1144, signal_772}), .a ({signal_2713, signal_2712}), .c ({signal_1152, signal_868}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_3 ( .s (signal_2707), .b ({signal_1143, signal_771}), .a ({signal_2715, signal_2714}), .c ({signal_1154, signal_867}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_4 ( .s (signal_2707), .b ({signal_1142, signal_770}), .a ({signal_2717, signal_2716}), .c ({signal_1156, signal_866}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_5 ( .s (signal_2707), .b ({signal_1141, signal_769}), .a ({signal_2719, signal_2718}), .c ({signal_1158, signal_865}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_6 ( .s (signal_2707), .b ({signal_1140, signal_768}), .a ({signal_2721, signal_2720}), .c ({signal_1160, signal_864}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_7 ( .s (signal_2707), .b ({signal_1139, signal_767}), .a ({signal_2723, signal_2722}), .c ({signal_1162, signal_863}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_8 ( .s (signal_2707), .b ({signal_1138, signal_766}), .a ({signal_2725, signal_2724}), .c ({signal_1164, signal_862}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_9 ( .s (signal_2707), .b ({signal_1137, signal_765}), .a ({signal_2727, signal_2726}), .c ({signal_1166, signal_861}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_10 ( .s (signal_2707), .b ({signal_1136, signal_764}), .a ({signal_2729, signal_2728}), .c ({signal_1168, signal_860}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_11 ( .s (signal_2707), .b ({signal_1135, signal_763}), .a ({signal_2731, signal_2730}), .c ({signal_1170, signal_859}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_12 ( .s (signal_2707), .b ({signal_1134, signal_762}), .a ({signal_2733, signal_2732}), .c ({signal_1172, signal_858}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_13 ( .s (signal_2707), .b ({signal_1133, signal_761}), .a ({signal_2735, signal_2734}), .c ({signal_1174, signal_857}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_14 ( .s (signal_2707), .b ({signal_1132, signal_760}), .a ({signal_2737, signal_2736}), .c ({signal_1176, signal_856}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_15 ( .s (signal_2707), .b ({signal_1131, signal_759}), .a ({signal_2739, signal_2738}), .c ({signal_1178, signal_855}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_16 ( .s (signal_2707), .b ({signal_1130, signal_758}), .a ({signal_2741, signal_2740}), .c ({signal_1180, signal_854}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_17 ( .s (signal_2707), .b ({signal_1129, signal_757}), .a ({signal_2743, signal_2742}), .c ({signal_1182, signal_853}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_18 ( .s (signal_2707), .b ({signal_1128, signal_756}), .a ({signal_2745, signal_2744}), .c ({signal_1184, signal_852}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_19 ( .s (signal_2707), .b ({signal_1127, signal_755}), .a ({signal_2747, signal_2746}), .c ({signal_1186, signal_851}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_20 ( .s (signal_2707), .b ({signal_1126, signal_754}), .a ({signal_2749, signal_2748}), .c ({signal_1188, signal_850}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_21 ( .s (signal_2707), .b ({signal_1125, signal_753}), .a ({signal_2751, signal_2750}), .c ({signal_1190, signal_849}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_22 ( .s (signal_2707), .b ({signal_1124, signal_752}), .a ({signal_2753, signal_2752}), .c ({signal_1192, signal_848}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_23 ( .s (signal_2707), .b ({signal_1123, signal_751}), .a ({signal_2755, signal_2754}), .c ({signal_1194, signal_847}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_24 ( .s (signal_2707), .b ({signal_1122, signal_750}), .a ({signal_2757, signal_2756}), .c ({signal_1196, signal_846}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_25 ( .s (signal_2707), .b ({signal_1121, signal_749}), .a ({signal_2759, signal_2758}), .c ({signal_1198, signal_845}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_26 ( .s (signal_2707), .b ({signal_1120, signal_748}), .a ({signal_2761, signal_2760}), .c ({signal_1200, signal_844}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_27 ( .s (signal_2707), .b ({signal_1119, signal_747}), .a ({signal_2763, signal_2762}), .c ({signal_1202, signal_843}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_28 ( .s (signal_2707), .b ({signal_1118, signal_746}), .a ({signal_2765, signal_2764}), .c ({signal_1204, signal_842}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_29 ( .s (signal_2707), .b ({signal_1117, signal_745}), .a ({signal_2767, signal_2766}), .c ({signal_1206, signal_841}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_30 ( .s (signal_2707), .b ({signal_1116, signal_744}), .a ({signal_2769, signal_2768}), .c ({signal_1208, signal_840}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_31 ( .s (signal_2707), .b ({signal_1115, signal_743}), .a ({signal_2771, signal_2770}), .c ({signal_1210, signal_839}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_32 ( .s (signal_2707), .b ({signal_1114, signal_742}), .a ({signal_2773, signal_2772}), .c ({signal_1212, signal_806}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_33 ( .s (signal_2707), .b ({signal_1113, signal_741}), .a ({signal_2775, signal_2774}), .c ({signal_1214, signal_805}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_34 ( .s (signal_2707), .b ({signal_1112, signal_740}), .a ({signal_2777, signal_2776}), .c ({signal_1216, signal_804}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_35 ( .s (signal_2707), .b ({signal_1111, signal_739}), .a ({signal_2779, signal_2778}), .c ({signal_1218, signal_803}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_36 ( .s (signal_2707), .b ({signal_1110, signal_738}), .a ({signal_2781, signal_2780}), .c ({signal_1220, signal_802}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_37 ( .s (signal_2707), .b ({signal_1109, signal_737}), .a ({signal_2783, signal_2782}), .c ({signal_1222, signal_801}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_38 ( .s (signal_2707), .b ({signal_1108, signal_736}), .a ({signal_2785, signal_2784}), .c ({signal_1224, signal_800}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_39 ( .s (signal_2707), .b ({signal_1107, signal_735}), .a ({signal_2787, signal_2786}), .c ({signal_1226, signal_799}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_40 ( .s (signal_2707), .b ({signal_1106, signal_734}), .a ({signal_2789, signal_2788}), .c ({signal_1228, signal_798}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_41 ( .s (signal_2707), .b ({signal_1105, signal_733}), .a ({signal_2791, signal_2790}), .c ({signal_1230, signal_797}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_42 ( .s (signal_2707), .b ({signal_1104, signal_732}), .a ({signal_2793, signal_2792}), .c ({signal_1232, signal_796}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_43 ( .s (signal_2707), .b ({signal_1103, signal_731}), .a ({signal_2795, signal_2794}), .c ({signal_1234, signal_795}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_44 ( .s (signal_2707), .b ({signal_1102, signal_730}), .a ({signal_2797, signal_2796}), .c ({signal_1236, signal_794}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_45 ( .s (signal_2707), .b ({signal_1101, signal_729}), .a ({signal_2799, signal_2798}), .c ({signal_1238, signal_793}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_46 ( .s (signal_2707), .b ({signal_1100, signal_728}), .a ({signal_2801, signal_2800}), .c ({signal_1240, signal_792}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_47 ( .s (signal_2707), .b ({signal_1099, signal_727}), .a ({signal_2803, signal_2802}), .c ({signal_1242, signal_791}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_48 ( .s (signal_2707), .b ({signal_1098, signal_726}), .a ({signal_2805, signal_2804}), .c ({signal_1244, signal_790}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_49 ( .s (signal_2707), .b ({signal_1097, signal_725}), .a ({signal_2807, signal_2806}), .c ({signal_1246, signal_789}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_50 ( .s (signal_2707), .b ({signal_1096, signal_724}), .a ({signal_2809, signal_2808}), .c ({signal_1248, signal_788}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_51 ( .s (signal_2707), .b ({signal_1095, signal_723}), .a ({signal_2811, signal_2810}), .c ({signal_1250, signal_787}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_52 ( .s (signal_2707), .b ({signal_1094, signal_722}), .a ({signal_2813, signal_2812}), .c ({signal_1252, signal_786}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_53 ( .s (signal_2707), .b ({signal_1093, signal_721}), .a ({signal_2815, signal_2814}), .c ({signal_1254, signal_785}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_54 ( .s (signal_2707), .b ({signal_1092, signal_720}), .a ({signal_2817, signal_2816}), .c ({signal_1256, signal_784}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_55 ( .s (signal_2707), .b ({signal_1091, signal_719}), .a ({signal_2819, signal_2818}), .c ({signal_1258, signal_783}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_56 ( .s (signal_2707), .b ({signal_1090, signal_718}), .a ({signal_2821, signal_2820}), .c ({signal_1260, signal_782}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_57 ( .s (signal_2707), .b ({signal_1089, signal_717}), .a ({signal_2823, signal_2822}), .c ({signal_1262, signal_781}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_58 ( .s (signal_2707), .b ({signal_1088, signal_716}), .a ({signal_2825, signal_2824}), .c ({signal_1264, signal_780}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_59 ( .s (signal_2707), .b ({signal_1087, signal_715}), .a ({signal_2827, signal_2826}), .c ({signal_1266, signal_779}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_60 ( .s (signal_2707), .b ({signal_1086, signal_714}), .a ({signal_2829, signal_2828}), .c ({signal_1268, signal_778}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_61 ( .s (signal_2707), .b ({signal_1085, signal_713}), .a ({signal_2831, signal_2830}), .c ({signal_1270, signal_777}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_62 ( .s (signal_2707), .b ({signal_1084, signal_712}), .a ({signal_2833, signal_2832}), .c ({signal_1272, signal_776}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_63 ( .s (signal_2707), .b ({signal_1083, signal_711}), .a ({signal_2835, signal_2834}), .c ({signal_1274, signal_775}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_64 ( .a ({signal_1324, signal_268}), .b ({signal_1323, signal_269}), .c ({signal_1403, signal_822}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_65 ( .a ({signal_1180, signal_854}), .b ({signal_1148, signal_870}), .c ({signal_1323, signal_269}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_66 ( .a ({1'b0, 1'b0}), .b ({signal_1244, signal_790}), .c ({signal_1324, signal_268}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_67 ( .a ({signal_1325, signal_270}), .b ({signal_1148, signal_870}), .c ({signal_1404, signal_838}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_68 ( .a ({1'b0, 1'b0}), .b ({signal_1212, signal_806}), .c ({signal_1325, signal_270}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_69 ( .a ({signal_1327, signal_271}), .b ({signal_1326, signal_272}), .c ({signal_1405, signal_821}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_70 ( .a ({signal_1182, signal_853}), .b ({signal_1150, signal_869}), .c ({signal_1326, signal_272}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_71 ( .a ({1'b0, 1'b0}), .b ({signal_1246, signal_789}), .c ({signal_1327, signal_271}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_72 ( .a ({signal_1328, signal_273}), .b ({signal_1150, signal_869}), .c ({signal_1406, signal_837}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_73 ( .a ({1'b0, 1'b0}), .b ({signal_1214, signal_805}), .c ({signal_1328, signal_273}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_74 ( .a ({signal_1330, signal_274}), .b ({signal_1329, signal_275}), .c ({signal_1407, signal_820}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_75 ( .a ({signal_1184, signal_852}), .b ({signal_1152, signal_868}), .c ({signal_1329, signal_275}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_76 ( .a ({1'b0, 1'b0}), .b ({signal_1248, signal_788}), .c ({signal_1330, signal_274}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_77 ( .a ({signal_1331, signal_276}), .b ({signal_1152, signal_868}), .c ({signal_1408, signal_836}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_78 ( .a ({1'b0, 1'b0}), .b ({signal_1216, signal_804}), .c ({signal_1331, signal_276}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_79 ( .a ({signal_1333, signal_277}), .b ({signal_1332, signal_278}), .c ({signal_1409, signal_819}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_80 ( .a ({signal_1186, signal_851}), .b ({signal_1154, signal_867}), .c ({signal_1332, signal_278}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_81 ( .a ({1'b0, 1'b0}), .b ({signal_1250, signal_787}), .c ({signal_1333, signal_277}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_82 ( .a ({signal_1334, signal_279}), .b ({signal_1154, signal_867}), .c ({signal_1410, signal_835}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_83 ( .a ({1'b0, 1'b0}), .b ({signal_1218, signal_803}), .c ({signal_1334, signal_279}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_84 ( .a ({signal_1336, signal_280}), .b ({signal_1335, signal_281}), .c ({signal_1411, signal_818}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_85 ( .a ({signal_1188, signal_850}), .b ({signal_1156, signal_866}), .c ({signal_1335, signal_281}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_86 ( .a ({1'b0, 1'b0}), .b ({signal_1252, signal_786}), .c ({signal_1336, signal_280}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_87 ( .a ({signal_1337, signal_282}), .b ({signal_1156, signal_866}), .c ({signal_1412, signal_834}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_88 ( .a ({1'b0, 1'b0}), .b ({signal_1220, signal_802}), .c ({signal_1337, signal_282}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_89 ( .a ({signal_1339, signal_283}), .b ({signal_1338, signal_284}), .c ({signal_1413, signal_817}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_90 ( .a ({signal_1190, signal_849}), .b ({signal_1158, signal_865}), .c ({signal_1338, signal_284}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_91 ( .a ({1'b0, 1'b0}), .b ({signal_1254, signal_785}), .c ({signal_1339, signal_283}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_92 ( .a ({signal_1340, signal_285}), .b ({signal_1158, signal_865}), .c ({signal_1414, signal_833}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_93 ( .a ({1'b0, 1'b0}), .b ({signal_1222, signal_801}), .c ({signal_1340, signal_285}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_94 ( .a ({signal_1342, signal_286}), .b ({signal_1341, signal_287}), .c ({signal_1415, signal_816}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_95 ( .a ({signal_1192, signal_848}), .b ({signal_1160, signal_864}), .c ({signal_1341, signal_287}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_96 ( .a ({1'b0, 1'b0}), .b ({signal_1256, signal_784}), .c ({signal_1342, signal_286}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_97 ( .a ({signal_1343, signal_288}), .b ({signal_1160, signal_864}), .c ({signal_1416, signal_832}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_98 ( .a ({1'b0, 1'b0}), .b ({signal_1224, signal_800}), .c ({signal_1343, signal_288}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_99 ( .a ({signal_1345, signal_289}), .b ({signal_1344, signal_290}), .c ({signal_1417, signal_815}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_100 ( .a ({signal_1194, signal_847}), .b ({signal_1162, signal_863}), .c ({signal_1344, signal_290}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_101 ( .a ({1'b0, 1'b0}), .b ({signal_1258, signal_783}), .c ({signal_1345, signal_289}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_102 ( .a ({signal_1346, signal_291}), .b ({signal_1162, signal_863}), .c ({signal_1418, signal_831}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_103 ( .a ({1'b0, 1'b0}), .b ({signal_1226, signal_799}), .c ({signal_1346, signal_291}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_104 ( .a ({signal_1348, signal_292}), .b ({signal_1347, signal_293}), .c ({signal_1419, signal_814}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_105 ( .a ({signal_1196, signal_846}), .b ({signal_1164, signal_862}), .c ({signal_1347, signal_293}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_106 ( .a ({1'b0, 1'b0}), .b ({signal_1260, signal_782}), .c ({signal_1348, signal_292}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_107 ( .a ({signal_1349, signal_294}), .b ({signal_1164, signal_862}), .c ({signal_1420, signal_830}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_108 ( .a ({1'b0, 1'b0}), .b ({signal_1228, signal_798}), .c ({signal_1349, signal_294}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_109 ( .a ({signal_1351, signal_295}), .b ({signal_1350, signal_296}), .c ({signal_1421, signal_813}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_110 ( .a ({signal_1198, signal_845}), .b ({signal_1166, signal_861}), .c ({signal_1350, signal_296}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_111 ( .a ({1'b0, 1'b0}), .b ({signal_1262, signal_781}), .c ({signal_1351, signal_295}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_112 ( .a ({signal_1352, signal_297}), .b ({signal_1166, signal_861}), .c ({signal_1422, signal_829}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_113 ( .a ({1'b0, 1'b0}), .b ({signal_1230, signal_797}), .c ({signal_1352, signal_297}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_114 ( .a ({signal_1354, signal_298}), .b ({signal_1353, signal_299}), .c ({signal_1423, signal_812}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_115 ( .a ({signal_1200, signal_844}), .b ({signal_1168, signal_860}), .c ({signal_1353, signal_299}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_116 ( .a ({1'b0, 1'b0}), .b ({signal_1264, signal_780}), .c ({signal_1354, signal_298}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_117 ( .a ({signal_1355, signal_300}), .b ({signal_1168, signal_860}), .c ({signal_1424, signal_828}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_118 ( .a ({1'b0, 1'b0}), .b ({signal_1232, signal_796}), .c ({signal_1355, signal_300}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_119 ( .a ({signal_1357, signal_301}), .b ({signal_1356, signal_302}), .c ({signal_1425, signal_811}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_120 ( .a ({signal_1202, signal_843}), .b ({signal_1170, signal_859}), .c ({signal_1356, signal_302}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_121 ( .a ({1'b0, 1'b0}), .b ({signal_1266, signal_779}), .c ({signal_1357, signal_301}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_122 ( .a ({signal_1358, signal_303}), .b ({signal_1170, signal_859}), .c ({signal_1426, signal_827}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_123 ( .a ({1'b0, 1'b0}), .b ({signal_1234, signal_795}), .c ({signal_1358, signal_303}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_124 ( .a ({signal_1360, signal_304}), .b ({signal_1359, signal_305}), .c ({signal_1427, signal_810}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_125 ( .a ({signal_1204, signal_842}), .b ({signal_1172, signal_858}), .c ({signal_1359, signal_305}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_126 ( .a ({1'b0, 1'b0}), .b ({signal_1268, signal_778}), .c ({signal_1360, signal_304}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_127 ( .a ({signal_1361, signal_306}), .b ({signal_1172, signal_858}), .c ({signal_1428, signal_826}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_128 ( .a ({1'b0, 1'b0}), .b ({signal_1236, signal_794}), .c ({signal_1361, signal_306}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_129 ( .a ({signal_1363, signal_307}), .b ({signal_1362, signal_308}), .c ({signal_1429, signal_809}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_130 ( .a ({signal_1206, signal_841}), .b ({signal_1174, signal_857}), .c ({signal_1362, signal_308}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_131 ( .a ({1'b0, 1'b0}), .b ({signal_1270, signal_777}), .c ({signal_1363, signal_307}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_132 ( .a ({signal_1364, signal_309}), .b ({signal_1174, signal_857}), .c ({signal_1430, signal_825}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_133 ( .a ({1'b0, 1'b0}), .b ({signal_1238, signal_793}), .c ({signal_1364, signal_309}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_134 ( .a ({signal_1366, signal_310}), .b ({signal_1365, signal_311}), .c ({signal_1431, signal_808}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_135 ( .a ({signal_1208, signal_840}), .b ({signal_1176, signal_856}), .c ({signal_1365, signal_311}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_136 ( .a ({1'b0, 1'b0}), .b ({signal_1272, signal_776}), .c ({signal_1366, signal_310}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_137 ( .a ({signal_1367, signal_312}), .b ({signal_1176, signal_856}), .c ({signal_1432, signal_824}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_138 ( .a ({1'b0, 1'b0}), .b ({signal_1240, signal_792}), .c ({signal_1367, signal_312}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_139 ( .a ({signal_1369, signal_313}), .b ({signal_1368, signal_314}), .c ({signal_1433, signal_807}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_140 ( .a ({signal_1210, signal_839}), .b ({signal_1178, signal_855}), .c ({signal_1368, signal_314}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_141 ( .a ({1'b0, 1'b0}), .b ({signal_1274, signal_775}), .c ({signal_1369, signal_313}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_142 ( .a ({signal_1370, signal_315}), .b ({signal_1178, signal_855}), .c ({signal_1434, signal_823}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_143 ( .a ({1'b0, 1'b0}), .b ({signal_1242, signal_791}), .c ({signal_1370, signal_315}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_144 ( .a ({signal_1587, signal_316}), .b ({signal_2837, signal_2836}), .c ({signal_1651, signal_950}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_145 ( .a ({1'b0, 1'b0}), .b ({signal_1403, signal_822}), .c ({signal_1587, signal_316}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_146 ( .a ({signal_1588, signal_317}), .b ({signal_2839, signal_2838}), .c ({signal_1652, signal_949}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_147 ( .a ({1'b0, 1'b0}), .b ({signal_1405, signal_821}), .c ({signal_1588, signal_317}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_148 ( .a ({signal_1589, signal_318}), .b ({signal_2841, signal_2840}), .c ({signal_1653, signal_948}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_149 ( .a ({1'b0, 1'b0}), .b ({signal_1407, signal_820}), .c ({signal_1589, signal_318}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_150 ( .a ({signal_1590, signal_319}), .b ({signal_2843, signal_2842}), .c ({signal_1654, signal_947}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_151 ( .a ({1'b0, 1'b0}), .b ({signal_1409, signal_819}), .c ({signal_1590, signal_319}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_152 ( .a ({signal_1591, signal_320}), .b ({signal_2845, signal_2844}), .c ({signal_1655, signal_946}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_153 ( .a ({1'b0, 1'b0}), .b ({signal_1411, signal_818}), .c ({signal_1591, signal_320}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_154 ( .a ({signal_1592, signal_321}), .b ({signal_2847, signal_2846}), .c ({signal_1656, signal_945}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_155 ( .a ({1'b0, 1'b0}), .b ({signal_1413, signal_817}), .c ({signal_1592, signal_321}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_156 ( .a ({signal_1593, signal_322}), .b ({signal_2849, signal_2848}), .c ({signal_1657, signal_944}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_157 ( .a ({1'b0, 1'b0}), .b ({signal_1415, signal_816}), .c ({signal_1593, signal_322}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_158 ( .a ({signal_1594, signal_323}), .b ({signal_2851, signal_2850}), .c ({signal_1658, signal_943}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_159 ( .a ({1'b0, 1'b0}), .b ({signal_1417, signal_815}), .c ({signal_1594, signal_323}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_160 ( .a ({signal_1595, signal_324}), .b ({signal_2853, signal_2852}), .c ({signal_1659, signal_942}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_161 ( .a ({1'b0, 1'b0}), .b ({signal_1419, signal_814}), .c ({signal_1595, signal_324}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_162 ( .a ({signal_1596, signal_325}), .b ({signal_2855, signal_2854}), .c ({signal_1660, signal_941}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_163 ( .a ({1'b0, 1'b0}), .b ({signal_1421, signal_813}), .c ({signal_1596, signal_325}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_164 ( .a ({signal_1597, signal_326}), .b ({signal_2857, signal_2856}), .c ({signal_1661, signal_940}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_165 ( .a ({1'b0, 1'b0}), .b ({signal_1423, signal_812}), .c ({signal_1597, signal_326}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_166 ( .a ({signal_1598, signal_327}), .b ({signal_2859, signal_2858}), .c ({signal_1662, signal_939}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_167 ( .a ({1'b0, 1'b0}), .b ({signal_1425, signal_811}), .c ({signal_1598, signal_327}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_168 ( .a ({signal_1599, signal_328}), .b ({signal_2861, signal_2860}), .c ({signal_1663, signal_938}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_169 ( .a ({1'b0, 1'b0}), .b ({signal_1427, signal_810}), .c ({signal_1599, signal_328}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_170 ( .a ({signal_1600, signal_329}), .b ({signal_2863, signal_2862}), .c ({signal_1664, signal_937}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_171 ( .a ({1'b0, 1'b0}), .b ({signal_1429, signal_809}), .c ({signal_1600, signal_329}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_172 ( .a ({signal_1601, signal_330}), .b ({signal_2865, signal_2864}), .c ({signal_1665, signal_936}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_173 ( .a ({1'b0, 1'b0}), .b ({signal_1431, signal_808}), .c ({signal_1601, signal_330}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_174 ( .a ({signal_1602, signal_331}), .b ({signal_2867, signal_2866}), .c ({signal_1666, signal_935}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_175 ( .a ({1'b0, 1'b0}), .b ({signal_1433, signal_807}), .c ({signal_1602, signal_331}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_176 ( .a ({signal_1604, signal_332}), .b ({signal_2869, signal_2868}), .c ({signal_1667, signal_958}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_178 ( .a ({1'b0, 1'b0}), .b ({signal_1420, signal_830}), .c ({signal_1604, signal_332}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_179 ( .a ({signal_1606, signal_334}), .b ({signal_2871, signal_2870}), .c ({signal_1668, signal_957}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_181 ( .a ({1'b0, 1'b0}), .b ({signal_1422, signal_829}), .c ({signal_1606, signal_334}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_182 ( .a ({signal_1608, signal_336}), .b ({signal_2873, signal_2872}), .c ({signal_1669, signal_956}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_184 ( .a ({1'b0, 1'b0}), .b ({signal_1424, signal_828}), .c ({signal_1608, signal_336}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_185 ( .a ({signal_1610, signal_338}), .b ({signal_2875, signal_2874}), .c ({signal_1670, signal_955}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_187 ( .a ({1'b0, 1'b0}), .b ({signal_1426, signal_827}), .c ({signal_1610, signal_338}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_188 ( .a ({signal_1612, signal_340}), .b ({signal_2877, signal_2876}), .c ({signal_1671, signal_954}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_190 ( .a ({1'b0, 1'b0}), .b ({signal_1428, signal_826}), .c ({signal_1612, signal_340}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_191 ( .a ({signal_1614, signal_342}), .b ({signal_2879, signal_2878}), .c ({signal_1672, signal_953}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_193 ( .a ({1'b0, 1'b0}), .b ({signal_1430, signal_825}), .c ({signal_1614, signal_342}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_194 ( .a ({signal_1616, signal_344}), .b ({signal_2881, signal_2880}), .c ({signal_1673, signal_952}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_196 ( .a ({1'b0, 1'b0}), .b ({signal_1432, signal_824}), .c ({signal_1616, signal_344}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_197 ( .a ({signal_1618, signal_346}), .b ({signal_2883, signal_2882}), .c ({signal_1674, signal_951}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_199 ( .a ({1'b0, 1'b0}), .b ({signal_1434, signal_823}), .c ({signal_1618, signal_346}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_200 ( .a ({signal_1371, signal_348}), .b ({signal_2885, signal_2884}), .c ({signal_1435, signal_998}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_201 ( .a ({1'b0, 1'b0}), .b ({signal_1148, signal_870}), .c ({signal_1371, signal_348}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_202 ( .a ({signal_1372, signal_349}), .b ({signal_2887, signal_2886}), .c ({signal_1619, signal_997}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_203 ( .a ({1'b0, 1'b0}), .b ({signal_1150, signal_869}), .c ({signal_1372, signal_349}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_204 ( .a ({signal_1373, signal_350}), .b ({signal_2889, signal_2888}), .c ({signal_1436, signal_996}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_205 ( .a ({1'b0, 1'b0}), .b ({signal_1152, signal_868}), .c ({signal_1373, signal_350}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_206 ( .a ({signal_1374, signal_351}), .b ({signal_2891, signal_2890}), .c ({signal_1620, signal_995}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_207 ( .a ({1'b0, 1'b0}), .b ({signal_1154, signal_867}), .c ({signal_1374, signal_351}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_208 ( .a ({signal_1375, signal_352}), .b ({signal_2893, signal_2892}), .c ({signal_1621, signal_994}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_209 ( .a ({1'b0, 1'b0}), .b ({signal_1156, signal_866}), .c ({signal_1375, signal_352}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_210 ( .a ({signal_1376, signal_353}), .b ({signal_2895, signal_2894}), .c ({signal_1622, signal_993}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_211 ( .a ({1'b0, 1'b0}), .b ({signal_1158, signal_865}), .c ({signal_1376, signal_353}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_212 ( .a ({signal_1377, signal_354}), .b ({signal_2897, signal_2896}), .c ({signal_1623, signal_992}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_213 ( .a ({1'b0, 1'b0}), .b ({signal_1160, signal_864}), .c ({signal_1377, signal_354}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_214 ( .a ({signal_1378, signal_355}), .b ({signal_2899, signal_2898}), .c ({signal_1624, signal_991}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_215 ( .a ({1'b0, 1'b0}), .b ({signal_1162, signal_863}), .c ({signal_1378, signal_355}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_216 ( .a ({signal_1379, signal_356}), .b ({signal_2901, signal_2900}), .c ({signal_1625, signal_990}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_217 ( .a ({1'b0, 1'b0}), .b ({signal_1164, signal_862}), .c ({signal_1379, signal_356}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_218 ( .a ({signal_1380, signal_357}), .b ({signal_2903, signal_2902}), .c ({signal_1626, signal_989}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_219 ( .a ({1'b0, 1'b0}), .b ({signal_1166, signal_861}), .c ({signal_1380, signal_357}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_220 ( .a ({signal_1381, signal_358}), .b ({signal_2905, signal_2904}), .c ({signal_1627, signal_988}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_221 ( .a ({1'b0, 1'b0}), .b ({signal_1168, signal_860}), .c ({signal_1381, signal_358}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_222 ( .a ({signal_1382, signal_359}), .b ({signal_2907, signal_2906}), .c ({signal_1628, signal_987}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_223 ( .a ({1'b0, 1'b0}), .b ({signal_1170, signal_859}), .c ({signal_1382, signal_359}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_224 ( .a ({signal_1383, signal_360}), .b ({signal_2909, signal_2908}), .c ({signal_1629, signal_986}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_225 ( .a ({1'b0, 1'b0}), .b ({signal_1172, signal_858}), .c ({signal_1383, signal_360}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_226 ( .a ({signal_1384, signal_361}), .b ({signal_2911, signal_2910}), .c ({signal_1630, signal_985}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_227 ( .a ({1'b0, 1'b0}), .b ({signal_1174, signal_857}), .c ({signal_1384, signal_361}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_228 ( .a ({signal_1385, signal_362}), .b ({signal_2913, signal_2912}), .c ({signal_1631, signal_984}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_229 ( .a ({1'b0, 1'b0}), .b ({signal_1176, signal_856}), .c ({signal_1385, signal_362}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_230 ( .a ({signal_1386, signal_363}), .b ({signal_2915, signal_2914}), .c ({signal_1632, signal_983}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_231 ( .a ({1'b0, 1'b0}), .b ({signal_1178, signal_855}), .c ({signal_1386, signal_363}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_232 ( .a ({signal_1387, signal_364}), .b ({signal_2917, signal_2916}), .c ({signal_1633, signal_982}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_233 ( .a ({1'b0, 1'b0}), .b ({signal_1180, signal_854}), .c ({signal_1387, signal_364}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_234 ( .a ({signal_1388, signal_365}), .b ({signal_2919, signal_2918}), .c ({signal_1634, signal_981}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_235 ( .a ({1'b0, 1'b0}), .b ({signal_1182, signal_853}), .c ({signal_1388, signal_365}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_236 ( .a ({signal_1389, signal_366}), .b ({signal_2921, signal_2920}), .c ({signal_1635, signal_980}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_237 ( .a ({1'b0, 1'b0}), .b ({signal_1184, signal_852}), .c ({signal_1389, signal_366}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_238 ( .a ({signal_1390, signal_367}), .b ({signal_2923, signal_2922}), .c ({signal_1636, signal_979}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_239 ( .a ({1'b0, 1'b0}), .b ({signal_1186, signal_851}), .c ({signal_1390, signal_367}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_240 ( .a ({signal_1391, signal_368}), .b ({signal_2925, signal_2924}), .c ({signal_1637, signal_978}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_241 ( .a ({1'b0, 1'b0}), .b ({signal_1188, signal_850}), .c ({signal_1391, signal_368}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_242 ( .a ({signal_1392, signal_369}), .b ({signal_2927, signal_2926}), .c ({signal_1638, signal_977}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_243 ( .a ({1'b0, 1'b0}), .b ({signal_1190, signal_849}), .c ({signal_1392, signal_369}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_244 ( .a ({signal_1393, signal_370}), .b ({signal_2929, signal_2928}), .c ({signal_1437, signal_976}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_245 ( .a ({1'b0, 1'b0}), .b ({signal_1192, signal_848}), .c ({signal_1393, signal_370}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_246 ( .a ({signal_1394, signal_371}), .b ({signal_2931, signal_2930}), .c ({signal_1438, signal_975}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_247 ( .a ({1'b0, 1'b0}), .b ({signal_1194, signal_847}), .c ({signal_1394, signal_371}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_248 ( .a ({signal_1395, signal_372}), .b ({signal_2933, signal_2932}), .c ({signal_1439, signal_974}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_249 ( .a ({1'b0, 1'b0}), .b ({signal_1196, signal_846}), .c ({signal_1395, signal_372}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_250 ( .a ({signal_1396, signal_373}), .b ({signal_2935, signal_2934}), .c ({signal_1440, signal_973}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_251 ( .a ({1'b0, 1'b0}), .b ({signal_1198, signal_845}), .c ({signal_1396, signal_373}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_252 ( .a ({signal_1397, signal_374}), .b ({signal_2937, signal_2936}), .c ({signal_1441, signal_972}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_253 ( .a ({1'b0, 1'b0}), .b ({signal_1200, signal_844}), .c ({signal_1397, signal_374}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_254 ( .a ({signal_1398, signal_375}), .b ({signal_2939, signal_2938}), .c ({signal_1442, signal_971}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_255 ( .a ({1'b0, 1'b0}), .b ({signal_1202, signal_843}), .c ({signal_1398, signal_375}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_256 ( .a ({signal_1399, signal_376}), .b ({signal_2941, signal_2940}), .c ({signal_1639, signal_970}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_257 ( .a ({1'b0, 1'b0}), .b ({signal_1204, signal_842}), .c ({signal_1399, signal_376}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_258 ( .a ({signal_1400, signal_377}), .b ({signal_2943, signal_2942}), .c ({signal_1640, signal_969}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_259 ( .a ({1'b0, 1'b0}), .b ({signal_1206, signal_841}), .c ({signal_1400, signal_377}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_260 ( .a ({signal_1401, signal_378}), .b ({signal_2945, signal_2944}), .c ({signal_1641, signal_968}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_261 ( .a ({1'b0, 1'b0}), .b ({signal_1208, signal_840}), .c ({signal_1401, signal_378}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_262 ( .a ({signal_1402, signal_379}), .b ({signal_2947, signal_2946}), .c ({signal_1642, signal_967}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_263 ( .a ({1'b0, 1'b0}), .b ({signal_1210, signal_839}), .c ({signal_1402, signal_379}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_264 ( .a ({signal_1643, signal_380}), .b ({signal_2949, signal_2948}), .c ({signal_1675, signal_966}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_265 ( .a ({1'b0, 1'b0}), .b ({signal_1404, signal_838}), .c ({signal_1643, signal_380}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_266 ( .a ({signal_1644, signal_381}), .b ({signal_2951, signal_2950}), .c ({signal_1676, signal_965}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_267 ( .a ({1'b0, 1'b0}), .b ({signal_1406, signal_837}), .c ({signal_1644, signal_381}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_268 ( .a ({signal_1645, signal_382}), .b ({signal_2953, signal_2952}), .c ({signal_1677, signal_964}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_269 ( .a ({1'b0, 1'b0}), .b ({signal_1408, signal_836}), .c ({signal_1645, signal_382}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_270 ( .a ({signal_1646, signal_383}), .b ({signal_2955, signal_2954}), .c ({signal_1678, signal_963}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_271 ( .a ({1'b0, 1'b0}), .b ({signal_1410, signal_835}), .c ({signal_1646, signal_383}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_272 ( .a ({signal_1647, signal_384}), .b ({signal_2957, signal_2956}), .c ({signal_1679, signal_962}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_273 ( .a ({1'b0, 1'b0}), .b ({signal_1412, signal_834}), .c ({signal_1647, signal_384}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_274 ( .a ({signal_1648, signal_385}), .b ({signal_2959, signal_2958}), .c ({signal_1680, signal_961}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_275 ( .a ({1'b0, 1'b0}), .b ({signal_1414, signal_833}), .c ({signal_1648, signal_385}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_276 ( .a ({signal_1649, signal_386}), .b ({signal_2961, signal_2960}), .c ({signal_1681, signal_960}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_277 ( .a ({1'b0, 1'b0}), .b ({signal_1416, signal_832}), .c ({signal_1649, signal_386}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_278 ( .a ({signal_1650, signal_387}), .b ({signal_2963, signal_2962}), .c ({signal_1682, signal_959}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_279 ( .a ({1'b0, 1'b0}), .b ({signal_1418, signal_831}), .c ({signal_1650, signal_387}) ) ;
    CRAFT_step2_ANF #(.low_latency(1), .pipeline(1)) cell_819 ( .in0 ({ciphertext_s0[0], ciphertext_s0[1], ciphertext_s0[2], ciphertext_s0[3], ciphertext_s0[4], ciphertext_s0[5], ciphertext_s0[6], ciphertext_s0[7], ciphertext_s0[8], ciphertext_s0[9], ciphertext_s0[10], ciphertext_s0[11], ciphertext_s0[12], ciphertext_s0[13], ciphertext_s0[14], ciphertext_s0[15], ciphertext_s0[16], ciphertext_s0[17], ciphertext_s0[18], ciphertext_s0[19], ciphertext_s0[20], ciphertext_s0[21], ciphertext_s0[22], ciphertext_s0[23], ciphertext_s0[24], ciphertext_s0[25], ciphertext_s0[26], ciphertext_s0[27], ciphertext_s0[28], ciphertext_s0[29], ciphertext_s0[30], ciphertext_s0[31], ciphertext_s0[32], ciphertext_s0[33], ciphertext_s0[34], ciphertext_s0[35], ciphertext_s0[36], ciphertext_s0[37], ciphertext_s0[38], ciphertext_s0[39], ciphertext_s0[40], ciphertext_s0[41], ciphertext_s0[42], ciphertext_s0[43], ciphertext_s0[44], ciphertext_s0[45], ciphertext_s0[46], ciphertext_s0[47], ciphertext_s0[48], ciphertext_s0[49], ciphertext_s0[50], ciphertext_s0[51], ciphertext_s0[52], ciphertext_s0[53], ciphertext_s0[54], ciphertext_s0[55], ciphertext_s0[56], ciphertext_s0[57], ciphertext_s0[58], ciphertext_s0[59], ciphertext_s0[60], ciphertext_s0[61], ciphertext_s0[62], ciphertext_s0[63]}), .in1 ({ciphertext_s1[0], ciphertext_s1[1], ciphertext_s1[2], ciphertext_s1[3], ciphertext_s1[4], ciphertext_s1[5], ciphertext_s1[6], ciphertext_s1[7], ciphertext_s1[8], ciphertext_s1[9], ciphertext_s1[10], ciphertext_s1[11], ciphertext_s1[12], ciphertext_s1[13], ciphertext_s1[14], ciphertext_s1[15], ciphertext_s1[16], ciphertext_s1[17], ciphertext_s1[18], ciphertext_s1[19], ciphertext_s1[20], ciphertext_s1[21], ciphertext_s1[22], ciphertext_s1[23], ciphertext_s1[24], ciphertext_s1[25], ciphertext_s1[26], ciphertext_s1[27], ciphertext_s1[28], ciphertext_s1[29], ciphertext_s1[30], ciphertext_s1[31], ciphertext_s1[32], ciphertext_s1[33], ciphertext_s1[34], ciphertext_s1[35], ciphertext_s1[36], ciphertext_s1[37], ciphertext_s1[38], ciphertext_s1[39], ciphertext_s1[40], ciphertext_s1[41], ciphertext_s1[42], ciphertext_s1[43], ciphertext_s1[44], ciphertext_s1[45], ciphertext_s1[46], ciphertext_s1[47], ciphertext_s1[48], ciphertext_s1[49], ciphertext_s1[50], ciphertext_s1[51], ciphertext_s1[52], ciphertext_s1[53], ciphertext_s1[54], ciphertext_s1[55], ciphertext_s1[56], ciphertext_s1[57], ciphertext_s1[58], ciphertext_s1[59], ciphertext_s1[60], ciphertext_s1[61], ciphertext_s1[62], ciphertext_s1[63]}), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960], Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720], Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480], Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240], Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_774, signal_773, signal_772, signal_771, signal_770, signal_769, signal_768, signal_767, signal_766, signal_765, signal_764, signal_763, signal_762, signal_761, signal_760, signal_759, signal_758, signal_757, signal_756, signal_755, signal_754, signal_753, signal_752, signal_751, signal_750, signal_749, signal_748, signal_747, signal_746, signal_745, signal_744, signal_743, signal_742, signal_741, signal_740, signal_739, signal_738, signal_737, signal_736, signal_735, signal_734, signal_733, signal_732, signal_731, signal_730, signal_729, signal_728, signal_727, signal_726, signal_725, signal_724, signal_723, signal_722, signal_721, signal_720, signal_719, signal_718, signal_717, signal_716, signal_715, signal_714, signal_713, signal_712, signal_711}), .out1 ({signal_1146, signal_1145, signal_1144, signal_1143, signal_1142, signal_1141, signal_1140, signal_1139, signal_1138, signal_1137, signal_1136, signal_1135, signal_1134, signal_1133, signal_1132, signal_1131, signal_1130, signal_1129, signal_1128, signal_1127, signal_1126, signal_1125, signal_1124, signal_1123, signal_1122, signal_1121, signal_1120, signal_1119, signal_1118, signal_1117, signal_1116, signal_1115, signal_1114, signal_1113, signal_1112, signal_1111, signal_1110, signal_1109, signal_1108, signal_1107, signal_1106, signal_1105, signal_1104, signal_1103, signal_1102, signal_1101, signal_1100, signal_1099, signal_1098, signal_1097, signal_1096, signal_1095, signal_1094, signal_1093, signal_1092, signal_1091, signal_1090, signal_1089, signal_1088, signal_1087, signal_1086, signal_1085, signal_1084, signal_1083}) ) ;
    buf_clk cell_820 ( .C (clk), .D (rst), .Q (signal_2707) ) ;
    buf_clk cell_821 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_2708) ) ;
    buf_clk cell_822 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_2709) ) ;
    buf_clk cell_823 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_2710) ) ;
    buf_clk cell_824 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_2711) ) ;
    buf_clk cell_825 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_2712) ) ;
    buf_clk cell_826 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_2713) ) ;
    buf_clk cell_827 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_2714) ) ;
    buf_clk cell_828 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_2715) ) ;
    buf_clk cell_829 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_2716) ) ;
    buf_clk cell_830 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_2717) ) ;
    buf_clk cell_831 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_2718) ) ;
    buf_clk cell_832 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_2719) ) ;
    buf_clk cell_833 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_2720) ) ;
    buf_clk cell_834 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_2721) ) ;
    buf_clk cell_835 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_2722) ) ;
    buf_clk cell_836 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_2723) ) ;
    buf_clk cell_837 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_2724) ) ;
    buf_clk cell_838 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_2725) ) ;
    buf_clk cell_839 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_2726) ) ;
    buf_clk cell_840 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_2727) ) ;
    buf_clk cell_841 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_2728) ) ;
    buf_clk cell_842 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_2729) ) ;
    buf_clk cell_843 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_2730) ) ;
    buf_clk cell_844 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_2731) ) ;
    buf_clk cell_845 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_2732) ) ;
    buf_clk cell_846 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_2733) ) ;
    buf_clk cell_847 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_2734) ) ;
    buf_clk cell_848 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_2735) ) ;
    buf_clk cell_849 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_2736) ) ;
    buf_clk cell_850 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_2737) ) ;
    buf_clk cell_851 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_2738) ) ;
    buf_clk cell_852 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_2739) ) ;
    buf_clk cell_853 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_2740) ) ;
    buf_clk cell_854 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_2741) ) ;
    buf_clk cell_855 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_2742) ) ;
    buf_clk cell_856 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_2743) ) ;
    buf_clk cell_857 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_2744) ) ;
    buf_clk cell_858 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_2745) ) ;
    buf_clk cell_859 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_2746) ) ;
    buf_clk cell_860 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_2747) ) ;
    buf_clk cell_861 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_2748) ) ;
    buf_clk cell_862 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_2749) ) ;
    buf_clk cell_863 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_2750) ) ;
    buf_clk cell_864 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_2751) ) ;
    buf_clk cell_865 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_2752) ) ;
    buf_clk cell_866 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_2753) ) ;
    buf_clk cell_867 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_2754) ) ;
    buf_clk cell_868 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_2755) ) ;
    buf_clk cell_869 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_2756) ) ;
    buf_clk cell_870 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_2757) ) ;
    buf_clk cell_871 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_2758) ) ;
    buf_clk cell_872 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_2759) ) ;
    buf_clk cell_873 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_2760) ) ;
    buf_clk cell_874 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_2761) ) ;
    buf_clk cell_875 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_2762) ) ;
    buf_clk cell_876 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_2763) ) ;
    buf_clk cell_877 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_2764) ) ;
    buf_clk cell_878 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_2765) ) ;
    buf_clk cell_879 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_2766) ) ;
    buf_clk cell_880 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_2767) ) ;
    buf_clk cell_881 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_2768) ) ;
    buf_clk cell_882 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_2769) ) ;
    buf_clk cell_883 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_2770) ) ;
    buf_clk cell_884 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_2771) ) ;
    buf_clk cell_885 ( .C (clk), .D (plaintext_s0[32]), .Q (signal_2772) ) ;
    buf_clk cell_886 ( .C (clk), .D (plaintext_s1[32]), .Q (signal_2773) ) ;
    buf_clk cell_887 ( .C (clk), .D (plaintext_s0[33]), .Q (signal_2774) ) ;
    buf_clk cell_888 ( .C (clk), .D (plaintext_s1[33]), .Q (signal_2775) ) ;
    buf_clk cell_889 ( .C (clk), .D (plaintext_s0[34]), .Q (signal_2776) ) ;
    buf_clk cell_890 ( .C (clk), .D (plaintext_s1[34]), .Q (signal_2777) ) ;
    buf_clk cell_891 ( .C (clk), .D (plaintext_s0[35]), .Q (signal_2778) ) ;
    buf_clk cell_892 ( .C (clk), .D (plaintext_s1[35]), .Q (signal_2779) ) ;
    buf_clk cell_893 ( .C (clk), .D (plaintext_s0[36]), .Q (signal_2780) ) ;
    buf_clk cell_894 ( .C (clk), .D (plaintext_s1[36]), .Q (signal_2781) ) ;
    buf_clk cell_895 ( .C (clk), .D (plaintext_s0[37]), .Q (signal_2782) ) ;
    buf_clk cell_896 ( .C (clk), .D (plaintext_s1[37]), .Q (signal_2783) ) ;
    buf_clk cell_897 ( .C (clk), .D (plaintext_s0[38]), .Q (signal_2784) ) ;
    buf_clk cell_898 ( .C (clk), .D (plaintext_s1[38]), .Q (signal_2785) ) ;
    buf_clk cell_899 ( .C (clk), .D (plaintext_s0[39]), .Q (signal_2786) ) ;
    buf_clk cell_900 ( .C (clk), .D (plaintext_s1[39]), .Q (signal_2787) ) ;
    buf_clk cell_901 ( .C (clk), .D (plaintext_s0[40]), .Q (signal_2788) ) ;
    buf_clk cell_902 ( .C (clk), .D (plaintext_s1[40]), .Q (signal_2789) ) ;
    buf_clk cell_903 ( .C (clk), .D (plaintext_s0[41]), .Q (signal_2790) ) ;
    buf_clk cell_904 ( .C (clk), .D (plaintext_s1[41]), .Q (signal_2791) ) ;
    buf_clk cell_905 ( .C (clk), .D (plaintext_s0[42]), .Q (signal_2792) ) ;
    buf_clk cell_906 ( .C (clk), .D (plaintext_s1[42]), .Q (signal_2793) ) ;
    buf_clk cell_907 ( .C (clk), .D (plaintext_s0[43]), .Q (signal_2794) ) ;
    buf_clk cell_908 ( .C (clk), .D (plaintext_s1[43]), .Q (signal_2795) ) ;
    buf_clk cell_909 ( .C (clk), .D (plaintext_s0[44]), .Q (signal_2796) ) ;
    buf_clk cell_910 ( .C (clk), .D (plaintext_s1[44]), .Q (signal_2797) ) ;
    buf_clk cell_911 ( .C (clk), .D (plaintext_s0[45]), .Q (signal_2798) ) ;
    buf_clk cell_912 ( .C (clk), .D (plaintext_s1[45]), .Q (signal_2799) ) ;
    buf_clk cell_913 ( .C (clk), .D (plaintext_s0[46]), .Q (signal_2800) ) ;
    buf_clk cell_914 ( .C (clk), .D (plaintext_s1[46]), .Q (signal_2801) ) ;
    buf_clk cell_915 ( .C (clk), .D (plaintext_s0[47]), .Q (signal_2802) ) ;
    buf_clk cell_916 ( .C (clk), .D (plaintext_s1[47]), .Q (signal_2803) ) ;
    buf_clk cell_917 ( .C (clk), .D (plaintext_s0[48]), .Q (signal_2804) ) ;
    buf_clk cell_918 ( .C (clk), .D (plaintext_s1[48]), .Q (signal_2805) ) ;
    buf_clk cell_919 ( .C (clk), .D (plaintext_s0[49]), .Q (signal_2806) ) ;
    buf_clk cell_920 ( .C (clk), .D (plaintext_s1[49]), .Q (signal_2807) ) ;
    buf_clk cell_921 ( .C (clk), .D (plaintext_s0[50]), .Q (signal_2808) ) ;
    buf_clk cell_922 ( .C (clk), .D (plaintext_s1[50]), .Q (signal_2809) ) ;
    buf_clk cell_923 ( .C (clk), .D (plaintext_s0[51]), .Q (signal_2810) ) ;
    buf_clk cell_924 ( .C (clk), .D (plaintext_s1[51]), .Q (signal_2811) ) ;
    buf_clk cell_925 ( .C (clk), .D (plaintext_s0[52]), .Q (signal_2812) ) ;
    buf_clk cell_926 ( .C (clk), .D (plaintext_s1[52]), .Q (signal_2813) ) ;
    buf_clk cell_927 ( .C (clk), .D (plaintext_s0[53]), .Q (signal_2814) ) ;
    buf_clk cell_928 ( .C (clk), .D (plaintext_s1[53]), .Q (signal_2815) ) ;
    buf_clk cell_929 ( .C (clk), .D (plaintext_s0[54]), .Q (signal_2816) ) ;
    buf_clk cell_930 ( .C (clk), .D (plaintext_s1[54]), .Q (signal_2817) ) ;
    buf_clk cell_931 ( .C (clk), .D (plaintext_s0[55]), .Q (signal_2818) ) ;
    buf_clk cell_932 ( .C (clk), .D (plaintext_s1[55]), .Q (signal_2819) ) ;
    buf_clk cell_933 ( .C (clk), .D (plaintext_s0[56]), .Q (signal_2820) ) ;
    buf_clk cell_934 ( .C (clk), .D (plaintext_s1[56]), .Q (signal_2821) ) ;
    buf_clk cell_935 ( .C (clk), .D (plaintext_s0[57]), .Q (signal_2822) ) ;
    buf_clk cell_936 ( .C (clk), .D (plaintext_s1[57]), .Q (signal_2823) ) ;
    buf_clk cell_937 ( .C (clk), .D (plaintext_s0[58]), .Q (signal_2824) ) ;
    buf_clk cell_938 ( .C (clk), .D (plaintext_s1[58]), .Q (signal_2825) ) ;
    buf_clk cell_939 ( .C (clk), .D (plaintext_s0[59]), .Q (signal_2826) ) ;
    buf_clk cell_940 ( .C (clk), .D (plaintext_s1[59]), .Q (signal_2827) ) ;
    buf_clk cell_941 ( .C (clk), .D (plaintext_s0[60]), .Q (signal_2828) ) ;
    buf_clk cell_942 ( .C (clk), .D (plaintext_s1[60]), .Q (signal_2829) ) ;
    buf_clk cell_943 ( .C (clk), .D (plaintext_s0[61]), .Q (signal_2830) ) ;
    buf_clk cell_944 ( .C (clk), .D (plaintext_s1[61]), .Q (signal_2831) ) ;
    buf_clk cell_945 ( .C (clk), .D (plaintext_s0[62]), .Q (signal_2832) ) ;
    buf_clk cell_946 ( .C (clk), .D (plaintext_s1[62]), .Q (signal_2833) ) ;
    buf_clk cell_947 ( .C (clk), .D (plaintext_s0[63]), .Q (signal_2834) ) ;
    buf_clk cell_948 ( .C (clk), .D (plaintext_s1[63]), .Q (signal_2835) ) ;
    buf_clk cell_949 ( .C (clk), .D (signal_886), .Q (signal_2836) ) ;
    buf_clk cell_950 ( .C (clk), .D (signal_1556), .Q (signal_2837) ) ;
    buf_clk cell_951 ( .C (clk), .D (signal_885), .Q (signal_2838) ) ;
    buf_clk cell_952 ( .C (clk), .D (signal_1559), .Q (signal_2839) ) ;
    buf_clk cell_953 ( .C (clk), .D (signal_884), .Q (signal_2840) ) ;
    buf_clk cell_954 ( .C (clk), .D (signal_1562), .Q (signal_2841) ) ;
    buf_clk cell_955 ( .C (clk), .D (signal_883), .Q (signal_2842) ) ;
    buf_clk cell_956 ( .C (clk), .D (signal_1565), .Q (signal_2843) ) ;
    buf_clk cell_957 ( .C (clk), .D (signal_882), .Q (signal_2844) ) ;
    buf_clk cell_958 ( .C (clk), .D (signal_1568), .Q (signal_2845) ) ;
    buf_clk cell_959 ( .C (clk), .D (signal_881), .Q (signal_2846) ) ;
    buf_clk cell_960 ( .C (clk), .D (signal_1310), .Q (signal_2847) ) ;
    buf_clk cell_961 ( .C (clk), .D (signal_880), .Q (signal_2848) ) ;
    buf_clk cell_962 ( .C (clk), .D (signal_1313), .Q (signal_2849) ) ;
    buf_clk cell_963 ( .C (clk), .D (signal_879), .Q (signal_2850) ) ;
    buf_clk cell_964 ( .C (clk), .D (signal_1571), .Q (signal_2851) ) ;
    buf_clk cell_965 ( .C (clk), .D (signal_878), .Q (signal_2852) ) ;
    buf_clk cell_966 ( .C (clk), .D (signal_1316), .Q (signal_2853) ) ;
    buf_clk cell_967 ( .C (clk), .D (signal_877), .Q (signal_2854) ) ;
    buf_clk cell_968 ( .C (clk), .D (signal_1574), .Q (signal_2855) ) ;
    buf_clk cell_969 ( .C (clk), .D (signal_876), .Q (signal_2856) ) ;
    buf_clk cell_970 ( .C (clk), .D (signal_1577), .Q (signal_2857) ) ;
    buf_clk cell_971 ( .C (clk), .D (signal_875), .Q (signal_2858) ) ;
    buf_clk cell_972 ( .C (clk), .D (signal_1319), .Q (signal_2859) ) ;
    buf_clk cell_973 ( .C (clk), .D (signal_874), .Q (signal_2860) ) ;
    buf_clk cell_974 ( .C (clk), .D (signal_1580), .Q (signal_2861) ) ;
    buf_clk cell_975 ( .C (clk), .D (signal_873), .Q (signal_2862) ) ;
    buf_clk cell_976 ( .C (clk), .D (signal_1583), .Q (signal_2863) ) ;
    buf_clk cell_977 ( .C (clk), .D (signal_872), .Q (signal_2864) ) ;
    buf_clk cell_978 ( .C (clk), .D (signal_1322), .Q (signal_2865) ) ;
    buf_clk cell_979 ( .C (clk), .D (signal_871), .Q (signal_2866) ) ;
    buf_clk cell_980 ( .C (clk), .D (signal_1586), .Q (signal_2867) ) ;
    buf_clk cell_981 ( .C (clk), .D (signal_333), .Q (signal_2868) ) ;
    buf_clk cell_982 ( .C (clk), .D (signal_1603), .Q (signal_2869) ) ;
    buf_clk cell_983 ( .C (clk), .D (signal_335), .Q (signal_2870) ) ;
    buf_clk cell_984 ( .C (clk), .D (signal_1605), .Q (signal_2871) ) ;
    buf_clk cell_985 ( .C (clk), .D (signal_337), .Q (signal_2872) ) ;
    buf_clk cell_986 ( .C (clk), .D (signal_1607), .Q (signal_2873) ) ;
    buf_clk cell_987 ( .C (clk), .D (signal_339), .Q (signal_2874) ) ;
    buf_clk cell_988 ( .C (clk), .D (signal_1609), .Q (signal_2875) ) ;
    buf_clk cell_989 ( .C (clk), .D (signal_341), .Q (signal_2876) ) ;
    buf_clk cell_990 ( .C (clk), .D (signal_1611), .Q (signal_2877) ) ;
    buf_clk cell_991 ( .C (clk), .D (signal_343), .Q (signal_2878) ) ;
    buf_clk cell_992 ( .C (clk), .D (signal_1613), .Q (signal_2879) ) ;
    buf_clk cell_993 ( .C (clk), .D (signal_345), .Q (signal_2880) ) ;
    buf_clk cell_994 ( .C (clk), .D (signal_1615), .Q (signal_2881) ) ;
    buf_clk cell_995 ( .C (clk), .D (signal_347), .Q (signal_2882) ) ;
    buf_clk cell_996 ( .C (clk), .D (signal_1617), .Q (signal_2883) ) ;
    buf_clk cell_997 ( .C (clk), .D (signal_934), .Q (signal_2884) ) ;
    buf_clk cell_998 ( .C (clk), .D (signal_1277), .Q (signal_2885) ) ;
    buf_clk cell_999 ( .C (clk), .D (signal_933), .Q (signal_2886) ) ;
    buf_clk cell_1000 ( .C (clk), .D (signal_1445), .Q (signal_2887) ) ;
    buf_clk cell_1001 ( .C (clk), .D (signal_932), .Q (signal_2888) ) ;
    buf_clk cell_1002 ( .C (clk), .D (signal_1280), .Q (signal_2889) ) ;
    buf_clk cell_1003 ( .C (clk), .D (signal_931), .Q (signal_2890) ) ;
    buf_clk cell_1004 ( .C (clk), .D (signal_1448), .Q (signal_2891) ) ;
    buf_clk cell_1005 ( .C (clk), .D (signal_930), .Q (signal_2892) ) ;
    buf_clk cell_1006 ( .C (clk), .D (signal_1451), .Q (signal_2893) ) ;
    buf_clk cell_1007 ( .C (clk), .D (signal_929), .Q (signal_2894) ) ;
    buf_clk cell_1008 ( .C (clk), .D (signal_1454), .Q (signal_2895) ) ;
    buf_clk cell_1009 ( .C (clk), .D (signal_928), .Q (signal_2896) ) ;
    buf_clk cell_1010 ( .C (clk), .D (signal_1457), .Q (signal_2897) ) ;
    buf_clk cell_1011 ( .C (clk), .D (signal_927), .Q (signal_2898) ) ;
    buf_clk cell_1012 ( .C (clk), .D (signal_1460), .Q (signal_2899) ) ;
    buf_clk cell_1013 ( .C (clk), .D (signal_926), .Q (signal_2900) ) ;
    buf_clk cell_1014 ( .C (clk), .D (signal_1463), .Q (signal_2901) ) ;
    buf_clk cell_1015 ( .C (clk), .D (signal_925), .Q (signal_2902) ) ;
    buf_clk cell_1016 ( .C (clk), .D (signal_1466), .Q (signal_2903) ) ;
    buf_clk cell_1017 ( .C (clk), .D (signal_924), .Q (signal_2904) ) ;
    buf_clk cell_1018 ( .C (clk), .D (signal_1469), .Q (signal_2905) ) ;
    buf_clk cell_1019 ( .C (clk), .D (signal_923), .Q (signal_2906) ) ;
    buf_clk cell_1020 ( .C (clk), .D (signal_1472), .Q (signal_2907) ) ;
    buf_clk cell_1021 ( .C (clk), .D (signal_922), .Q (signal_2908) ) ;
    buf_clk cell_1022 ( .C (clk), .D (signal_1475), .Q (signal_2909) ) ;
    buf_clk cell_1023 ( .C (clk), .D (signal_921), .Q (signal_2910) ) ;
    buf_clk cell_1024 ( .C (clk), .D (signal_1478), .Q (signal_2911) ) ;
    buf_clk cell_1025 ( .C (clk), .D (signal_920), .Q (signal_2912) ) ;
    buf_clk cell_1026 ( .C (clk), .D (signal_1481), .Q (signal_2913) ) ;
    buf_clk cell_1027 ( .C (clk), .D (signal_919), .Q (signal_2914) ) ;
    buf_clk cell_1028 ( .C (clk), .D (signal_1484), .Q (signal_2915) ) ;
    buf_clk cell_1029 ( .C (clk), .D (signal_918), .Q (signal_2916) ) ;
    buf_clk cell_1030 ( .C (clk), .D (signal_1487), .Q (signal_2917) ) ;
    buf_clk cell_1031 ( .C (clk), .D (signal_917), .Q (signal_2918) ) ;
    buf_clk cell_1032 ( .C (clk), .D (signal_1490), .Q (signal_2919) ) ;
    buf_clk cell_1033 ( .C (clk), .D (signal_916), .Q (signal_2920) ) ;
    buf_clk cell_1034 ( .C (clk), .D (signal_1493), .Q (signal_2921) ) ;
    buf_clk cell_1035 ( .C (clk), .D (signal_915), .Q (signal_2922) ) ;
    buf_clk cell_1036 ( .C (clk), .D (signal_1496), .Q (signal_2923) ) ;
    buf_clk cell_1037 ( .C (clk), .D (signal_914), .Q (signal_2924) ) ;
    buf_clk cell_1038 ( .C (clk), .D (signal_1499), .Q (signal_2925) ) ;
    buf_clk cell_1039 ( .C (clk), .D (signal_913), .Q (signal_2926) ) ;
    buf_clk cell_1040 ( .C (clk), .D (signal_1502), .Q (signal_2927) ) ;
    buf_clk cell_1041 ( .C (clk), .D (signal_912), .Q (signal_2928) ) ;
    buf_clk cell_1042 ( .C (clk), .D (signal_1283), .Q (signal_2929) ) ;
    buf_clk cell_1043 ( .C (clk), .D (signal_911), .Q (signal_2930) ) ;
    buf_clk cell_1044 ( .C (clk), .D (signal_1286), .Q (signal_2931) ) ;
    buf_clk cell_1045 ( .C (clk), .D (signal_910), .Q (signal_2932) ) ;
    buf_clk cell_1046 ( .C (clk), .D (signal_1289), .Q (signal_2933) ) ;
    buf_clk cell_1047 ( .C (clk), .D (signal_909), .Q (signal_2934) ) ;
    buf_clk cell_1048 ( .C (clk), .D (signal_1292), .Q (signal_2935) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_908), .Q (signal_2936) ) ;
    buf_clk cell_1050 ( .C (clk), .D (signal_1295), .Q (signal_2937) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_907), .Q (signal_2938) ) ;
    buf_clk cell_1052 ( .C (clk), .D (signal_1298), .Q (signal_2939) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_906), .Q (signal_2940) ) ;
    buf_clk cell_1054 ( .C (clk), .D (signal_1505), .Q (signal_2941) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_905), .Q (signal_2942) ) ;
    buf_clk cell_1056 ( .C (clk), .D (signal_1508), .Q (signal_2943) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_904), .Q (signal_2944) ) ;
    buf_clk cell_1058 ( .C (clk), .D (signal_1511), .Q (signal_2945) ) ;
    buf_clk cell_1059 ( .C (clk), .D (signal_903), .Q (signal_2946) ) ;
    buf_clk cell_1060 ( .C (clk), .D (signal_1514), .Q (signal_2947) ) ;
    buf_clk cell_1061 ( .C (clk), .D (signal_902), .Q (signal_2948) ) ;
    buf_clk cell_1062 ( .C (clk), .D (signal_1517), .Q (signal_2949) ) ;
    buf_clk cell_1063 ( .C (clk), .D (signal_901), .Q (signal_2950) ) ;
    buf_clk cell_1064 ( .C (clk), .D (signal_1301), .Q (signal_2951) ) ;
    buf_clk cell_1065 ( .C (clk), .D (signal_900), .Q (signal_2952) ) ;
    buf_clk cell_1066 ( .C (clk), .D (signal_1520), .Q (signal_2953) ) ;
    buf_clk cell_1067 ( .C (clk), .D (signal_899), .Q (signal_2954) ) ;
    buf_clk cell_1068 ( .C (clk), .D (signal_1523), .Q (signal_2955) ) ;
    buf_clk cell_1069 ( .C (clk), .D (signal_898), .Q (signal_2956) ) ;
    buf_clk cell_1070 ( .C (clk), .D (signal_1304), .Q (signal_2957) ) ;
    buf_clk cell_1071 ( .C (clk), .D (signal_897), .Q (signal_2958) ) ;
    buf_clk cell_1072 ( .C (clk), .D (signal_1526), .Q (signal_2959) ) ;
    buf_clk cell_1073 ( .C (clk), .D (signal_896), .Q (signal_2960) ) ;
    buf_clk cell_1074 ( .C (clk), .D (signal_1529), .Q (signal_2961) ) ;
    buf_clk cell_1075 ( .C (clk), .D (signal_895), .Q (signal_2962) ) ;
    buf_clk cell_1076 ( .C (clk), .D (signal_1307), .Q (signal_2963) ) ;
    buf_clk cell_1077 ( .C (clk), .D (signal_1008), .Q (signal_2964) ) ;
    buf_clk cell_1078 ( .C (clk), .D (signal_1009), .Q (signal_2965) ) ;
    buf_clk cell_1079 ( .C (clk), .D (signal_1010), .Q (signal_2966) ) ;
    buf_clk cell_1080 ( .C (clk), .D (signal_1011), .Q (signal_2967) ) ;
    buf_clk cell_1081 ( .C (clk), .D (signal_1012), .Q (signal_2968) ) ;
    buf_clk cell_1082 ( .C (clk), .D (signal_1013), .Q (signal_2969) ) ;
    buf_clk cell_1083 ( .C (clk), .D (signal_1014), .Q (signal_2970) ) ;
    buf_clk cell_1084 ( .C (clk), .D (signal_1017), .Q (signal_2971) ) ;
    buf_clk cell_1085 ( .C (clk), .D (signal_1018), .Q (signal_2972) ) ;
    buf_clk cell_1086 ( .C (clk), .D (signal_267), .Q (signal_2973) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(1)) cell_281 ( .clk (clk), .D ({signal_1666, signal_935}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_283 ( .clk (clk), .D ({signal_1665, signal_936}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_285 ( .clk (clk), .D ({signal_1664, signal_937}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_287 ( .clk (clk), .D ({signal_1663, signal_938}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_289 ( .clk (clk), .D ({signal_1662, signal_939}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_291 ( .clk (clk), .D ({signal_1661, signal_940}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_293 ( .clk (clk), .D ({signal_1660, signal_941}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_295 ( .clk (clk), .D ({signal_1659, signal_942}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_297 ( .clk (clk), .D ({signal_1658, signal_943}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_299 ( .clk (clk), .D ({signal_1657, signal_944}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_301 ( .clk (clk), .D ({signal_1656, signal_945}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_303 ( .clk (clk), .D ({signal_1655, signal_946}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_305 ( .clk (clk), .D ({signal_1654, signal_947}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_307 ( .clk (clk), .D ({signal_1653, signal_948}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_309 ( .clk (clk), .D ({signal_1652, signal_949}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_311 ( .clk (clk), .D ({signal_1651, signal_950}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_313 ( .clk (clk), .D ({signal_1674, signal_951}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_315 ( .clk (clk), .D ({signal_1673, signal_952}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_317 ( .clk (clk), .D ({signal_1672, signal_953}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_319 ( .clk (clk), .D ({signal_1671, signal_954}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_321 ( .clk (clk), .D ({signal_1670, signal_955}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_323 ( .clk (clk), .D ({signal_1669, signal_956}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_325 ( .clk (clk), .D ({signal_1668, signal_957}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_327 ( .clk (clk), .D ({signal_1667, signal_958}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_329 ( .clk (clk), .D ({signal_1682, signal_959}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_331 ( .clk (clk), .D ({signal_1681, signal_960}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_333 ( .clk (clk), .D ({signal_1680, signal_961}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_335 ( .clk (clk), .D ({signal_1679, signal_962}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_337 ( .clk (clk), .D ({signal_1678, signal_963}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_339 ( .clk (clk), .D ({signal_1677, signal_964}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_341 ( .clk (clk), .D ({signal_1676, signal_965}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_343 ( .clk (clk), .D ({signal_1675, signal_966}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_345 ( .clk (clk), .D ({signal_1642, signal_967}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_347 ( .clk (clk), .D ({signal_1641, signal_968}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_349 ( .clk (clk), .D ({signal_1640, signal_969}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_351 ( .clk (clk), .D ({signal_1639, signal_970}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_353 ( .clk (clk), .D ({signal_1442, signal_971}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_355 ( .clk (clk), .D ({signal_1441, signal_972}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_357 ( .clk (clk), .D ({signal_1440, signal_973}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_359 ( .clk (clk), .D ({signal_1439, signal_974}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_361 ( .clk (clk), .D ({signal_1438, signal_975}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_363 ( .clk (clk), .D ({signal_1437, signal_976}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_365 ( .clk (clk), .D ({signal_1638, signal_977}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_367 ( .clk (clk), .D ({signal_1637, signal_978}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_369 ( .clk (clk), .D ({signal_1636, signal_979}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_371 ( .clk (clk), .D ({signal_1635, signal_980}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_373 ( .clk (clk), .D ({signal_1634, signal_981}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_375 ( .clk (clk), .D ({signal_1633, signal_982}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_377 ( .clk (clk), .D ({signal_1632, signal_983}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_379 ( .clk (clk), .D ({signal_1631, signal_984}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_381 ( .clk (clk), .D ({signal_1630, signal_985}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_383 ( .clk (clk), .D ({signal_1629, signal_986}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_385 ( .clk (clk), .D ({signal_1628, signal_987}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_387 ( .clk (clk), .D ({signal_1627, signal_988}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_389 ( .clk (clk), .D ({signal_1626, signal_989}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_391 ( .clk (clk), .D ({signal_1625, signal_990}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_393 ( .clk (clk), .D ({signal_1624, signal_991}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_395 ( .clk (clk), .D ({signal_1623, signal_992}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_397 ( .clk (clk), .D ({signal_1622, signal_993}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_399 ( .clk (clk), .D ({signal_1621, signal_994}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_401 ( .clk (clk), .D ({signal_1620, signal_995}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_403 ( .clk (clk), .D ({signal_1436, signal_996}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_405 ( .clk (clk), .D ({signal_1619, signal_997}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_407 ( .clk (clk), .D ({signal_1435, signal_998}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 cell_789 ( .CK (clk), .D (signal_2964), .Q (signal_1001), .QN () ) ;
    DFF_X1 cell_791 ( .CK (clk), .D (signal_2965), .Q (signal_1002), .QN () ) ;
    DFF_X1 cell_793 ( .CK (clk), .D (signal_2966), .Q (signal_1003), .QN () ) ;
    DFF_X1 cell_795 ( .CK (clk), .D (signal_2967), .Q (signal_1004), .QN () ) ;
    DFF_X1 cell_797 ( .CK (clk), .D (signal_2968), .Q (signal_1005), .QN () ) ;
    DFF_X1 cell_799 ( .CK (clk), .D (signal_2969), .Q (signal_1006), .QN () ) ;
    DFF_X1 cell_801 ( .CK (clk), .D (signal_2970), .Q (signal_1007), .QN () ) ;
    DFF_X1 cell_814 ( .CK (clk), .D (signal_2971), .Q (signal_1015), .QN () ) ;
    DFF_X1 cell_816 ( .CK (clk), .D (signal_2972), .Q (signal_1016), .QN () ) ;
    DFF_X1 cell_818 ( .CK (clk), .D (signal_2973), .Q (done), .QN () ) ;
endmodule
