/* modified netlist. Source: module CRAFT in file ../CaseStudies/09_CRAFT_round_based_encryption/netlists/CRAFT.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module CRAFT_LMDPL_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, Po_rst, Fresh, plaintext_s1, key_s1, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input Po_rst ;
    input [63:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [255:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire LMDPL_pre1 ;
    wire LMDPL_pre2 ;
    wire mid_rst ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;

    /* cells in depth 0 */
    mux2_masked_LMDPL InputMUX_MUXInst_0_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[0]}), .a ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, plaintext_s0[0]}), .c ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[0]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_1_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[1]}), .a ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, plaintext_s0[1]}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[1]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_2_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[2]}), .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, plaintext_s0[2]}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[2]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_3_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[3]}), .a ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, plaintext_s0[3]}), .c ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[3]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_4_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[4]}), .a ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, plaintext_s0[4]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[4]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_5_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[5]}), .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, plaintext_s0[5]}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[5]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_6_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[6]}), .a ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, plaintext_s0[6]}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[6]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_7_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[7]}), .a ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, plaintext_s0[7]}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[7]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_8_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[8]}), .a ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, plaintext_s0[8]}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[8]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_9_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[9]}), .a ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, plaintext_s0[9]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[9]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_10_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[10]}), .a ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, plaintext_s0[10]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[10]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_11_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[11]}), .a ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, plaintext_s0[11]}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[11]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_12_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[12]}), .a ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, plaintext_s0[12]}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[12]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_13_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[13]}), .a ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, plaintext_s0[13]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[13]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_14_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[14]}), .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, plaintext_s0[14]}), .c ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[14]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_15_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[15]}), .a ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, plaintext_s0[15]}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[15]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_16_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[16]}), .a ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, plaintext_s0[16]}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[16]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_17_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[17]}), .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, plaintext_s0[17]}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[17]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_18_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[18]}), .a ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, plaintext_s0[18]}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[18]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_19_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[19]}), .a ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, plaintext_s0[19]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[19]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_20_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[20]}), .a ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, plaintext_s0[20]}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[20]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_21_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[21]}), .a ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, plaintext_s0[21]}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[21]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_22_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[22]}), .a ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, plaintext_s0[22]}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[22]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_23_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[23]}), .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, plaintext_s0[23]}), .c ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[23]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_24_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[24]}), .a ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, plaintext_s0[24]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[24]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_25_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[25]}), .a ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, plaintext_s0[25]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[25]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_26_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[26]}), .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, plaintext_s0[26]}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[26]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_27_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[27]}), .a ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, plaintext_s0[27]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[27]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_28_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[28]}), .a ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, plaintext_s0[28]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[28]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_29_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[29]}), .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, plaintext_s0[29]}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCOutput[29]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_30_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[30]}), .a ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, plaintext_s0[30]}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCOutput[30]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_31_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[31]}), .a ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, plaintext_s0[31]}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCOutput[31]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_32_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[32]}), .a ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, plaintext_s0[32]}), .c ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[32]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_33_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[33]}), .a ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, plaintext_s0[33]}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[33]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_34_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[34]}), .a ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, plaintext_s0[34]}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[34]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_35_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[35]}), .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, plaintext_s0[35]}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[35]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_36_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[36]}), .a ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, plaintext_s0[36]}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[36]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_37_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[37]}), .a ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, plaintext_s0[37]}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[37]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_38_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[38]}), .a ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, plaintext_s0[38]}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[38]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_39_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[39]}), .a ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, plaintext_s0[39]}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[39]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_40_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[40]}), .a ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, plaintext_s0[40]}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[40]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_41_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[41]}), .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, plaintext_s0[41]}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[41]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_42_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[42]}), .a ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, plaintext_s0[42]}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[42]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_43_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[43]}), .a ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, plaintext_s0[43]}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[43]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_44_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[44]}), .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, plaintext_s0[44]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[44]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_45_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[45]}), .a ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, plaintext_s0[45]}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[45]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_46_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[46]}), .a ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, plaintext_s0[46]}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[46]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_47_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[47]}), .a ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, plaintext_s0[47]}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[47]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_48_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[48]}), .a ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, plaintext_s0[48]}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[48]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_49_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[49]}), .a ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, plaintext_s0[49]}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[49]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_50_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[50]}), .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, plaintext_s0[50]}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[50]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_51_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[51]}), .a ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, plaintext_s0[51]}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[51]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_52_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[52]}), .a ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, plaintext_s0[52]}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[52]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_53_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[53]}), .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, plaintext_s0[53]}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[53]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_54_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[54]}), .a ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, plaintext_s0[54]}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[54]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_55_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[55]}), .a ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, plaintext_s0[55]}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[55]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_56_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[56]}), .a ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, plaintext_s0[56]}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[56]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_57_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[57]}), .a ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, plaintext_s0[57]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[57]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_58_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[58]}), .a ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, plaintext_s0[58]}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[58]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_59_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[59]}), .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, plaintext_s0[59]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[59]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_60_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, Feedback[60]}), .a ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, plaintext_s0[60]}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[60]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_61_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, Feedback[61]}), .a ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, plaintext_s0[61]}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, MCInput[61]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_62_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, Feedback[62]}), .a ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, plaintext_s0[62]}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, MCInput[62]}) ) ;
    mux2_masked_LMDPL InputMUX_MUXInst_63_U1 ( .s ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, rst}), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[63]}), .a ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, plaintext_s0[63]}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, MCInput[63]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[48]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[16]}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[0]}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, MCInst_XOR_r0_Inst_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, MCInput[48]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, MCInst_XOR_r0_Inst_0_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[0]}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[32]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, MCInput[32]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, MCInst_XOR_r1_Inst_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[49]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[17]}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[1]}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, MCInst_XOR_r0_Inst_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, MCInput[49]}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, MCInst_XOR_r0_Inst_1_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[1]}), .c ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[33]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, MCInput[33]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, MCInst_XOR_r1_Inst_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[50]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[18]}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[2]}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, MCInst_XOR_r0_Inst_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, MCInput[50]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, MCInst_XOR_r0_Inst_2_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[2]}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[34]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, MCInput[34]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, MCInst_XOR_r1_Inst_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[51]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[19]}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[3]}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, MCInst_XOR_r0_Inst_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, MCInput[51]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, MCInst_XOR_r0_Inst_3_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[3]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[35]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, MCInput[35]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, MCInst_XOR_r1_Inst_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[52]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[20]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[4]}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, MCInst_XOR_r0_Inst_4_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_4_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, MCInput[52]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, MCInst_XOR_r0_Inst_4_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[4]}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[36]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_4_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, MCInput[36]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, MCInst_XOR_r1_Inst_4_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[53]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[21]}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[5]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, MCInst_XOR_r0_Inst_5_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_5_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, MCInput[53]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, MCInst_XOR_r0_Inst_5_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[5]}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[37]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_5_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, MCInput[37]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, MCInst_XOR_r1_Inst_5_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[54]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[22]}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[6]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, MCInst_XOR_r0_Inst_6_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_6_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, MCInput[54]}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, MCInst_XOR_r0_Inst_6_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[6]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[38]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_6_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, MCInput[38]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, MCInst_XOR_r1_Inst_6_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[55]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[23]}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[7]}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, MCInst_XOR_r0_Inst_7_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_7_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, MCInput[55]}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, MCInst_XOR_r0_Inst_7_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[7]}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[39]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_7_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, MCInput[39]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, MCInst_XOR_r1_Inst_7_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[56]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[24]}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[8]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, MCInst_XOR_r0_Inst_8_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_8_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, MCInput[56]}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, MCInst_XOR_r0_Inst_8_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[8]}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[40]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_8_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, MCInput[40]}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, MCInst_XOR_r1_Inst_8_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[57]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[25]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[9]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, MCInst_XOR_r0_Inst_9_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_9_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, MCInput[57]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, MCInst_XOR_r0_Inst_9_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[9]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[41]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_9_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, MCInput[41]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, MCInst_XOR_r1_Inst_9_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[58]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[26]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[10]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, MCInst_XOR_r0_Inst_10_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_10_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, MCInput[58]}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, MCInst_XOR_r0_Inst_10_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[10]}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[42]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_10_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, MCInput[42]}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, MCInst_XOR_r1_Inst_10_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[59]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[27]}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[11]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, MCInst_XOR_r0_Inst_11_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_11_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, MCInput[59]}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, MCInst_XOR_r0_Inst_11_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[11]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[43]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_11_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, MCInput[43]}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, MCInst_XOR_r1_Inst_11_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[60]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[28]}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[12]}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, MCInst_XOR_r0_Inst_12_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_12_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, MCInput[60]}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, MCInst_XOR_r0_Inst_12_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[12]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[44]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_12_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, MCInput[44]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, MCInst_XOR_r1_Inst_12_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, MCOutput[61]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCOutput[29]}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[13]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, MCInst_XOR_r0_Inst_13_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_13_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, MCInput[61]}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, MCInst_XOR_r0_Inst_13_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[13]}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, MCOutput[45]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_13_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, MCInput[45]}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, MCInst_XOR_r1_Inst_13_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, MCOutput[62]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCOutput[30]}), .b ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[14]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, MCInst_XOR_r0_Inst_14_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_14_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, MCInput[62]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, MCInst_XOR_r0_Inst_14_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[14]}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, MCOutput[46]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_14_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, MCInput[46]}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, MCInst_XOR_r1_Inst_14_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, MCOutput[63]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCOutput[31]}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[15]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, MCInst_XOR_r0_Inst_15_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MCInst_XOR_r0_Inst_15_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, MCInput[63]}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, MCInst_XOR_r0_Inst_15_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[15]}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, MCOutput[47]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MCInst_XOR_r1_Inst_15_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, MCInput[47]}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, MCInst_XOR_r1_Inst_15_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, SelectedKey[48]}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[48]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, MCOutput[48]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, SelectedKey[49]}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, AddRoundKeyOutput[49]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, MCOutput[49]}), .c ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, SelectedKey[50]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[50]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, MCOutput[50]}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, SelectedKey[51]}), .c ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, AddRoundKeyOutput[51]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, MCOutput[51]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, SelectedKey[52]}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[52]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, MCOutput[52]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SelectedKey[53]}), .c ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, AddRoundKeyOutput[53]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, MCOutput[53]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SelectedKey[54]}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[54]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, MCOutput[54]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, SelectedKey[55]}), .c ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, AddRoundKeyOutput[55]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, MCOutput[55]}), .c ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SelectedKey[56]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[56]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, MCOutput[56]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, SelectedKey[57]}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, AddRoundKeyOutput[57]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, MCOutput[57]}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, SelectedKey[58]}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[58]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, MCOutput[58]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SelectedKey[59]}), .c ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, AddRoundKeyOutput[59]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, MCOutput[59]}), .c ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, SelectedKey[60]}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[60]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, MCOutput[60]}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, SelectedKey[61]}), .c ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, AddRoundKeyOutput[61]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, MCOutput[61]}), .c ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SelectedKey[62]}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[62]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, MCOutput[62]}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, SelectedKey[63]}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, AddRoundKeyOutput[63]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, MCOutput[63]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, AddKeyConstXOR_XORInst_0_0_n1}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[40]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, SelectedKey[40]}), .b ({LMDPL_pre1, 1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, MCOutput[40]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, AddKeyConstXOR_XORInst_0_1_n1}), .c ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, AddRoundKeyOutput[41]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, SelectedKey[41]}), .b ({LMDPL_pre1, 1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, MCOutput[41]}), .c ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, AddKeyConstXOR_XORInst_0_2_n1}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[42]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, SelectedKey[42]}), .b ({LMDPL_pre1, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, MCOutput[42]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, AddKeyConstXOR_XORInst_0_3_n1}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, AddRoundKeyOutput[43]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, SelectedKey[43]}), .b ({LMDPL_pre1, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, MCOutput[43]}), .c ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, AddKeyConstXOR_XORInst_1_0_n1}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[44]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, SelectedKey[44]}), .b ({LMDPL_pre1, 1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, MCOutput[44]}), .c ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, AddKeyConstXOR_XORInst_1_1_n1}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, AddRoundKeyOutput[45]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, SelectedKey[45]}), .b ({LMDPL_pre1, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, MCOutput[45]}), .c ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, AddKeyConstXOR_XORInst_1_2_n1}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[46]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, SelectedKey[46]}), .b ({LMDPL_pre1, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, MCOutput[46]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, AddKeyConstXOR_XORInst_1_3_n1}), .c ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, AddRoundKeyOutput[47]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, SelectedKey[47]}), .b ({LMDPL_pre1, 1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, MCOutput[47]}), .c ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SelectedKey[0]}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[0]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, MCOutput[0]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, SelectedKey[1]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, AddRoundKeyOutput[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, MCOutput[1]}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SelectedKey[2]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[2]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, MCOutput[2]}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, SelectedKey[3]}), .c ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, AddRoundKeyOutput[3]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, MCOutput[3]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, SelectedKey[4]}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[4]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, MCOutput[4]}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, SelectedKey[5]}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, AddRoundKeyOutput[5]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, MCOutput[5]}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, SelectedKey[6]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[6]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, MCOutput[6]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, SelectedKey[7]}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, AddRoundKeyOutput[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, MCOutput[7]}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, SelectedKey[8]}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[8]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, MCOutput[8]}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, SelectedKey[9]}), .c ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, AddRoundKeyOutput[9]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, MCOutput[9]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, SelectedKey[10]}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[10]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, MCOutput[10]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, SelectedKey[11]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, AddRoundKeyOutput[11]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, MCOutput[11]}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, SelectedKey[12]}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[12]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, MCOutput[12]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, SelectedKey[13]}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, AddRoundKeyOutput[13]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, MCOutput[13]}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, SelectedKey[14]}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[14]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, MCOutput[14]}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, SelectedKey[15]}), .c ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, AddRoundKeyOutput[15]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, MCOutput[15]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, SelectedKey[16]}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[16]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, MCOutput[16]}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, SelectedKey[17]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, AddRoundKeyOutput[17]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, MCOutput[17]}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, SelectedKey[18]}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[18]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, MCOutput[18]}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, SelectedKey[19]}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, AddRoundKeyOutput[19]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, MCOutput[19]}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, SelectedKey[20]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[20]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, MCOutput[20]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, SelectedKey[21]}), .c ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, AddRoundKeyOutput[21]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, MCOutput[21]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SelectedKey[22]}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[22]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, MCOutput[22]}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SelectedKey[23]}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, AddRoundKeyOutput[23]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, MCOutput[23]}), .c ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SelectedKey[24]}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[24]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, MCOutput[24]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SelectedKey[25]}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, AddRoundKeyOutput[25]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, MCOutput[25]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SelectedKey[26]}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddRoundKeyOutput[26]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, MCOutput[26]}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SelectedKey[27]}), .c ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddRoundKeyOutput[27]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, MCOutput[27]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, SelectedKey[28]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddRoundKeyOutput[28]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, MCOutput[28]}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, SelectedKey[29]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddRoundKeyOutput[29]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, MCOutput[29]}), .c ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, SelectedKey[30]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddRoundKeyOutput[30]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, MCOutput[30]}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, SelectedKey[31]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddRoundKeyOutput[31]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, MCOutput[31]}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, SelectedKey[32]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[32]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, MCOutput[32]}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SelectedKey[33]}), .c ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, AddRoundKeyOutput[33]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, MCOutput[33]}), .c ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, SelectedKey[34]}), .c ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, AddRoundKeyOutput[34]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, MCOutput[34]}), .c ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, SelectedKey[35]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, AddRoundKeyOutput[35]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, MCOutput[35]}), .c ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SelectedKey[36]}), .c ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, AddRoundKeyOutput[36]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, MCOutput[36]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, SelectedKey[37]}), .c ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, AddRoundKeyOutput[37]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, MCOutput[37]}), .c ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, SelectedKey[38]}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, AddRoundKeyOutput[38]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, MCOutput[38]}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SelectedKey[39]}), .c ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, AddRoundKeyOutput[39]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({LMDPL_pre1, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, MCOutput[39]}), .c ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, Feedback[3]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_1570, ciphertext_s1[61], ciphertext_s0[61]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_0_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, SubCellInst_SboxInst_0_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, Feedback[2]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n11}), .b ({new_AGEMA_signal_1570, ciphertext_s1[61], ciphertext_s0[61]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, SubCellInst_SboxInst_0_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, SubCellInst_SboxInst_0_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U14 ( .a ({new_AGEMA_signal_1024, ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1026, ciphertext_s1[63], ciphertext_s0[63]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, SubCellInst_SboxInst_0_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_0_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n6}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_0_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, Feedback[1]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U11 ( .a ({new_AGEMA_signal_1024, ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SubCellInst_SboxInst_0_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U10 ( .a ({new_AGEMA_signal_1026, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SubCellInst_SboxInst_0_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_0_U9 ( .a ({new_AGEMA_signal_1030, ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SubCellInst_SboxInst_0_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, SubCellInst_SboxInst_0_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_0_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, Feedback[0]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_0_U7 ( .a ({new_AGEMA_signal_1570, ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_0_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_0_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n7}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_0_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_0_U5 ( .a ({new_AGEMA_signal_1030, ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1026, ciphertext_s1[63], ciphertext_s0[63]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_0_U4 ( .x ({new_AGEMA_signal_1024, ciphertext_s1[60], ciphertext_s0[60]}), .y ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SubCellInst_SboxInst_0_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SubCellInst_SboxInst_0_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_0_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_0_U2 ( .x ({new_AGEMA_signal_1026, ciphertext_s1[63], ciphertext_s0[63]}), .y ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SubCellInst_SboxInst_0_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_0_U1 ( .x ({new_AGEMA_signal_1030, ciphertext_s1[62], ciphertext_s0[62]}), .y ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, Feedback[7]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_1580, ciphertext_s1[49], ciphertext_s0[49]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SubCellInst_SboxInst_1_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, SubCellInst_SboxInst_1_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, Feedback[6]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n11}), .b ({new_AGEMA_signal_1580, ciphertext_s1[49], ciphertext_s0[49]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, SubCellInst_SboxInst_1_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SubCellInst_SboxInst_1_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SubCellInst_SboxInst_1_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U14 ( .a ({new_AGEMA_signal_1040, ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1042, ciphertext_s1[51], ciphertext_s0[51]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SubCellInst_SboxInst_1_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_1_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n6}), .b ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_1_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, Feedback[5]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U11 ( .a ({new_AGEMA_signal_1040, ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SubCellInst_SboxInst_1_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U10 ( .a ({new_AGEMA_signal_1042, ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SubCellInst_SboxInst_1_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_1_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_1_U9 ( .a ({new_AGEMA_signal_1046, ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SubCellInst_SboxInst_1_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_1_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, Feedback[4]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_1_U7 ( .a ({new_AGEMA_signal_1580, ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SubCellInst_SboxInst_1_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n7}), .b ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_1_U5 ( .a ({new_AGEMA_signal_1046, ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1042, ciphertext_s1[51], ciphertext_s0[51]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, SubCellInst_SboxInst_1_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_1_U4 ( .x ({new_AGEMA_signal_1040, ciphertext_s1[48], ciphertext_s0[48]}), .y ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SubCellInst_SboxInst_1_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_1_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_1_U2 ( .x ({new_AGEMA_signal_1042, ciphertext_s1[51], ciphertext_s0[51]}), .y ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SubCellInst_SboxInst_1_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_1_U1 ( .x ({new_AGEMA_signal_1046, ciphertext_s1[50], ciphertext_s0[50]}), .y ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SubCellInst_SboxInst_1_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, Feedback[11]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_1590, ciphertext_s1[53], ciphertext_s0[53]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SubCellInst_SboxInst_2_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, SubCellInst_SboxInst_2_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, Feedback[10]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n11}), .b ({new_AGEMA_signal_1590, ciphertext_s1[53], ciphertext_s0[53]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, SubCellInst_SboxInst_2_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SubCellInst_SboxInst_2_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U14 ( .a ({new_AGEMA_signal_1056, ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1058, ciphertext_s1[55], ciphertext_s0[55]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, SubCellInst_SboxInst_2_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n6}), .b ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_2_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, Feedback[9]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U11 ( .a ({new_AGEMA_signal_1056, ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_2_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U10 ( .a ({new_AGEMA_signal_1058, ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SubCellInst_SboxInst_2_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, SubCellInst_SboxInst_2_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_2_U9 ( .a ({new_AGEMA_signal_1062, ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, SubCellInst_SboxInst_2_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SubCellInst_SboxInst_2_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_2_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, Feedback[8]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_2_U7 ( .a ({new_AGEMA_signal_1590, ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_2_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SubCellInst_SboxInst_2_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n7}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_2_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_2_U5 ( .a ({new_AGEMA_signal_1062, ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1058, ciphertext_s1[55], ciphertext_s0[55]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SubCellInst_SboxInst_2_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_2_U4 ( .x ({new_AGEMA_signal_1056, ciphertext_s1[52], ciphertext_s0[52]}), .y ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, SubCellInst_SboxInst_2_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, SubCellInst_SboxInst_2_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_2_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_2_U2 ( .x ({new_AGEMA_signal_1058, ciphertext_s1[55], ciphertext_s0[55]}), .y ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, SubCellInst_SboxInst_2_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_2_U1 ( .x ({new_AGEMA_signal_1062, ciphertext_s1[54], ciphertext_s0[54]}), .y ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SubCellInst_SboxInst_2_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, Feedback[15]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_1600, ciphertext_s1[57], ciphertext_s0[57]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_3_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, SubCellInst_SboxInst_3_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, Feedback[14]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n11}), .b ({new_AGEMA_signal_1600, ciphertext_s1[57], ciphertext_s0[57]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, SubCellInst_SboxInst_3_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_3_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SubCellInst_SboxInst_3_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U14 ( .a ({new_AGEMA_signal_1072, ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1074, ciphertext_s1[59], ciphertext_s0[59]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SubCellInst_SboxInst_3_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_3_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n6}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_3_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, Feedback[13]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U11 ( .a ({new_AGEMA_signal_1072, ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SubCellInst_SboxInst_3_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U10 ( .a ({new_AGEMA_signal_1074, ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_3_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_3_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_3_U9 ( .a ({new_AGEMA_signal_1078, ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SubCellInst_SboxInst_3_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SubCellInst_SboxInst_3_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_3_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, Feedback[12]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_3_U7 ( .a ({new_AGEMA_signal_1600, ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_3_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_3_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n7}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_3_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_3_U5 ( .a ({new_AGEMA_signal_1078, ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1074, ciphertext_s1[59], ciphertext_s0[59]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_3_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_3_U4 ( .x ({new_AGEMA_signal_1072, ciphertext_s1[56], ciphertext_s0[56]}), .y ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, SubCellInst_SboxInst_3_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SubCellInst_SboxInst_3_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_3_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_3_U2 ( .x ({new_AGEMA_signal_1074, ciphertext_s1[59], ciphertext_s0[59]}), .y ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SubCellInst_SboxInst_3_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_3_U1 ( .x ({new_AGEMA_signal_1078, ciphertext_s1[58], ciphertext_s0[58]}), .y ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_3_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, Feedback[19]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_1610, ciphertext_s1[33], ciphertext_s0[33]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SubCellInst_SboxInst_4_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, SubCellInst_SboxInst_4_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, Feedback[18]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n11}), .b ({new_AGEMA_signal_1610, ciphertext_s1[33], ciphertext_s0[33]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, SubCellInst_SboxInst_4_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, SubCellInst_SboxInst_4_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SubCellInst_SboxInst_4_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U14 ( .a ({new_AGEMA_signal_1088, ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1090, ciphertext_s1[35], ciphertext_s0[35]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SubCellInst_SboxInst_4_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_4_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n6}), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_4_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, Feedback[17]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U11 ( .a ({new_AGEMA_signal_1088, ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SubCellInst_SboxInst_4_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U10 ( .a ({new_AGEMA_signal_1090, ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, SubCellInst_SboxInst_4_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SubCellInst_SboxInst_4_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_4_U9 ( .a ({new_AGEMA_signal_1094, ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, SubCellInst_SboxInst_4_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SubCellInst_SboxInst_4_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_4_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, Feedback[16]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_4_U7 ( .a ({new_AGEMA_signal_1610, ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_4_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SubCellInst_SboxInst_4_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n7}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_4_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_4_U5 ( .a ({new_AGEMA_signal_1094, ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1090, ciphertext_s1[35], ciphertext_s0[35]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SubCellInst_SboxInst_4_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_4_U4 ( .x ({new_AGEMA_signal_1088, ciphertext_s1[32], ciphertext_s0[32]}), .y ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_4_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, SubCellInst_SboxInst_4_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_4_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_4_U2 ( .x ({new_AGEMA_signal_1090, ciphertext_s1[35], ciphertext_s0[35]}), .y ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, SubCellInst_SboxInst_4_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_4_U1 ( .x ({new_AGEMA_signal_1094, ciphertext_s1[34], ciphertext_s0[34]}), .y ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, SubCellInst_SboxInst_4_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, Feedback[23]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_1620, ciphertext_s1[45], ciphertext_s0[45]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SubCellInst_SboxInst_5_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, SubCellInst_SboxInst_5_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, Feedback[22]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n11}), .b ({new_AGEMA_signal_1620, ciphertext_s1[45], ciphertext_s0[45]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, SubCellInst_SboxInst_5_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SubCellInst_SboxInst_5_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SubCellInst_SboxInst_5_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U14 ( .a ({new_AGEMA_signal_1104, ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1106, ciphertext_s1[47], ciphertext_s0[47]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, SubCellInst_SboxInst_5_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_5_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n6}), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_5_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, Feedback[21]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U11 ( .a ({new_AGEMA_signal_1104, ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_5_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U10 ( .a ({new_AGEMA_signal_1106, ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SubCellInst_SboxInst_5_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_5_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_5_U9 ( .a ({new_AGEMA_signal_1110, ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SubCellInst_SboxInst_5_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SubCellInst_SboxInst_5_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_5_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, Feedback[20]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_5_U7 ( .a ({new_AGEMA_signal_1620, ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_5_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SubCellInst_SboxInst_5_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n7}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_5_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_5_U5 ( .a ({new_AGEMA_signal_1110, ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1106, ciphertext_s1[47], ciphertext_s0[47]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SubCellInst_SboxInst_5_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_5_U4 ( .x ({new_AGEMA_signal_1104, ciphertext_s1[44], ciphertext_s0[44]}), .y ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SubCellInst_SboxInst_5_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SubCellInst_SboxInst_5_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_5_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_5_U2 ( .x ({new_AGEMA_signal_1106, ciphertext_s1[47], ciphertext_s0[47]}), .y ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SubCellInst_SboxInst_5_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_5_U1 ( .x ({new_AGEMA_signal_1110, ciphertext_s1[46], ciphertext_s0[46]}), .y ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SubCellInst_SboxInst_5_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, Feedback[27]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_1630, ciphertext_s1[41], ciphertext_s0[41]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_6_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, SubCellInst_SboxInst_6_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, Feedback[26]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n11}), .b ({new_AGEMA_signal_1630, ciphertext_s1[41], ciphertext_s0[41]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, SubCellInst_SboxInst_6_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_6_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SubCellInst_SboxInst_6_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U14 ( .a ({new_AGEMA_signal_1120, ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1122, ciphertext_s1[43], ciphertext_s0[43]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SubCellInst_SboxInst_6_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_6_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n6}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_6_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, Feedback[25]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U11 ( .a ({new_AGEMA_signal_1120, ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SubCellInst_SboxInst_6_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U10 ( .a ({new_AGEMA_signal_1122, ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_6_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SubCellInst_SboxInst_6_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_6_U9 ( .a ({new_AGEMA_signal_1126, ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SubCellInst_SboxInst_6_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SubCellInst_SboxInst_6_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_6_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, Feedback[24]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_6_U7 ( .a ({new_AGEMA_signal_1630, ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_6_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_6_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n7}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_6_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_6_U5 ( .a ({new_AGEMA_signal_1126, ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1122, ciphertext_s1[43], ciphertext_s0[43]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_6_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_6_U4 ( .x ({new_AGEMA_signal_1120, ciphertext_s1[40], ciphertext_s0[40]}), .y ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SubCellInst_SboxInst_6_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SubCellInst_SboxInst_6_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_6_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_6_U2 ( .x ({new_AGEMA_signal_1122, ciphertext_s1[43], ciphertext_s0[43]}), .y ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SubCellInst_SboxInst_6_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_6_U1 ( .x ({new_AGEMA_signal_1126, ciphertext_s1[42], ciphertext_s0[42]}), .y ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_6_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, Feedback[31]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_1640, ciphertext_s1[37], ciphertext_s0[37]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SubCellInst_SboxInst_7_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, SubCellInst_SboxInst_7_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, Feedback[30]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n11}), .b ({new_AGEMA_signal_1640, ciphertext_s1[37], ciphertext_s0[37]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, SubCellInst_SboxInst_7_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SubCellInst_SboxInst_7_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SubCellInst_SboxInst_7_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U14 ( .a ({new_AGEMA_signal_1136, ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1138, ciphertext_s1[39], ciphertext_s0[39]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, SubCellInst_SboxInst_7_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_7_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n6}), .b ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_7_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, Feedback[29]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U11 ( .a ({new_AGEMA_signal_1136, ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, SubCellInst_SboxInst_7_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U10 ( .a ({new_AGEMA_signal_1138, ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SubCellInst_SboxInst_7_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_7_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_7_U9 ( .a ({new_AGEMA_signal_1142, ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, SubCellInst_SboxInst_7_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SubCellInst_SboxInst_7_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_7_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, Feedback[28]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_7_U7 ( .a ({new_AGEMA_signal_1640, ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_7_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, SubCellInst_SboxInst_7_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n7}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_7_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_7_U5 ( .a ({new_AGEMA_signal_1142, ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1138, ciphertext_s1[39], ciphertext_s0[39]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SubCellInst_SboxInst_7_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_7_U4 ( .x ({new_AGEMA_signal_1136, ciphertext_s1[36], ciphertext_s0[36]}), .y ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_7_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, SubCellInst_SboxInst_7_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_7_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_7_U2 ( .x ({new_AGEMA_signal_1138, ciphertext_s1[39], ciphertext_s0[39]}), .y ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, SubCellInst_SboxInst_7_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_7_U1 ( .x ({new_AGEMA_signal_1142, ciphertext_s1[38], ciphertext_s0[38]}), .y ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SubCellInst_SboxInst_7_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, Feedback[35]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_1650, ciphertext_s1[17], ciphertext_s0[17]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SubCellInst_SboxInst_8_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, SubCellInst_SboxInst_8_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, Feedback[34]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n11}), .b ({new_AGEMA_signal_1650, ciphertext_s1[17], ciphertext_s0[17]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, SubCellInst_SboxInst_8_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, SubCellInst_SboxInst_8_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SubCellInst_SboxInst_8_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U14 ( .a ({new_AGEMA_signal_1152, ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1154, ciphertext_s1[19], ciphertext_s0[19]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SubCellInst_SboxInst_8_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_8_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n6}), .b ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_8_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, Feedback[33]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U11 ( .a ({new_AGEMA_signal_1152, ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_8_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U10 ( .a ({new_AGEMA_signal_1154, ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, SubCellInst_SboxInst_8_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SubCellInst_SboxInst_8_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_8_U9 ( .a ({new_AGEMA_signal_1158, ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SubCellInst_SboxInst_8_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SubCellInst_SboxInst_8_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_8_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, Feedback[32]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_8_U7 ( .a ({new_AGEMA_signal_1650, ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_8_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SubCellInst_SboxInst_8_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n7}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_8_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_8_U5 ( .a ({new_AGEMA_signal_1158, ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1154, ciphertext_s1[19], ciphertext_s0[19]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, SubCellInst_SboxInst_8_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_8_U4 ( .x ({new_AGEMA_signal_1152, ciphertext_s1[16], ciphertext_s0[16]}), .y ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, SubCellInst_SboxInst_8_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SubCellInst_SboxInst_8_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_8_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_8_U2 ( .x ({new_AGEMA_signal_1154, ciphertext_s1[19], ciphertext_s0[19]}), .y ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SubCellInst_SboxInst_8_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_8_U1 ( .x ({new_AGEMA_signal_1158, ciphertext_s1[18], ciphertext_s0[18]}), .y ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, SubCellInst_SboxInst_8_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, Feedback[39]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_1660, ciphertext_s1[29], ciphertext_s0[29]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_9_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, SubCellInst_SboxInst_9_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, Feedback[38]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n11}), .b ({new_AGEMA_signal_1660, ciphertext_s1[29], ciphertext_s0[29]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, SubCellInst_SboxInst_9_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_9_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SubCellInst_SboxInst_9_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U14 ( .a ({new_AGEMA_signal_1168, ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1170, ciphertext_s1[31], ciphertext_s0[31]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SubCellInst_SboxInst_9_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_9_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n6}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_9_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, Feedback[37]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U11 ( .a ({new_AGEMA_signal_1168, ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SubCellInst_SboxInst_9_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U10 ( .a ({new_AGEMA_signal_1170, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_9_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_9_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_9_U9 ( .a ({new_AGEMA_signal_1174, ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_9_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SubCellInst_SboxInst_9_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_9_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, Feedback[36]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_9_U7 ( .a ({new_AGEMA_signal_1660, ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_9_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_9_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n7}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_9_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_9_U5 ( .a ({new_AGEMA_signal_1174, ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1170, ciphertext_s1[31], ciphertext_s0[31]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_9_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_9_U4 ( .x ({new_AGEMA_signal_1168, ciphertext_s1[28], ciphertext_s0[28]}), .y ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SubCellInst_SboxInst_9_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_9_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_9_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_9_U2 ( .x ({new_AGEMA_signal_1170, ciphertext_s1[31], ciphertext_s0[31]}), .y ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_9_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_9_U1 ( .x ({new_AGEMA_signal_1174, ciphertext_s1[30], ciphertext_s0[30]}), .y ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_9_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, Feedback[43]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_1670, ciphertext_s1[25], ciphertext_s0[25]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, SubCellInst_SboxInst_10_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, SubCellInst_SboxInst_10_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, Feedback[42]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n11}), .b ({new_AGEMA_signal_1670, ciphertext_s1[25], ciphertext_s0[25]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, SubCellInst_SboxInst_10_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_10_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SubCellInst_SboxInst_10_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U14 ( .a ({new_AGEMA_signal_1184, ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1186, ciphertext_s1[27], ciphertext_s0[27]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, SubCellInst_SboxInst_10_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_10_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n6}), .b ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_10_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, Feedback[41]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U11 ( .a ({new_AGEMA_signal_1184, ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SubCellInst_SboxInst_10_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U10 ( .a ({new_AGEMA_signal_1186, ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_10_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_10_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_10_U9 ( .a ({new_AGEMA_signal_1190, ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SubCellInst_SboxInst_10_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SubCellInst_SboxInst_10_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_10_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, Feedback[40]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_10_U7 ( .a ({new_AGEMA_signal_1670, ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_10_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, SubCellInst_SboxInst_10_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n7}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_10_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_10_U5 ( .a ({new_AGEMA_signal_1190, ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1186, ciphertext_s1[27], ciphertext_s0[27]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_10_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_10_U4 ( .x ({new_AGEMA_signal_1184, ciphertext_s1[24], ciphertext_s0[24]}), .y ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_10_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SubCellInst_SboxInst_10_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_10_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_10_U2 ( .x ({new_AGEMA_signal_1186, ciphertext_s1[27], ciphertext_s0[27]}), .y ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SubCellInst_SboxInst_10_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_10_U1 ( .x ({new_AGEMA_signal_1190, ciphertext_s1[26], ciphertext_s0[26]}), .y ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_10_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, Feedback[47]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_1680, ciphertext_s1[21], ciphertext_s0[21]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SubCellInst_SboxInst_11_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, SubCellInst_SboxInst_11_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, Feedback[46]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n11}), .b ({new_AGEMA_signal_1680, ciphertext_s1[21], ciphertext_s0[21]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, SubCellInst_SboxInst_11_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SubCellInst_SboxInst_11_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U14 ( .a ({new_AGEMA_signal_1200, ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1202, ciphertext_s1[23], ciphertext_s0[23]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_11_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_11_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n6}), .b ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_11_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, Feedback[45]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U11 ( .a ({new_AGEMA_signal_1200, ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_11_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U10 ( .a ({new_AGEMA_signal_1202, ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_11_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_11_U9 ( .a ({new_AGEMA_signal_1206, ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SubCellInst_SboxInst_11_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SubCellInst_SboxInst_11_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_11_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, Feedback[44]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_11_U7 ( .a ({new_AGEMA_signal_1680, ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_11_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, SubCellInst_SboxInst_11_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n7}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_11_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_11_U5 ( .a ({new_AGEMA_signal_1206, ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1202, ciphertext_s1[23], ciphertext_s0[23]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, SubCellInst_SboxInst_11_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_11_U4 ( .x ({new_AGEMA_signal_1200, ciphertext_s1[20], ciphertext_s0[20]}), .y ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_11_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SubCellInst_SboxInst_11_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_11_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_11_U2 ( .x ({new_AGEMA_signal_1202, ciphertext_s1[23], ciphertext_s0[23]}), .y ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SubCellInst_SboxInst_11_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_11_U1 ( .x ({new_AGEMA_signal_1206, ciphertext_s1[22], ciphertext_s0[22]}), .y ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, Feedback[51]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_1690, ciphertext_s1[5], ciphertext_s0[5]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SubCellInst_SboxInst_12_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, SubCellInst_SboxInst_12_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, Feedback[50]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n11}), .b ({new_AGEMA_signal_1690, ciphertext_s1[5], ciphertext_s0[5]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, SubCellInst_SboxInst_12_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_12_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SubCellInst_SboxInst_12_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U14 ( .a ({new_AGEMA_signal_1216, ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1218, ciphertext_s1[7], ciphertext_s0[7]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_12_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n6}), .b ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_12_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, Feedback[49]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U11 ( .a ({new_AGEMA_signal_1216, ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, SubCellInst_SboxInst_12_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U10 ( .a ({new_AGEMA_signal_1218, ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_12_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_12_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_12_U9 ( .a ({new_AGEMA_signal_1222, ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_12_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SubCellInst_SboxInst_12_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_12_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, Feedback[48]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_12_U7 ( .a ({new_AGEMA_signal_1690, ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_12_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SubCellInst_SboxInst_12_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n7}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_12_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_12_U5 ( .a ({new_AGEMA_signal_1222, ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1218, ciphertext_s1[7], ciphertext_s0[7]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_12_U4 ( .x ({new_AGEMA_signal_1216, ciphertext_s1[4], ciphertext_s0[4]}), .y ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, SubCellInst_SboxInst_12_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_12_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_12_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_12_U2 ( .x ({new_AGEMA_signal_1218, ciphertext_s1[7], ciphertext_s0[7]}), .y ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_12_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_12_U1 ( .x ({new_AGEMA_signal_1222, ciphertext_s1[6], ciphertext_s0[6]}), .y ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_12_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, Feedback[55]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_1700, ciphertext_s1[9], ciphertext_s0[9]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, SubCellInst_SboxInst_13_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, SubCellInst_SboxInst_13_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, Feedback[54]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n11}), .b ({new_AGEMA_signal_1700, ciphertext_s1[9], ciphertext_s0[9]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, SubCellInst_SboxInst_13_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_13_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SubCellInst_SboxInst_13_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U14 ( .a ({new_AGEMA_signal_1232, ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1234, ciphertext_s1[11], ciphertext_s0[11]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SubCellInst_SboxInst_13_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_13_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n6}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_13_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, Feedback[53]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U11 ( .a ({new_AGEMA_signal_1232, ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SubCellInst_SboxInst_13_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U10 ( .a ({new_AGEMA_signal_1234, ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_13_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_13_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_13_U9 ( .a ({new_AGEMA_signal_1238, ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SubCellInst_SboxInst_13_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_13_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, Feedback[52]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_13_U7 ( .a ({new_AGEMA_signal_1700, ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_13_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SubCellInst_SboxInst_13_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n7}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_13_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_13_U5 ( .a ({new_AGEMA_signal_1238, ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1234, ciphertext_s1[11], ciphertext_s0[11]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_13_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_13_U4 ( .x ({new_AGEMA_signal_1232, ciphertext_s1[8], ciphertext_s0[8]}), .y ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_13_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_13_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_13_U2 ( .x ({new_AGEMA_signal_1234, ciphertext_s1[11], ciphertext_s0[11]}), .y ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SubCellInst_SboxInst_13_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_13_U1 ( .x ({new_AGEMA_signal_1238, ciphertext_s1[10], ciphertext_s0[10]}), .y ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_13_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, Feedback[59]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_1710, ciphertext_s1[13], ciphertext_s0[13]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, SubCellInst_SboxInst_14_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, SubCellInst_SboxInst_14_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, Feedback[58]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n11}), .b ({new_AGEMA_signal_1710, ciphertext_s1[13], ciphertext_s0[13]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, SubCellInst_SboxInst_14_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, SubCellInst_SboxInst_14_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SubCellInst_SboxInst_14_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U14 ( .a ({new_AGEMA_signal_1248, ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1250, ciphertext_s1[15], ciphertext_s0[15]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_14_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_14_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n6}), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_14_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, Feedback[57]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U11 ( .a ({new_AGEMA_signal_1248, ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SubCellInst_SboxInst_14_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U10 ( .a ({new_AGEMA_signal_1250, ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, SubCellInst_SboxInst_14_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_14_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_14_U9 ( .a ({new_AGEMA_signal_1254, ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, SubCellInst_SboxInst_14_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SubCellInst_SboxInst_14_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_14_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, Feedback[56]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_14_U7 ( .a ({new_AGEMA_signal_1710, ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_14_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, SubCellInst_SboxInst_14_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n7}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SubCellInst_SboxInst_14_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_14_U5 ( .a ({new_AGEMA_signal_1254, ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1250, ciphertext_s1[15], ciphertext_s0[15]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SubCellInst_SboxInst_14_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_14_U4 ( .x ({new_AGEMA_signal_1248, ciphertext_s1[12], ciphertext_s0[12]}), .y ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_14_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, SubCellInst_SboxInst_14_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_14_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_14_U2 ( .x ({new_AGEMA_signal_1250, ciphertext_s1[15], ciphertext_s0[15]}), .y ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, SubCellInst_SboxInst_14_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_14_U1 ( .x ({new_AGEMA_signal_1254, ciphertext_s1[14], ciphertext_s0[14]}), .y ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, SubCellInst_SboxInst_14_n9}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n14}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, Feedback[63]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b11)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_1720, ciphertext_s1[1], ciphertext_s0[1]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SubCellInst_SboxInst_15_n14}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, SubCellInst_SboxInst_15_n12}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, Feedback[62]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n11}), .b ({new_AGEMA_signal_1720, ciphertext_s1[1], ciphertext_s0[1]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, SubCellInst_SboxInst_15_n12}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_15_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SubCellInst_SboxInst_15_n11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U14 ( .a ({new_AGEMA_signal_1264, ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1266, ciphertext_s1[3], ciphertext_s0[3]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, SubCellInst_SboxInst_15_n10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n7}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SubCellInst_SboxInst_15_n15}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n6}), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, SubCellInst_SboxInst_15_n5}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, Feedback[61]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U11 ( .a ({new_AGEMA_signal_1264, ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, SubCellInst_SboxInst_15_n5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U10 ( .a ({new_AGEMA_signal_1266, ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_15_n9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_15_n4}) ) ;
    nonlinear_LMDPL #(.CONF(2'b01)) SubCellInst_SboxInst_15_U9 ( .a ({new_AGEMA_signal_1270, ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_15_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SubCellInst_SboxInst_15_n6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, SubCellInst_SboxInst_15_n3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, Feedback[60]}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_15_U7 ( .a ({new_AGEMA_signal_1720, ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, SubCellInst_SboxInst_15_n2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, SubCellInst_SboxInst_15_n3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n7}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, SubCellInst_SboxInst_15_n2}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_15_U5 ( .a ({new_AGEMA_signal_1270, ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1266, ciphertext_s1[3], ciphertext_s0[3]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_15_n1}) ) ;
    not_LMDPL SubCellInst_SboxInst_15_U4 ( .x ({new_AGEMA_signal_1264, ciphertext_s1[0], ciphertext_s0[0]}), .y ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SubCellInst_SboxInst_15_n7}) ) ;
    nonlinear_LMDPL #(.CONF(2'b10)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_15_n8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, SubCellInst_SboxInst_15_n13}) ) ;
    not_LMDPL SubCellInst_SboxInst_15_U2 ( .x ({new_AGEMA_signal_1266, ciphertext_s1[3], ciphertext_s0[3]}), .y ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_15_n8}) ) ;
    not_LMDPL SubCellInst_SboxInst_15_U1 ( .x ({new_AGEMA_signal_1270, ciphertext_s1[2], ciphertext_s0[2]}), .y ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_0_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, key_s0[64]}), .a ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, key_s0[0]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SelectedKey[0]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_1_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, key_s0[65]}), .a ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, key_s0[1]}), .c ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, SelectedKey[1]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_2_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, key_s0[66]}), .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, key_s0[2]}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SelectedKey[2]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_3_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, key_s0[67]}), .a ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, key_s0[3]}), .c ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, SelectedKey[3]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_4_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, key_s0[68]}), .a ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, key_s0[4]}), .c ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, SelectedKey[4]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_5_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, key_s0[69]}), .a ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, key_s0[5]}), .c ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, SelectedKey[5]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_6_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, key_s0[70]}), .a ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, key_s0[6]}), .c ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, SelectedKey[6]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_7_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, key_s0[71]}), .a ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, key_s0[7]}), .c ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, SelectedKey[7]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_8_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, key_s0[72]}), .a ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, key_s0[8]}), .c ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, SelectedKey[8]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_9_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, key_s0[73]}), .a ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, key_s0[9]}), .c ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, SelectedKey[9]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_10_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, key_s0[74]}), .a ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, key_s0[10]}), .c ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, SelectedKey[10]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_11_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, key_s0[75]}), .a ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, key_s0[11]}), .c ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, SelectedKey[11]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_12_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, key_s0[76]}), .a ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, key_s0[12]}), .c ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, SelectedKey[12]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_13_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1926, new_AGEMA_signal_1925, key_s0[77]}), .a ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, key_s0[13]}), .c ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, SelectedKey[13]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_14_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, key_s0[78]}), .a ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, key_s0[14]}), .c ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, SelectedKey[14]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_15_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, key_s0[79]}), .a ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, key_s0[15]}), .c ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, SelectedKey[15]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_16_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, key_s0[80]}), .a ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, key_s0[16]}), .c ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, SelectedKey[16]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_17_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, key_s0[81]}), .a ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, key_s0[17]}), .c ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, SelectedKey[17]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_18_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, key_s0[82]}), .a ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, key_s0[18]}), .c ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, SelectedKey[18]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_19_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, key_s0[83]}), .a ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, key_s0[19]}), .c ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, SelectedKey[19]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_20_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, key_s0[84]}), .a ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, key_s0[20]}), .c ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, SelectedKey[20]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_21_U1 ( .s ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, KeyMUX_n8}), .b ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, key_s0[85]}), .a ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, key_s0[21]}), .c ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, SelectedKey[21]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_22_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, key_s0[86]}), .a ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, key_s0[22]}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SelectedKey[22]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_23_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, key_s0[87]}), .a ({new_AGEMA_signal_1494, new_AGEMA_signal_1493, key_s0[23]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SelectedKey[23]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_24_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, key_s0[88]}), .a ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, key_s0[24]}), .c ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SelectedKey[24]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_25_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, key_s0[89]}), .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, key_s0[25]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SelectedKey[25]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_26_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, key_s0[90]}), .a ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, key_s0[26]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SelectedKey[26]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_27_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, key_s0[91]}), .a ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, key_s0[27]}), .c ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SelectedKey[27]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_28_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, key_s0[92]}), .a ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, key_s0[28]}), .c ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, SelectedKey[28]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_29_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, key_s0[93]}), .a ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, key_s0[29]}), .c ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, SelectedKey[29]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_30_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, key_s0[94]}), .a ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, key_s0[30]}), .c ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, SelectedKey[30]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_31_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, key_s0[95]}), .a ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, key_s0[31]}), .c ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, SelectedKey[31]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_32_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, key_s0[96]}), .a ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, key_s0[32]}), .c ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, SelectedKey[32]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_33_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, key_s0[97]}), .a ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, key_s0[33]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SelectedKey[33]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_34_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, key_s0[98]}), .a ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, key_s0[34]}), .c ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, SelectedKey[34]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_35_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, key_s0[99]}), .a ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, key_s0[35]}), .c ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, SelectedKey[35]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_36_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, key_s0[100]}), .a ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, key_s0[36]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SelectedKey[36]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_37_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, key_s0[101]}), .a ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, key_s0[37]}), .c ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, SelectedKey[37]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_38_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, key_s0[102]}), .a ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, key_s0[38]}), .c ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, SelectedKey[38]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_39_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, key_s0[103]}), .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, key_s0[39]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SelectedKey[39]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_40_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, key_s0[104]}), .a ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, key_s0[40]}), .c ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, SelectedKey[40]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_41_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, key_s0[105]}), .a ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, key_s0[41]}), .c ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, SelectedKey[41]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_42_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, key_s0[106]}), .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, key_s0[42]}), .c ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, SelectedKey[42]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_43_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, key_s0[107]}), .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, key_s0[43]}), .c ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, SelectedKey[43]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_44_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, key_s0[108]}), .a ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, key_s0[44]}), .c ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, SelectedKey[44]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_45_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, key_s0[109]}), .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, key_s0[45]}), .c ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, SelectedKey[45]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_46_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, key_s0[110]}), .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, key_s0[46]}), .c ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, SelectedKey[46]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_47_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, key_s0[111]}), .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, key_s0[47]}), .c ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, SelectedKey[47]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_48_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, key_s0[112]}), .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, key_s0[48]}), .c ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, SelectedKey[48]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_49_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, key_s0[113]}), .a ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, key_s0[49]}), .c ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, SelectedKey[49]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_50_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, key_s0[114]}), .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, key_s0[50]}), .c ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, SelectedKey[50]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_51_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, key_s0[115]}), .a ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, key_s0[51]}), .c ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, SelectedKey[51]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_52_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, key_s0[116]}), .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, key_s0[52]}), .c ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, SelectedKey[52]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_53_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, key_s0[117]}), .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, key_s0[53]}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SelectedKey[53]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_54_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, key_s0[118]}), .a ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, key_s0[54]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SelectedKey[54]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_55_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, key_s0[119]}), .a ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, key_s0[55]}), .c ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, SelectedKey[55]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_56_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, key_s0[120]}), .a ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, key_s0[56]}), .c ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SelectedKey[56]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_57_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, key_s0[121]}), .a ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, key_s0[57]}), .c ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, SelectedKey[57]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_58_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, key_s0[122]}), .a ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, key_s0[58]}), .c ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, SelectedKey[58]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_59_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, key_s0[123]}), .a ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, key_s0[59]}), .c ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SelectedKey[59]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_60_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, key_s0[124]}), .a ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, key_s0[60]}), .c ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, SelectedKey[60]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_61_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, key_s0[125]}), .a ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, key_s0[61]}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, SelectedKey[61]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_62_U1 ( .s ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, selects[0]}), .b ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, key_s0[126]}), .a ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, key_s0[62]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SelectedKey[62]}) ) ;
    mux2_masked_LMDPL KeyMUX_MUXInst_63_U1 ( .s ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, KeyMUX_n7}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, key_s0[127]}), .a ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, key_s0[63]}), .c ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;
    Precharger_reg new_AGEMA_gate_819 ( .D (selects[0]), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1472, new_AGEMA_signal_1471}) ) ;
    Precharger_reg new_AGEMA_gate_820 ( .D (KeyMUX_n8), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1858, new_AGEMA_signal_1857}) ) ;
    Precharger_reg new_AGEMA_gate_821 ( .D (KeyMUX_n7), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_1980, new_AGEMA_signal_1979}) ) ;
    Precharger_reg new_AGEMA_gate_822 ( .D (rst), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2150, new_AGEMA_signal_2149}) ) ;
    ClockController_LMDPL ClockControllerInst ( .clk (clk), .Po_rst (Po_rst), .pre1 (LMDPL_pre1), .pre2 (LMDPL_pre2), .mid_rst (mid_rst) ) ;
    Precharger PrechargeCell_0 ( .D (plaintext_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2404, new_AGEMA_signal_2403}) ) ;
    Precharger PrechargeCell_1 ( .D (plaintext_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2400, new_AGEMA_signal_2399}) ) ;
    Precharger PrechargeCell_2 ( .D (plaintext_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2396, new_AGEMA_signal_2395}) ) ;
    Precharger PrechargeCell_3 ( .D (plaintext_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2392, new_AGEMA_signal_2391}) ) ;
    Precharger PrechargeCell_4 ( .D (plaintext_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2388, new_AGEMA_signal_2387}) ) ;
    Precharger PrechargeCell_5 ( .D (plaintext_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2384, new_AGEMA_signal_2383}) ) ;
    Precharger PrechargeCell_6 ( .D (plaintext_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2380, new_AGEMA_signal_2379}) ) ;
    Precharger PrechargeCell_7 ( .D (plaintext_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2376, new_AGEMA_signal_2375}) ) ;
    Precharger PrechargeCell_8 ( .D (plaintext_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2372, new_AGEMA_signal_2371}) ) ;
    Precharger PrechargeCell_9 ( .D (plaintext_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2368, new_AGEMA_signal_2367}) ) ;
    Precharger PrechargeCell_10 ( .D (plaintext_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2364, new_AGEMA_signal_2363}) ) ;
    Precharger PrechargeCell_11 ( .D (plaintext_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2360, new_AGEMA_signal_2359}) ) ;
    Precharger PrechargeCell_12 ( .D (plaintext_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2356, new_AGEMA_signal_2355}) ) ;
    Precharger PrechargeCell_13 ( .D (plaintext_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2352, new_AGEMA_signal_2351}) ) ;
    Precharger PrechargeCell_14 ( .D (plaintext_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2348, new_AGEMA_signal_2347}) ) ;
    Precharger PrechargeCell_15 ( .D (plaintext_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2344, new_AGEMA_signal_2343}) ) ;
    Precharger PrechargeCell_16 ( .D (plaintext_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2340, new_AGEMA_signal_2339}) ) ;
    Precharger PrechargeCell_17 ( .D (plaintext_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2336, new_AGEMA_signal_2335}) ) ;
    Precharger PrechargeCell_18 ( .D (plaintext_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2332, new_AGEMA_signal_2331}) ) ;
    Precharger PrechargeCell_19 ( .D (plaintext_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2328, new_AGEMA_signal_2327}) ) ;
    Precharger PrechargeCell_20 ( .D (plaintext_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2324, new_AGEMA_signal_2323}) ) ;
    Precharger PrechargeCell_21 ( .D (plaintext_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2320, new_AGEMA_signal_2319}) ) ;
    Precharger PrechargeCell_22 ( .D (plaintext_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2316, new_AGEMA_signal_2315}) ) ;
    Precharger PrechargeCell_23 ( .D (plaintext_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2312, new_AGEMA_signal_2311}) ) ;
    Precharger PrechargeCell_24 ( .D (plaintext_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2308, new_AGEMA_signal_2307}) ) ;
    Precharger PrechargeCell_25 ( .D (plaintext_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2304, new_AGEMA_signal_2303}) ) ;
    Precharger PrechargeCell_26 ( .D (plaintext_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2300, new_AGEMA_signal_2299}) ) ;
    Precharger PrechargeCell_27 ( .D (plaintext_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2296, new_AGEMA_signal_2295}) ) ;
    Precharger PrechargeCell_28 ( .D (plaintext_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2292, new_AGEMA_signal_2291}) ) ;
    Precharger PrechargeCell_29 ( .D (plaintext_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2288, new_AGEMA_signal_2287}) ) ;
    Precharger PrechargeCell_30 ( .D (plaintext_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2284, new_AGEMA_signal_2283}) ) ;
    Precharger PrechargeCell_31 ( .D (plaintext_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2280, new_AGEMA_signal_2279}) ) ;
    Precharger PrechargeCell_32 ( .D (plaintext_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2276, new_AGEMA_signal_2275}) ) ;
    Precharger PrechargeCell_33 ( .D (plaintext_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2272, new_AGEMA_signal_2271}) ) ;
    Precharger PrechargeCell_34 ( .D (plaintext_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2268, new_AGEMA_signal_2267}) ) ;
    Precharger PrechargeCell_35 ( .D (plaintext_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2264, new_AGEMA_signal_2263}) ) ;
    Precharger PrechargeCell_36 ( .D (plaintext_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2260, new_AGEMA_signal_2259}) ) ;
    Precharger PrechargeCell_37 ( .D (plaintext_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2256, new_AGEMA_signal_2255}) ) ;
    Precharger PrechargeCell_38 ( .D (plaintext_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2252, new_AGEMA_signal_2251}) ) ;
    Precharger PrechargeCell_39 ( .D (plaintext_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2248, new_AGEMA_signal_2247}) ) ;
    Precharger PrechargeCell_40 ( .D (plaintext_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2244, new_AGEMA_signal_2243}) ) ;
    Precharger PrechargeCell_41 ( .D (plaintext_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2240, new_AGEMA_signal_2239}) ) ;
    Precharger PrechargeCell_42 ( .D (plaintext_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2236, new_AGEMA_signal_2235}) ) ;
    Precharger PrechargeCell_43 ( .D (plaintext_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2232, new_AGEMA_signal_2231}) ) ;
    Precharger PrechargeCell_44 ( .D (plaintext_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2228, new_AGEMA_signal_2227}) ) ;
    Precharger PrechargeCell_45 ( .D (plaintext_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2224, new_AGEMA_signal_2223}) ) ;
    Precharger PrechargeCell_46 ( .D (plaintext_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2220, new_AGEMA_signal_2219}) ) ;
    Precharger PrechargeCell_47 ( .D (plaintext_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2216, new_AGEMA_signal_2215}) ) ;
    Precharger PrechargeCell_48 ( .D (plaintext_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2212, new_AGEMA_signal_2211}) ) ;
    Precharger PrechargeCell_49 ( .D (plaintext_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2208, new_AGEMA_signal_2207}) ) ;
    Precharger PrechargeCell_50 ( .D (plaintext_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2204, new_AGEMA_signal_2203}) ) ;
    Precharger PrechargeCell_51 ( .D (plaintext_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2200, new_AGEMA_signal_2199}) ) ;
    Precharger PrechargeCell_52 ( .D (plaintext_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2196, new_AGEMA_signal_2195}) ) ;
    Precharger PrechargeCell_53 ( .D (plaintext_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2192, new_AGEMA_signal_2191}) ) ;
    Precharger PrechargeCell_54 ( .D (plaintext_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2188, new_AGEMA_signal_2187}) ) ;
    Precharger PrechargeCell_55 ( .D (plaintext_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2184, new_AGEMA_signal_2183}) ) ;
    Precharger PrechargeCell_56 ( .D (plaintext_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2180, new_AGEMA_signal_2179}) ) ;
    Precharger PrechargeCell_57 ( .D (plaintext_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2176, new_AGEMA_signal_2175}) ) ;
    Precharger PrechargeCell_58 ( .D (plaintext_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2172, new_AGEMA_signal_2171}) ) ;
    Precharger PrechargeCell_59 ( .D (plaintext_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2168, new_AGEMA_signal_2167}) ) ;
    Precharger PrechargeCell_60 ( .D (plaintext_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2164, new_AGEMA_signal_2163}) ) ;
    Precharger PrechargeCell_61 ( .D (plaintext_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2160, new_AGEMA_signal_2159}) ) ;
    Precharger PrechargeCell_62 ( .D (plaintext_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2156, new_AGEMA_signal_2155}) ) ;
    Precharger PrechargeCell_63 ( .D (plaintext_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2152, new_AGEMA_signal_2151}) ) ;
    Precharger PrechargeCell_64 ( .D (key_s1[127]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2144, new_AGEMA_signal_2143}) ) ;
    Precharger PrechargeCell_65 ( .D (key_s1[126]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1564, new_AGEMA_signal_1563}) ) ;
    Precharger PrechargeCell_66 ( .D (key_s1[125]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2138, new_AGEMA_signal_2137}) ) ;
    Precharger PrechargeCell_67 ( .D (key_s1[124]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2132, new_AGEMA_signal_2131}) ) ;
    Precharger PrechargeCell_68 ( .D (key_s1[123]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1558, new_AGEMA_signal_1557}) ) ;
    Precharger PrechargeCell_69 ( .D (key_s1[122]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2126, new_AGEMA_signal_2125}) ) ;
    Precharger PrechargeCell_70 ( .D (key_s1[121]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2120, new_AGEMA_signal_2119}) ) ;
    Precharger PrechargeCell_71 ( .D (key_s1[120]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1552, new_AGEMA_signal_1551}) ) ;
    Precharger PrechargeCell_72 ( .D (key_s1[119]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2114, new_AGEMA_signal_2113}) ) ;
    Precharger PrechargeCell_73 ( .D (key_s1[118]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1546, new_AGEMA_signal_1545}) ) ;
    Precharger PrechargeCell_74 ( .D (key_s1[117]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1540, new_AGEMA_signal_1539}) ) ;
    Precharger PrechargeCell_75 ( .D (key_s1[116]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2108, new_AGEMA_signal_2107}) ) ;
    Precharger PrechargeCell_76 ( .D (key_s1[115]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2102, new_AGEMA_signal_2101}) ) ;
    Precharger PrechargeCell_77 ( .D (key_s1[114]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2096, new_AGEMA_signal_2095}) ) ;
    Precharger PrechargeCell_78 ( .D (key_s1[113]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2090, new_AGEMA_signal_2089}) ) ;
    Precharger PrechargeCell_79 ( .D (key_s1[112]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2084, new_AGEMA_signal_2083}) ) ;
    Precharger PrechargeCell_80 ( .D (key_s1[111]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2078, new_AGEMA_signal_2077}) ) ;
    Precharger PrechargeCell_81 ( .D (key_s1[110]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2072, new_AGEMA_signal_2071}) ) ;
    Precharger PrechargeCell_82 ( .D (key_s1[109]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2066, new_AGEMA_signal_2065}) ) ;
    Precharger PrechargeCell_83 ( .D (key_s1[108]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2060, new_AGEMA_signal_2059}) ) ;
    Precharger PrechargeCell_84 ( .D (key_s1[107]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2054, new_AGEMA_signal_2053}) ) ;
    Precharger PrechargeCell_85 ( .D (key_s1[106]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2048, new_AGEMA_signal_2047}) ) ;
    Precharger PrechargeCell_86 ( .D (key_s1[105]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2042, new_AGEMA_signal_2041}) ) ;
    Precharger PrechargeCell_87 ( .D (key_s1[104]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2036, new_AGEMA_signal_2035}) ) ;
    Precharger PrechargeCell_88 ( .D (key_s1[103]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1534, new_AGEMA_signal_1533}) ) ;
    Precharger PrechargeCell_89 ( .D (key_s1[102]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2030, new_AGEMA_signal_2029}) ) ;
    Precharger PrechargeCell_90 ( .D (key_s1[101]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2024, new_AGEMA_signal_2023}) ) ;
    Precharger PrechargeCell_91 ( .D (key_s1[100]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1528, new_AGEMA_signal_1527}) ) ;
    Precharger PrechargeCell_92 ( .D (key_s1[99]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2018, new_AGEMA_signal_2017}) ) ;
    Precharger PrechargeCell_93 ( .D (key_s1[98]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2012, new_AGEMA_signal_2011}) ) ;
    Precharger PrechargeCell_94 ( .D (key_s1[97]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1522, new_AGEMA_signal_1521}) ) ;
    Precharger PrechargeCell_95 ( .D (key_s1[96]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2006, new_AGEMA_signal_2005}) ) ;
    Precharger PrechargeCell_96 ( .D (key_s1[95]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2000, new_AGEMA_signal_1999}) ) ;
    Precharger PrechargeCell_97 ( .D (key_s1[94]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1994, new_AGEMA_signal_1993}) ) ;
    Precharger PrechargeCell_98 ( .D (key_s1[93]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1988, new_AGEMA_signal_1987}) ) ;
    Precharger PrechargeCell_99 ( .D (key_s1[92]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1982, new_AGEMA_signal_1981}) ) ;
    Precharger PrechargeCell_100 ( .D (key_s1[91]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1516, new_AGEMA_signal_1515}) ) ;
    Precharger PrechargeCell_101 ( .D (key_s1[90]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1510, new_AGEMA_signal_1509}) ) ;
    Precharger PrechargeCell_102 ( .D (key_s1[89]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1504, new_AGEMA_signal_1503}) ) ;
    Precharger PrechargeCell_103 ( .D (key_s1[88]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1498, new_AGEMA_signal_1497}) ) ;
    Precharger PrechargeCell_104 ( .D (key_s1[87]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1492, new_AGEMA_signal_1491}) ) ;
    Precharger PrechargeCell_105 ( .D (key_s1[86]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1486, new_AGEMA_signal_1485}) ) ;
    Precharger PrechargeCell_106 ( .D (key_s1[85]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1974, new_AGEMA_signal_1973}) ) ;
    Precharger PrechargeCell_107 ( .D (key_s1[84]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1968, new_AGEMA_signal_1967}) ) ;
    Precharger PrechargeCell_108 ( .D (key_s1[83]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1962, new_AGEMA_signal_1961}) ) ;
    Precharger PrechargeCell_109 ( .D (key_s1[82]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1956, new_AGEMA_signal_1955}) ) ;
    Precharger PrechargeCell_110 ( .D (key_s1[81]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1950, new_AGEMA_signal_1949}) ) ;
    Precharger PrechargeCell_111 ( .D (key_s1[80]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1944, new_AGEMA_signal_1943}) ) ;
    Precharger PrechargeCell_112 ( .D (key_s1[79]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1938, new_AGEMA_signal_1937}) ) ;
    Precharger PrechargeCell_113 ( .D (key_s1[78]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1932, new_AGEMA_signal_1931}) ) ;
    Precharger PrechargeCell_114 ( .D (key_s1[77]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1926, new_AGEMA_signal_1925}) ) ;
    Precharger PrechargeCell_115 ( .D (key_s1[76]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1920, new_AGEMA_signal_1919}) ) ;
    Precharger PrechargeCell_116 ( .D (key_s1[75]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1914, new_AGEMA_signal_1913}) ) ;
    Precharger PrechargeCell_117 ( .D (key_s1[74]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1908, new_AGEMA_signal_1907}) ) ;
    Precharger PrechargeCell_118 ( .D (key_s1[73]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1902, new_AGEMA_signal_1901}) ) ;
    Precharger PrechargeCell_119 ( .D (key_s1[72]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1896, new_AGEMA_signal_1895}) ) ;
    Precharger PrechargeCell_120 ( .D (key_s1[71]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1890, new_AGEMA_signal_1889}) ) ;
    Precharger PrechargeCell_121 ( .D (key_s1[70]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1884, new_AGEMA_signal_1883}) ) ;
    Precharger PrechargeCell_122 ( .D (key_s1[69]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1878, new_AGEMA_signal_1877}) ) ;
    Precharger PrechargeCell_123 ( .D (key_s1[68]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1872, new_AGEMA_signal_1871}) ) ;
    Precharger PrechargeCell_124 ( .D (key_s1[67]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1866, new_AGEMA_signal_1865}) ) ;
    Precharger PrechargeCell_125 ( .D (key_s1[66]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1480, new_AGEMA_signal_1479}) ) ;
    Precharger PrechargeCell_126 ( .D (key_s1[65]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1860, new_AGEMA_signal_1859}) ) ;
    Precharger PrechargeCell_127 ( .D (key_s1[64]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1474, new_AGEMA_signal_1473}) ) ;
    Precharger PrechargeCell_128 ( .D (key_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2146, new_AGEMA_signal_2145}) ) ;
    Precharger PrechargeCell_129 ( .D (key_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1566, new_AGEMA_signal_1565}) ) ;
    Precharger PrechargeCell_130 ( .D (key_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2140, new_AGEMA_signal_2139}) ) ;
    Precharger PrechargeCell_131 ( .D (key_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2134, new_AGEMA_signal_2133}) ) ;
    Precharger PrechargeCell_132 ( .D (key_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1560, new_AGEMA_signal_1559}) ) ;
    Precharger PrechargeCell_133 ( .D (key_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2128, new_AGEMA_signal_2127}) ) ;
    Precharger PrechargeCell_134 ( .D (key_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2122, new_AGEMA_signal_2121}) ) ;
    Precharger PrechargeCell_135 ( .D (key_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1554, new_AGEMA_signal_1553}) ) ;
    Precharger PrechargeCell_136 ( .D (key_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2116, new_AGEMA_signal_2115}) ) ;
    Precharger PrechargeCell_137 ( .D (key_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1548, new_AGEMA_signal_1547}) ) ;
    Precharger PrechargeCell_138 ( .D (key_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1542, new_AGEMA_signal_1541}) ) ;
    Precharger PrechargeCell_139 ( .D (key_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2110, new_AGEMA_signal_2109}) ) ;
    Precharger PrechargeCell_140 ( .D (key_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2104, new_AGEMA_signal_2103}) ) ;
    Precharger PrechargeCell_141 ( .D (key_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2098, new_AGEMA_signal_2097}) ) ;
    Precharger PrechargeCell_142 ( .D (key_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2092, new_AGEMA_signal_2091}) ) ;
    Precharger PrechargeCell_143 ( .D (key_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2086, new_AGEMA_signal_2085}) ) ;
    Precharger PrechargeCell_144 ( .D (key_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2080, new_AGEMA_signal_2079}) ) ;
    Precharger PrechargeCell_145 ( .D (key_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2074, new_AGEMA_signal_2073}) ) ;
    Precharger PrechargeCell_146 ( .D (key_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2068, new_AGEMA_signal_2067}) ) ;
    Precharger PrechargeCell_147 ( .D (key_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2062, new_AGEMA_signal_2061}) ) ;
    Precharger PrechargeCell_148 ( .D (key_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2056, new_AGEMA_signal_2055}) ) ;
    Precharger PrechargeCell_149 ( .D (key_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2050, new_AGEMA_signal_2049}) ) ;
    Precharger PrechargeCell_150 ( .D (key_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2044, new_AGEMA_signal_2043}) ) ;
    Precharger PrechargeCell_151 ( .D (key_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2038, new_AGEMA_signal_2037}) ) ;
    Precharger PrechargeCell_152 ( .D (key_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1536, new_AGEMA_signal_1535}) ) ;
    Precharger PrechargeCell_153 ( .D (key_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2032, new_AGEMA_signal_2031}) ) ;
    Precharger PrechargeCell_154 ( .D (key_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2026, new_AGEMA_signal_2025}) ) ;
    Precharger PrechargeCell_155 ( .D (key_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1530, new_AGEMA_signal_1529}) ) ;
    Precharger PrechargeCell_156 ( .D (key_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2020, new_AGEMA_signal_2019}) ) ;
    Precharger PrechargeCell_157 ( .D (key_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2014, new_AGEMA_signal_2013}) ) ;
    Precharger PrechargeCell_158 ( .D (key_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1524, new_AGEMA_signal_1523}) ) ;
    Precharger PrechargeCell_159 ( .D (key_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2008, new_AGEMA_signal_2007}) ) ;
    Precharger PrechargeCell_160 ( .D (key_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2002, new_AGEMA_signal_2001}) ) ;
    Precharger PrechargeCell_161 ( .D (key_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1996, new_AGEMA_signal_1995}) ) ;
    Precharger PrechargeCell_162 ( .D (key_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1990, new_AGEMA_signal_1989}) ) ;
    Precharger PrechargeCell_163 ( .D (key_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1984, new_AGEMA_signal_1983}) ) ;
    Precharger PrechargeCell_164 ( .D (key_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1518, new_AGEMA_signal_1517}) ) ;
    Precharger PrechargeCell_165 ( .D (key_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1512, new_AGEMA_signal_1511}) ) ;
    Precharger PrechargeCell_166 ( .D (key_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1506, new_AGEMA_signal_1505}) ) ;
    Precharger PrechargeCell_167 ( .D (key_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1500, new_AGEMA_signal_1499}) ) ;
    Precharger PrechargeCell_168 ( .D (key_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1494, new_AGEMA_signal_1493}) ) ;
    Precharger PrechargeCell_169 ( .D (key_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1488, new_AGEMA_signal_1487}) ) ;
    Precharger PrechargeCell_170 ( .D (key_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1976, new_AGEMA_signal_1975}) ) ;
    Precharger PrechargeCell_171 ( .D (key_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1970, new_AGEMA_signal_1969}) ) ;
    Precharger PrechargeCell_172 ( .D (key_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1964, new_AGEMA_signal_1963}) ) ;
    Precharger PrechargeCell_173 ( .D (key_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1958, new_AGEMA_signal_1957}) ) ;
    Precharger PrechargeCell_174 ( .D (key_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1952, new_AGEMA_signal_1951}) ) ;
    Precharger PrechargeCell_175 ( .D (key_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1946, new_AGEMA_signal_1945}) ) ;
    Precharger PrechargeCell_176 ( .D (key_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1940, new_AGEMA_signal_1939}) ) ;
    Precharger PrechargeCell_177 ( .D (key_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1934, new_AGEMA_signal_1933}) ) ;
    Precharger PrechargeCell_178 ( .D (key_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1928, new_AGEMA_signal_1927}) ) ;
    Precharger PrechargeCell_179 ( .D (key_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1922, new_AGEMA_signal_1921}) ) ;
    Precharger PrechargeCell_180 ( .D (key_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1916, new_AGEMA_signal_1915}) ) ;
    Precharger PrechargeCell_181 ( .D (key_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1910, new_AGEMA_signal_1909}) ) ;
    Precharger PrechargeCell_182 ( .D (key_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1904, new_AGEMA_signal_1903}) ) ;
    Precharger PrechargeCell_183 ( .D (key_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1898, new_AGEMA_signal_1897}) ) ;
    Precharger PrechargeCell_184 ( .D (key_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1892, new_AGEMA_signal_1891}) ) ;
    Precharger PrechargeCell_185 ( .D (key_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1886, new_AGEMA_signal_1885}) ) ;
    Precharger PrechargeCell_186 ( .D (key_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1880, new_AGEMA_signal_1879}) ) ;
    Precharger PrechargeCell_187 ( .D (key_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1874, new_AGEMA_signal_1873}) ) ;
    Precharger PrechargeCell_188 ( .D (key_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1868, new_AGEMA_signal_1867}) ) ;
    Precharger PrechargeCell_189 ( .D (key_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1482, new_AGEMA_signal_1481}) ) ;
    Precharger PrechargeCell_190 ( .D (key_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1862, new_AGEMA_signal_1861}) ) ;
    Precharger PrechargeCell_191 ( .D (key_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_1476, new_AGEMA_signal_1475}) ) ;

    /* register cells */
    reg_LMDPL StateReg_s_current_state_reg_63__FF_FF ( .D ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, AddRoundKeyOutput[63]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1026, ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_62__FF_FF ( .D ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, AddRoundKeyOutput[62]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1030, ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_61__FF_FF ( .D ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, AddRoundKeyOutput[61]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1570, ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_60__FF_FF ( .D ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, AddRoundKeyOutput[60]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1024, ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_59__FF_FF ( .D ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, AddRoundKeyOutput[59]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1074, ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_58__FF_FF ( .D ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, AddRoundKeyOutput[58]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1078, ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_57__FF_FF ( .D ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, AddRoundKeyOutput[57]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1600, ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_56__FF_FF ( .D ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, AddRoundKeyOutput[56]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1072, ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_55__FF_FF ( .D ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, AddRoundKeyOutput[55]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1058, ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_54__FF_FF ( .D ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, AddRoundKeyOutput[54]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1062, ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_53__FF_FF ( .D ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, AddRoundKeyOutput[53]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1590, ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_52__FF_FF ( .D ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, AddRoundKeyOutput[52]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1056, ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_51__FF_FF ( .D ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, AddRoundKeyOutput[51]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1042, ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_50__FF_FF ( .D ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, AddRoundKeyOutput[50]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1046, ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_49__FF_FF ( .D ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, AddRoundKeyOutput[49]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1580, ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_48__FF_FF ( .D ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, AddRoundKeyOutput[48]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1040, ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_47__FF_FF ( .D ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, AddRoundKeyOutput[47]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1106, ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_46__FF_FF ( .D ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, AddRoundKeyOutput[46]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1110, ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_45__FF_FF ( .D ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, AddRoundKeyOutput[45]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1620, ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_44__FF_FF ( .D ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, AddRoundKeyOutput[44]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1104, ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_43__FF_FF ( .D ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, AddRoundKeyOutput[43]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1122, ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_42__FF_FF ( .D ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, AddRoundKeyOutput[42]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1126, ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_41__FF_FF ( .D ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, AddRoundKeyOutput[41]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1630, ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_40__FF_FF ( .D ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, AddRoundKeyOutput[40]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1120, ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_39__FF_FF ( .D ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, AddRoundKeyOutput[39]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1138, ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_38__FF_FF ( .D ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, AddRoundKeyOutput[38]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1142, ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_37__FF_FF ( .D ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, AddRoundKeyOutput[37]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1640, ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_36__FF_FF ( .D ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, AddRoundKeyOutput[36]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1136, ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_35__FF_FF ( .D ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, AddRoundKeyOutput[35]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1090, ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_34__FF_FF ( .D ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, AddRoundKeyOutput[34]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1094, ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_33__FF_FF ( .D ({new_AGEMA_signal_2826, new_AGEMA_signal_2825, AddRoundKeyOutput[33]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1610, ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_32__FF_FF ( .D ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, AddRoundKeyOutput[32]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1088, ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_31__FF_FF ( .D ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, AddRoundKeyOutput[31]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1170, ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_30__FF_FF ( .D ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, AddRoundKeyOutput[30]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1174, ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_29__FF_FF ( .D ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, AddRoundKeyOutput[29]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1660, ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_28__FF_FF ( .D ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, AddRoundKeyOutput[28]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1168, ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_27__FF_FF ( .D ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, AddRoundKeyOutput[27]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1186, ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_26__FF_FF ( .D ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, AddRoundKeyOutput[26]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1190, ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_25__FF_FF ( .D ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, AddRoundKeyOutput[25]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1670, ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_24__FF_FF ( .D ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, AddRoundKeyOutput[24]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1184, ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_23__FF_FF ( .D ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, AddRoundKeyOutput[23]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1202, ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_22__FF_FF ( .D ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, AddRoundKeyOutput[22]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1206, ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_21__FF_FF ( .D ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, AddRoundKeyOutput[21]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1680, ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_20__FF_FF ( .D ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, AddRoundKeyOutput[20]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1200, ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_19__FF_FF ( .D ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, AddRoundKeyOutput[19]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1154, ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_18__FF_FF ( .D ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, AddRoundKeyOutput[18]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1158, ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_17__FF_FF ( .D ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, AddRoundKeyOutput[17]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1650, ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_16__FF_FF ( .D ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, AddRoundKeyOutput[16]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1152, ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_15__FF_FF ( .D ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, AddRoundKeyOutput[15]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1250, ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_14__FF_FF ( .D ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, AddRoundKeyOutput[14]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1254, ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_13__FF_FF ( .D ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, AddRoundKeyOutput[13]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1710, ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_12__FF_FF ( .D ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, AddRoundKeyOutput[12]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1248, ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_11__FF_FF ( .D ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, AddRoundKeyOutput[11]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1234, ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_10__FF_FF ( .D ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, AddRoundKeyOutput[10]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1238, ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_9__FF_FF ( .D ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, AddRoundKeyOutput[9]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1700, ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_8__FF_FF ( .D ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, AddRoundKeyOutput[8]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1232, ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_7__FF_FF ( .D ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, AddRoundKeyOutput[7]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1218, ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_6__FF_FF ( .D ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, AddRoundKeyOutput[6]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1222, ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_5__FF_FF ( .D ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, AddRoundKeyOutput[5]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1690, ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_4__FF_FF ( .D ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, AddRoundKeyOutput[4]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1216, ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_3__FF_FF ( .D ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, AddRoundKeyOutput[3]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1266, ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_2__FF_FF ( .D ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, AddRoundKeyOutput[2]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1270, ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_1__FF_FF ( .D ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, AddRoundKeyOutput[1]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1720, ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_LMDPL StateReg_s_current_state_reg_0__FF_FF ( .D ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, AddRoundKeyOutput[0]}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1264, ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_6__FF_FF ( .D (FSMUpdate[6]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[6]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_5__FF_FF ( .D (FSMUpdate[5]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[5]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_4__FF_FF ( .D (FSMUpdate[4]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[4]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_3__FF_FF ( .D (FSMUpdate[3]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[3]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_2__FF_FF ( .D (FSMUpdate[2]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[2]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_1__FF_FF ( .D (FSMUpdate[1]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[1]), .QN () ) ;
    reg_sr_LMDPL FSMRegInst_s_current_state_reg_0__FF_FF ( .D (FSMUpdate[0]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (FSMReg[0]), .QN () ) ;
    reg_sr_LMDPL selectsRegInst_s_current_state_reg_1__FF_FF ( .D (selectsNext[1]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (selectsReg[1]), .QN () ) ;
    reg_sr_LMDPL selectsRegInst_s_current_state_reg_0__FF_FF ( .D (selectsNext[0]), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (selectsReg[0]), .QN () ) ;
    reg_sr_LMDPL done_reg_FF_FF ( .D (done_internal), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (done), .QN () ) ;
endmodule
