/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC1_ClockGating_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [7:0] X_s4 ;
    input rst ;
    input [509:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output [7:0] Y_s4 ;
    output Synch ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_161 ;
    wire new_AGEMA_signal_162 ;
    wire new_AGEMA_signal_167 ;
    wire new_AGEMA_signal_168 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_181 ;
    wire new_AGEMA_signal_182 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;
    wire new_AGEMA_signal_593 ;
    wire new_AGEMA_signal_594 ;
    wire new_AGEMA_signal_595 ;
    wire new_AGEMA_signal_596 ;
    wire new_AGEMA_signal_597 ;
    wire new_AGEMA_signal_598 ;
    wire new_AGEMA_signal_599 ;
    wire new_AGEMA_signal_600 ;
    wire new_AGEMA_signal_601 ;
    wire new_AGEMA_signal_602 ;
    wire new_AGEMA_signal_603 ;
    wire new_AGEMA_signal_604 ;
    wire new_AGEMA_signal_605 ;
    wire new_AGEMA_signal_606 ;
    wire new_AGEMA_signal_607 ;
    wire new_AGEMA_signal_608 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;
    wire new_AGEMA_signal_656 ;
    wire new_AGEMA_signal_657 ;
    wire new_AGEMA_signal_658 ;
    wire new_AGEMA_signal_659 ;
    wire new_AGEMA_signal_660 ;
    wire new_AGEMA_signal_661 ;
    wire new_AGEMA_signal_662 ;
    wire new_AGEMA_signal_663 ;
    wire new_AGEMA_signal_664 ;
    wire new_AGEMA_signal_665 ;
    wire new_AGEMA_signal_666 ;
    wire new_AGEMA_signal_667 ;
    wire new_AGEMA_signal_668 ;
    wire new_AGEMA_signal_669 ;
    wire new_AGEMA_signal_670 ;
    wire new_AGEMA_signal_671 ;
    wire new_AGEMA_signal_672 ;
    wire new_AGEMA_signal_673 ;
    wire new_AGEMA_signal_674 ;
    wire new_AGEMA_signal_675 ;
    wire new_AGEMA_signal_676 ;
    wire new_AGEMA_signal_677 ;
    wire new_AGEMA_signal_678 ;
    wire new_AGEMA_signal_679 ;
    wire new_AGEMA_signal_680 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T1_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T2_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T3_U1 ( .a ({X_s4[7], X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T4_U1 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T5_U1 ( .a ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T6_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .c ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T7_U1 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T8_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .c ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, T8}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T9_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .c ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T10_U1 ( .a ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .b ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .c ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T11_U1 ( .a ({X_s4[6], X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T12_U1 ( .a ({X_s4[5], X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T13_U1 ( .a ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .b ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}), .c ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, new_AGEMA_signal_231, T13}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T14_U1 ( .a ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .b ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}), .c ({new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, new_AGEMA_signal_263, T14}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T15_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .b ({new_AGEMA_signal_206, new_AGEMA_signal_205, new_AGEMA_signal_204, new_AGEMA_signal_203, T11}), .c ({new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T15}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T16_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_189, new_AGEMA_signal_188, new_AGEMA_signal_187, T5}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}), .c ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T17_U1 ( .a ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}), .b ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .c ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T18_U1 ( .a ({X_s4[4], X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, new_AGEMA_signal_215, T18}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T19_U1 ( .a ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, new_AGEMA_signal_215, T18}), .c ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T20_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}), .c ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T21_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, T21}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T22_U1 ( .a ({new_AGEMA_signal_202, new_AGEMA_signal_201, new_AGEMA_signal_200, new_AGEMA_signal_199, T7}), .b ({new_AGEMA_signal_222, new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, T21}), .c ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T23_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .b ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}), .c ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, new_AGEMA_signal_275, T23}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T24_U1 ( .a ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .b ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}), .c ({new_AGEMA_signal_310, new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, T24}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T25_U1 ( .a ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}), .b ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}), .c ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, new_AGEMA_signal_311, T25}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T26_U1 ( .a ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .b ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .c ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, new_AGEMA_signal_279, T26}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_T27_U1 ( .a ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .b ({new_AGEMA_signal_210, new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, T12}), .c ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, new_AGEMA_signal_251, T27}) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M1_U1 ( .ina ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, new_AGEMA_signal_231, T13}), .inb ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .clk (clk), .rnd ({Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M2_U1 ( .ina ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, new_AGEMA_signal_275, T23}), .inb ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, T8}), .clk (clk), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15]}), .outt ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, M2}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M3_U1 ( .a ({new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, new_AGEMA_signal_263, T14}), .b ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}), .c ({new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M3}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M4_U1 ( .ina ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}), .inb ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .rnd ({Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, new_AGEMA_signal_287, M4}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M5_U1 ( .a ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, new_AGEMA_signal_287, M4}), .b ({new_AGEMA_signal_286, new_AGEMA_signal_285, new_AGEMA_signal_284, new_AGEMA_signal_283, M1}), .c ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, new_AGEMA_signal_323, M5}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M6_U1 ( .ina ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .inb ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .clk (clk), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45]}), .outt ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M7_U1 ( .ina ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}), .inb ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}), .clk (clk), .rnd ({Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M7}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M8_U1 ( .a ({new_AGEMA_signal_282, new_AGEMA_signal_281, new_AGEMA_signal_280, new_AGEMA_signal_279, T26}), .b ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}), .c ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, M8}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M9_U1 ( .ina ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}), .inb ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}), .clk (clk), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75]}), .outt ({new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M9}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M10_U1 ( .a ({new_AGEMA_signal_334, new_AGEMA_signal_333, new_AGEMA_signal_332, new_AGEMA_signal_331, M9}), .b ({new_AGEMA_signal_294, new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, M6}), .c ({new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M10}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M11_U1 ( .ina ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .inb ({new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T15}), .clk (clk), .rnd ({Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M12_U1 ( .ina ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}), .inb ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, new_AGEMA_signal_251, T27}), .clk (clk), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105]}), .outt ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, M12}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M13_U1 ( .a ({new_AGEMA_signal_306, new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, M12}), .b ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}), .c ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M14_U1 ( .ina ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .inb ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}), .clk (clk), .rnd ({Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, M14}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M15_U1 ( .a ({new_AGEMA_signal_342, new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, M14}), .b ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, new_AGEMA_signal_299, M11}), .c ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M16_U1 ( .a ({new_AGEMA_signal_322, new_AGEMA_signal_321, new_AGEMA_signal_320, new_AGEMA_signal_319, M3}), .b ({new_AGEMA_signal_318, new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, M2}), .c ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, M16}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M17_U1 ( .a ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, new_AGEMA_signal_323, M5}), .b ({new_AGEMA_signal_310, new_AGEMA_signal_309, new_AGEMA_signal_308, new_AGEMA_signal_307, T24}), .c ({new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M17}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M18_U1 ( .a ({new_AGEMA_signal_330, new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, M8}), .b ({new_AGEMA_signal_298, new_AGEMA_signal_297, new_AGEMA_signal_296, new_AGEMA_signal_295, M7}), .c ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, new_AGEMA_signal_359, M18}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M19_U1 ( .a ({new_AGEMA_signal_346, new_AGEMA_signal_345, new_AGEMA_signal_344, new_AGEMA_signal_343, M10}), .b ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}), .c ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, M19}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M20_U1 ( .a ({new_AGEMA_signal_354, new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, M16}), .b ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}), .c ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M21_U1 ( .a ({new_AGEMA_signal_358, new_AGEMA_signal_357, new_AGEMA_signal_356, new_AGEMA_signal_355, M17}), .b ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, new_AGEMA_signal_347, M15}), .c ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M22_U1 ( .a ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, new_AGEMA_signal_359, M18}), .b ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, new_AGEMA_signal_335, M13}), .c ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M23_U1 ( .a ({new_AGEMA_signal_366, new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, M19}), .b ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, new_AGEMA_signal_311, T25}), .c ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M24_U1 ( .a ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .b ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .c ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, new_AGEMA_signal_395, M24}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M27_U1 ( .a ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .b ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .c ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M25_U1 ( .ina ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .inb ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .clk (clk), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135]}), .outt ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M26_U1 ( .a ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, M26}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M28_U1 ( .a ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M28}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M31_U1 ( .ina ({new_AGEMA_signal_370, new_AGEMA_signal_369, new_AGEMA_signal_368, new_AGEMA_signal_367, M20}), .inb ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .clk (clk), .rnd ({Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, new_AGEMA_signal_407, M31}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M33_U1 ( .a ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, M27}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, M33}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M34_U1 ( .ina ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .inb ({new_AGEMA_signal_378, new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, M22}), .clk (clk), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165]}), .outt ({new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M34}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M36_U1 ( .a ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, new_AGEMA_signal_395, M24}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, new_AGEMA_signal_383, M25}), .c ({new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, new_AGEMA_signal_431, M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M29_U1 ( .ina ({new_AGEMA_signal_406, new_AGEMA_signal_405, new_AGEMA_signal_404, new_AGEMA_signal_403, M28}), .inb ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, M27}), .clk (clk), .rnd ({Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M29}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M30_U1 ( .ina ({new_AGEMA_signal_402, new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, M26}), .inb ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, new_AGEMA_signal_395, M24}), .clk (clk), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195]}), .outt ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, new_AGEMA_signal_419, M30}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M32_U1 ( .ina ({new_AGEMA_signal_390, new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, M27}), .inb ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, new_AGEMA_signal_407, M31}), .clk (clk), .rnd ({Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, M32}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M35_U1 ( .ina ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, new_AGEMA_signal_395, M24}), .inb ({new_AGEMA_signal_394, new_AGEMA_signal_393, new_AGEMA_signal_392, new_AGEMA_signal_391, M34}), .clk (clk), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225]}), .outt ({new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M35}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M37_U1 ( .a ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, new_AGEMA_signal_371, M21}), .b ({new_AGEMA_signal_418, new_AGEMA_signal_417, new_AGEMA_signal_416, new_AGEMA_signal_415, M29}), .c ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M38_U1 ( .a ({new_AGEMA_signal_426, new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, M32}), .b ({new_AGEMA_signal_414, new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, M33}), .c ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M39_U1 ( .a ({new_AGEMA_signal_382, new_AGEMA_signal_381, new_AGEMA_signal_380, new_AGEMA_signal_379, M23}), .b ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, new_AGEMA_signal_419, M30}), .c ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M40_U1 ( .a ({new_AGEMA_signal_430, new_AGEMA_signal_429, new_AGEMA_signal_428, new_AGEMA_signal_427, M35}), .b ({new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, new_AGEMA_signal_431, M36}), .c ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M41_U1 ( .a ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .c ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M42_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .c ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M43_U1 ( .a ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .b ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .c ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M44_U1 ( .a ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .b ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .c ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_M45_U1 ( .a ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .b ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .c ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M46_U1 ( .ina ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}), .inb ({new_AGEMA_signal_226, new_AGEMA_signal_225, new_AGEMA_signal_224, new_AGEMA_signal_223, T6}), .clk (clk), .rnd ({Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M47_U1 ( .ina ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .inb ({new_AGEMA_signal_258, new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, T8}), .clk (clk), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255]}), .outt ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, new_AGEMA_signal_467, M47}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M48_U1 ( .ina ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .inb ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .clk (clk), .rnd ({Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M49_U1 ( .ina ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}), .inb ({new_AGEMA_signal_242, new_AGEMA_signal_241, new_AGEMA_signal_240, new_AGEMA_signal_239, T16}), .clk (clk), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285]}), .outt ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, M49}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M50_U1 ( .ina ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .inb ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, new_AGEMA_signal_227, T9}), .clk (clk), .rnd ({Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M51_U1 ( .ina ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .inb ({new_AGEMA_signal_270, new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, T17}), .clk (clk), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315]}), .outt ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M52_U1 ( .ina ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .inb ({new_AGEMA_signal_238, new_AGEMA_signal_237, new_AGEMA_signal_236, new_AGEMA_signal_235, T15}), .clk (clk), .rnd ({Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M53_U1 ( .ina ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}), .inb ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, new_AGEMA_signal_251, T27}), .clk (clk), .rnd ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345]}), .outt ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M54_U1 ( .ina ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .inb ({new_AGEMA_signal_262, new_AGEMA_signal_261, new_AGEMA_signal_260, new_AGEMA_signal_259, T10}), .clk (clk), .rnd ({Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, new_AGEMA_signal_515, M54}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M55_U1 ( .ina ({new_AGEMA_signal_466, new_AGEMA_signal_465, new_AGEMA_signal_464, new_AGEMA_signal_463, M44}), .inb ({new_AGEMA_signal_234, new_AGEMA_signal_233, new_AGEMA_signal_232, new_AGEMA_signal_231, T13}), .clk (clk), .rnd ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375]}), .outt ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M56_U1 ( .ina ({new_AGEMA_signal_450, new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, M40}), .inb ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, new_AGEMA_signal_275, T23}), .clk (clk), .rnd ({Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M57_U1 ( .ina ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, new_AGEMA_signal_443, M39}), .inb ({new_AGEMA_signal_246, new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, T19}), .clk (clk), .rnd ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405]}), .outt ({new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, M57}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M58_U1 ( .ina ({new_AGEMA_signal_462, new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, M43}), .inb ({new_AGEMA_signal_178, new_AGEMA_signal_177, new_AGEMA_signal_176, new_AGEMA_signal_175, T3}), .clk (clk), .rnd ({Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .outt ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M59_U1 ( .ina ({new_AGEMA_signal_442, new_AGEMA_signal_441, new_AGEMA_signal_440, new_AGEMA_signal_439, M38}), .inb ({new_AGEMA_signal_250, new_AGEMA_signal_249, new_AGEMA_signal_248, new_AGEMA_signal_247, T22}), .clk (clk), .rnd ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435]}), .outt ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, new_AGEMA_signal_491, M59}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M60_U1 ( .ina ({new_AGEMA_signal_438, new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, M37}), .inb ({new_AGEMA_signal_274, new_AGEMA_signal_273, new_AGEMA_signal_272, new_AGEMA_signal_271, T20}), .clk (clk), .rnd ({Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .outt ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, M60}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M61_U1 ( .ina ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, new_AGEMA_signal_455, M42}), .inb ({new_AGEMA_signal_162, new_AGEMA_signal_161, new_AGEMA_signal_160, new_AGEMA_signal_159, T1}), .clk (clk), .rnd ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465]}), .outt ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M62_U1 ( .ina ({new_AGEMA_signal_502, new_AGEMA_signal_501, new_AGEMA_signal_500, new_AGEMA_signal_499, M45}), .inb ({new_AGEMA_signal_182, new_AGEMA_signal_181, new_AGEMA_signal_180, new_AGEMA_signal_179, T4}), .clk (clk), .rnd ({Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .outt ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(0)) AND_M63_U1 ( .ina ({new_AGEMA_signal_454, new_AGEMA_signal_453, new_AGEMA_signal_452, new_AGEMA_signal_451, M41}), .inb ({new_AGEMA_signal_170, new_AGEMA_signal_169, new_AGEMA_signal_168, new_AGEMA_signal_167, T2}), .clk (clk), .rnd ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495]}), .outt ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, M63}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L0_U1 ( .a ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .b ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}), .c ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L1_U1 ( .a ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}), .b ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}), .c ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L2_U1 ( .a ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}), .b ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}), .c ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L3_U1 ( .a ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, new_AGEMA_signal_467, M47}), .b ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}), .c ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L4_U1 ( .a ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, new_AGEMA_signal_515, M54}), .b ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}), .c ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L5_U1 ( .a ({new_AGEMA_signal_510, new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, M49}), .b ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .c ({new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, L5}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L6_U1 ( .a ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, new_AGEMA_signal_551, M62}), .b ({new_AGEMA_signal_570, new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, L5}), .c ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L7_U1 ( .a ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, new_AGEMA_signal_503, M46}), .b ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}), .c ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L8_U1 ( .a ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}), .b ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, new_AGEMA_signal_491, M59}), .c ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L9_U1 ( .a ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}), .b ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}), .c ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L10_U1 ( .a ({new_AGEMA_signal_550, new_AGEMA_signal_549, new_AGEMA_signal_548, new_AGEMA_signal_547, M53}), .b ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}), .c ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L11_U1 ( .a ({new_AGEMA_signal_498, new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, M60}), .b ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}), .c ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L12_U1 ( .a ({new_AGEMA_signal_474, new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, M48}), .b ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, new_AGEMA_signal_479, M51}), .c ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, L12}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L13_U1 ( .a ({new_AGEMA_signal_478, new_AGEMA_signal_477, new_AGEMA_signal_476, new_AGEMA_signal_475, M50}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .c ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, new_AGEMA_signal_623, L13}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L14_U1 ( .a ({new_AGEMA_signal_514, new_AGEMA_signal_513, new_AGEMA_signal_512, new_AGEMA_signal_511, M52}), .b ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, new_AGEMA_signal_527, M61}), .c ({new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, new_AGEMA_signal_571, L14}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L15_U1 ( .a ({new_AGEMA_signal_522, new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, M55}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, new_AGEMA_signal_575, L15}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L16_U1 ( .a ({new_AGEMA_signal_486, new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, M56}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .c ({new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, L16}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L17_U1 ( .a ({new_AGEMA_signal_490, new_AGEMA_signal_489, new_AGEMA_signal_488, new_AGEMA_signal_487, M57}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, L17}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L18_U1 ( .a ({new_AGEMA_signal_526, new_AGEMA_signal_525, new_AGEMA_signal_524, new_AGEMA_signal_523, M58}), .b ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}), .c ({new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, new_AGEMA_signal_583, L18}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L19_U1 ( .a ({new_AGEMA_signal_534, new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, M63}), .b ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, new_AGEMA_signal_563, L4}), .c ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, new_AGEMA_signal_611, L19}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L20_U1 ( .a ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, new_AGEMA_signal_587, L0}), .b ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .c ({new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, new_AGEMA_signal_631, L20}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L21_U1 ( .a ({new_AGEMA_signal_538, new_AGEMA_signal_537, new_AGEMA_signal_536, new_AGEMA_signal_535, L1}), .b ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}), .c ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, new_AGEMA_signal_635, L21}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L22_U1 ( .a ({new_AGEMA_signal_562, new_AGEMA_signal_561, new_AGEMA_signal_560, new_AGEMA_signal_559, L3}), .b ({new_AGEMA_signal_546, new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, L12}), .c ({new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, L22}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L23_U1 ( .a ({new_AGEMA_signal_586, new_AGEMA_signal_585, new_AGEMA_signal_584, new_AGEMA_signal_583, L18}), .b ({new_AGEMA_signal_558, new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, L2}), .c ({new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, new_AGEMA_signal_619, L23}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L24_U1 ( .a ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, new_AGEMA_signal_575, L15}), .b ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}), .c ({new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, L24}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L25_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}), .c ({new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, new_AGEMA_signal_643, L25}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L26_U1 ( .a ({new_AGEMA_signal_598, new_AGEMA_signal_597, new_AGEMA_signal_596, new_AGEMA_signal_595, L7}), .b ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, new_AGEMA_signal_599, L9}), .c ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, new_AGEMA_signal_647, L26}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L27_U1 ( .a ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, new_AGEMA_signal_539, L8}), .b ({new_AGEMA_signal_606, new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, L10}), .c ({new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, L27}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L28_U1 ( .a ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}), .b ({new_AGEMA_signal_574, new_AGEMA_signal_573, new_AGEMA_signal_572, new_AGEMA_signal_571, L14}), .c ({new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, new_AGEMA_signal_655, L28}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_L29_U1 ( .a ({new_AGEMA_signal_610, new_AGEMA_signal_609, new_AGEMA_signal_608, new_AGEMA_signal_607, L11}), .b ({new_AGEMA_signal_582, new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, L17}), .c ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, new_AGEMA_signal_659, L29}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S0_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_642, new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, L24}), .c ({new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, new_AGEMA_signal_667, O[7]}) ) ;
    xnor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S1_U1 ( .a ({new_AGEMA_signal_630, new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, L16}), .b ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, new_AGEMA_signal_647, L26}), .c ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, new_AGEMA_signal_671, O[6]}) ) ;
    xnor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S2_U1 ( .a ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, new_AGEMA_signal_611, L19}), .b ({new_AGEMA_signal_658, new_AGEMA_signal_657, new_AGEMA_signal_656, new_AGEMA_signal_655, L28}), .c ({new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, O[5]}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S3_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, new_AGEMA_signal_635, L21}), .c ({new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, new_AGEMA_signal_679, O[4]}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S4_U1 ( .a ({new_AGEMA_signal_634, new_AGEMA_signal_633, new_AGEMA_signal_632, new_AGEMA_signal_631, L20}), .b ({new_AGEMA_signal_618, new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, L22}), .c ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, new_AGEMA_signal_683, O[3]}) ) ;
    xor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S5_U1 ( .a ({new_AGEMA_signal_646, new_AGEMA_signal_645, new_AGEMA_signal_644, new_AGEMA_signal_643, L25}), .b ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, new_AGEMA_signal_659, L29}), .c ({new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, O[2]}) ) ;
    xnor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S6_U1 ( .a ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, new_AGEMA_signal_623, L13}), .b ({new_AGEMA_signal_654, new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, L27}), .c ({new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, new_AGEMA_signal_691, O[1]}) ) ;
    xnor_HPC1 #(.security_order(4), .pipeline(0)) XOR_S7_U1 ( .a ({new_AGEMA_signal_594, new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, L6}), .b ({new_AGEMA_signal_622, new_AGEMA_signal_621, new_AGEMA_signal_620, new_AGEMA_signal_619, L23}), .c ({new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, O[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_7_ ( .clk (clk_gated), .D ({new_AGEMA_signal_670, new_AGEMA_signal_669, new_AGEMA_signal_668, new_AGEMA_signal_667, O[7]}), .Q ({Y_s4[7], Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_6_ ( .clk (clk_gated), .D ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, new_AGEMA_signal_671, O[6]}), .Q ({Y_s4[6], Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_5_ ( .clk (clk_gated), .D ({new_AGEMA_signal_678, new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, O[5]}), .Q ({Y_s4[5], Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_4_ ( .clk (clk_gated), .D ({new_AGEMA_signal_682, new_AGEMA_signal_681, new_AGEMA_signal_680, new_AGEMA_signal_679, O[4]}), .Q ({Y_s4[4], Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_3_ ( .clk (clk_gated), .D ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, new_AGEMA_signal_683, O[3]}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_2_ ( .clk (clk_gated), .D ({new_AGEMA_signal_690, new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, O[2]}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_1_ ( .clk (clk_gated), .D ({new_AGEMA_signal_694, new_AGEMA_signal_693, new_AGEMA_signal_692, new_AGEMA_signal_691, O[1]}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) Y_reg_0_ ( .clk (clk_gated), .D ({new_AGEMA_signal_666, new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, O[0]}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
