library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.GHPC_pkg.all;

entity GHPC_Step1_0 is
   Generic (
      in_size	    : integer;
      out_size	    : integer; 
      fresh_size    : integer;
      low_latency   : integer;
      pipeline      : integer);
   Port(
	in0 		: in  std_logic_vector(in_size-1    downto 0);
	r   		: in  std_logic_vector(fresh_size-1 downto 0);
	clk 		: in  std_logic;
	Step1_reg	: out bus_array(0 to out_size-1, 2**in_size-1 downto 0));
end GHPC_Step1_0;


architecture Behavioral of GHPC_Step1_0 is


	type in_array  is array(natural range <>) of std_logic_vector(in_size-1  downto 0);
	type out_array is array(natural range <>) of std_logic_vector(out_size-1 downto 0);

	signal in0_comb		: in_array(0 to 2**in_size-1);
	signal FuncOut 		: out_array(0 to 2**in_size-1);
	signal Step1		: bus_array(0 to   out_size-1, 2**in_size-1 downto 0);

begin

	GEN_in0_comb: for I in 0 to 2**in_size-1 generate
		GEN_in0_bit: for J in 0 to in_size-1 generate
			in0_comb(I)(j) <= in0(J) when GetBit(I,in_size,J) = '0' else (not in0(J));
		end generate;
		
            FuncOut(I)(0) <= (in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(1) <= (in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(2) <= (in0_comb(I)(7)) xor (in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(3) <= (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(4) <= (in0_comb(I)(7)) xor (in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(6)) xor (in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(5) <= (in0_comb(I)(7)) xor (in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(6) <= (in0_comb(I)(7)) xor (in0_comb(I)(6)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
            FuncOut(I)(7) <= (in0_comb(I)(7)) xor (in0_comb(I)(7) and in0_comb(I)(5)) xor (in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5)) xor (in0_comb(I)(7) and in0_comb(I)(4)) xor (in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4)) xor (in0_comb(I)(5) and in0_comb(I)(4)) xor (in0_comb(I)(7) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3)) xor (in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3)) xor (in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2)) xor (in0_comb(I)(7) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1)) xor (in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1)) xor (in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(6) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(7) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0)) xor (in0_comb(I)(6) and in0_comb(I)(5) and in0_comb(I)(4) and in0_comb(I)(3) and in0_comb(I)(2) and in0_comb(I)(1) and in0_comb(I)(0));
                                                                    -- input:  in0_comb(I)
	end generate;

	---------------------------------

	GEN_out: for X in 0 to out_size-1 generate
		GEN_Step1_1: for I in 0 to 2**in_size-1 generate
		   GEN_normal: if (low_latency = 0) generate
                      Step1(X, I) <= r(X) xor FuncOut(I)(X);
                   end generate;

		   GEN_LL: if (low_latency /= 0) generate
                      Step1(X, I) <= r(I+X*(2**in_size)) xor FuncOut(I)(X);
                   end generate;
			
 		   reg_ins: entity work.reg
		   Port map(
		     clk	=> clk,
		     D		=> Step1(X, I),
		     Q		=> Step1_reg(X, I));
		end generate;	
	end generate;	
	
end Behavioral;
