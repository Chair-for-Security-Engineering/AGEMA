/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_Pipeline_d4 (X_s0, clk, X_s1, X_s2, X_s3, X_s4, Fresh, Y_s0, Y_s1, Y_s2, Y_s3, Y_s4);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [3:0] X_s3 ;
    input [3:0] X_s4 ;
    input [39:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    output [3:0] Y_s3 ;
    output [3:0] Y_s4 ;
    wire Q0 ;
    wire Q1 ;
    wire T0 ;
    wire Q2 ;
    wire T1 ;
    wire Q4 ;
    wire T2 ;
    wire L0 ;
    wire Q6 ;
    wire L1 ;
    wire Q7 ;
    wire T3 ;
    wire L2 ;
    wire L2_T1 ;
    wire L3 ;
    wire n2 ;
    wire [2:1] XX ;
    wire [3:0] YY ;
    wire new_AGEMA_signal_41 ;
    wire new_AGEMA_signal_42 ;
    wire new_AGEMA_signal_43 ;
    wire new_AGEMA_signal_44 ;
    wire new_AGEMA_signal_49 ;
    wire new_AGEMA_signal_50 ;
    wire new_AGEMA_signal_51 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_57 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_89 ;
    wire new_AGEMA_signal_90 ;
    wire new_AGEMA_signal_91 ;
    wire new_AGEMA_signal_92 ;
    wire new_AGEMA_signal_93 ;
    wire new_AGEMA_signal_94 ;
    wire new_AGEMA_signal_95 ;
    wire new_AGEMA_signal_96 ;
    wire new_AGEMA_signal_97 ;
    wire new_AGEMA_signal_98 ;
    wire new_AGEMA_signal_99 ;
    wire new_AGEMA_signal_100 ;
    wire new_AGEMA_signal_101 ;
    wire new_AGEMA_signal_102 ;
    wire new_AGEMA_signal_103 ;
    wire new_AGEMA_signal_104 ;
    wire new_AGEMA_signal_105 ;
    wire new_AGEMA_signal_106 ;
    wire new_AGEMA_signal_107 ;
    wire new_AGEMA_signal_108 ;
    wire new_AGEMA_signal_109 ;
    wire new_AGEMA_signal_110 ;
    wire new_AGEMA_signal_111 ;
    wire new_AGEMA_signal_112 ;
    wire new_AGEMA_signal_113 ;
    wire new_AGEMA_signal_114 ;
    wire new_AGEMA_signal_115 ;
    wire new_AGEMA_signal_116 ;
    wire new_AGEMA_signal_117 ;
    wire new_AGEMA_signal_118 ;
    wire new_AGEMA_signal_119 ;
    wire new_AGEMA_signal_120 ;
    wire new_AGEMA_signal_121 ;
    wire new_AGEMA_signal_122 ;
    wire new_AGEMA_signal_123 ;
    wire new_AGEMA_signal_124 ;
    wire new_AGEMA_signal_125 ;
    wire new_AGEMA_signal_126 ;
    wire new_AGEMA_signal_127 ;
    wire new_AGEMA_signal_128 ;
    wire new_AGEMA_signal_129 ;
    wire new_AGEMA_signal_130 ;
    wire new_AGEMA_signal_131 ;
    wire new_AGEMA_signal_132 ;
    wire new_AGEMA_signal_133 ;
    wire new_AGEMA_signal_134 ;
    wire new_AGEMA_signal_135 ;
    wire new_AGEMA_signal_136 ;
    wire new_AGEMA_signal_137 ;
    wire new_AGEMA_signal_138 ;
    wire new_AGEMA_signal_139 ;
    wire new_AGEMA_signal_140 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) U5 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_i1_U1 ( .a ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s4[3], X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .c ({new_AGEMA_signal_52, new_AGEMA_signal_51, new_AGEMA_signal_50, new_AGEMA_signal_49, XX[1]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR_i2_U1 ( .a ({X_s4[0], X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({X_s4[2], X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, new_AGEMA_signal_57, XX[2]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR0_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, new_AGEMA_signal_57, XX[2]}), .c ({new_AGEMA_signal_68, new_AGEMA_signal_67, new_AGEMA_signal_66, new_AGEMA_signal_65, Q0}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR1_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_52, new_AGEMA_signal_51, new_AGEMA_signal_50, new_AGEMA_signal_49, XX[1]}), .c ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, new_AGEMA_signal_69, Q1}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR3_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}), .c ({new_AGEMA_signal_76, new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, Q4}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR5_U1 ( .a ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, new_AGEMA_signal_57, XX[2]}), .b ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}), .c ({new_AGEMA_signal_80, new_AGEMA_signal_79, new_AGEMA_signal_78, new_AGEMA_signal_77, Q6}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR6_U1 ( .a ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, new_AGEMA_signal_69, Q1}), .b ({new_AGEMA_signal_80, new_AGEMA_signal_79, new_AGEMA_signal_78, new_AGEMA_signal_77, Q6}), .c ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, new_AGEMA_signal_93, L1}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR8_U1 ( .a ({X_s4[1], X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}), .c ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, new_AGEMA_signal_81, L2}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_26 ( .C (clk), .D (Q0), .Q (new_AGEMA_signal_197) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C (clk), .D (new_AGEMA_signal_65), .Q (new_AGEMA_signal_199) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C (clk), .D (new_AGEMA_signal_66), .Q (new_AGEMA_signal_201) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C (clk), .D (new_AGEMA_signal_67), .Q (new_AGEMA_signal_203) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C (clk), .D (new_AGEMA_signal_68), .Q (new_AGEMA_signal_205) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C (clk), .D (L1), .Q (new_AGEMA_signal_207) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C (clk), .D (new_AGEMA_signal_93), .Q (new_AGEMA_signal_209) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C (clk), .D (new_AGEMA_signal_94), .Q (new_AGEMA_signal_211) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C (clk), .D (new_AGEMA_signal_95), .Q (new_AGEMA_signal_213) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C (clk), .D (new_AGEMA_signal_96), .Q (new_AGEMA_signal_215) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C (clk), .D (XX[2]), .Q (new_AGEMA_signal_217) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C (clk), .D (new_AGEMA_signal_57), .Q (new_AGEMA_signal_219) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C (clk), .D (new_AGEMA_signal_58), .Q (new_AGEMA_signal_221) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C (clk), .D (new_AGEMA_signal_59), .Q (new_AGEMA_signal_223) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C (clk), .D (new_AGEMA_signal_60), .Q (new_AGEMA_signal_225) ) ;
    buf_clk new_AGEMA_reg_buffer_56 ( .C (clk), .D (XX[1]), .Q (new_AGEMA_signal_227) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C (clk), .D (new_AGEMA_signal_49), .Q (new_AGEMA_signal_229) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C (clk), .D (new_AGEMA_signal_50), .Q (new_AGEMA_signal_231) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C (clk), .D (new_AGEMA_signal_51), .Q (new_AGEMA_signal_233) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C (clk), .D (new_AGEMA_signal_52), .Q (new_AGEMA_signal_235) ) ;
    buf_clk new_AGEMA_reg_buffer_66 ( .C (clk), .D (X_s0[1]), .Q (new_AGEMA_signal_237) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C (clk), .D (X_s1[1]), .Q (new_AGEMA_signal_239) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C (clk), .D (X_s2[1]), .Q (new_AGEMA_signal_241) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C (clk), .D (X_s3[1]), .Q (new_AGEMA_signal_243) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C (clk), .D (X_s4[1]), .Q (new_AGEMA_signal_245) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C (clk), .D (Q6), .Q (new_AGEMA_signal_257) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C (clk), .D (new_AGEMA_signal_77), .Q (new_AGEMA_signal_259) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C (clk), .D (new_AGEMA_signal_78), .Q (new_AGEMA_signal_261) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C (clk), .D (new_AGEMA_signal_79), .Q (new_AGEMA_signal_263) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C (clk), .D (new_AGEMA_signal_80), .Q (new_AGEMA_signal_265) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C (clk), .D (L2), .Q (new_AGEMA_signal_267) ) ;
    buf_clk new_AGEMA_reg_buffer_100 ( .C (clk), .D (new_AGEMA_signal_81), .Q (new_AGEMA_signal_271) ) ;
    buf_clk new_AGEMA_reg_buffer_104 ( .C (clk), .D (new_AGEMA_signal_82), .Q (new_AGEMA_signal_275) ) ;
    buf_clk new_AGEMA_reg_buffer_108 ( .C (clk), .D (new_AGEMA_signal_83), .Q (new_AGEMA_signal_279) ) ;
    buf_clk new_AGEMA_reg_buffer_112 ( .C (clk), .D (new_AGEMA_signal_84), .Q (new_AGEMA_signal_283) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND1_U1 ( .a ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}), .b ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, new_AGEMA_signal_69, Q1}), .clk (clk), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_88, new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, T0}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR2_U1 ( .a ({new_AGEMA_signal_206, new_AGEMA_signal_204, new_AGEMA_signal_202, new_AGEMA_signal_200, new_AGEMA_signal_198}), .b ({new_AGEMA_signal_88, new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, T0}), .c ({new_AGEMA_signal_100, new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, Q2}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND3_U1 ( .a ({new_AGEMA_signal_44, new_AGEMA_signal_43, new_AGEMA_signal_42, new_AGEMA_signal_41, n2}), .b ({new_AGEMA_signal_76, new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, Q4}), .clk (clk), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, new_AGEMA_signal_89, T2}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR7_U1 ( .a ({new_AGEMA_signal_216, new_AGEMA_signal_214, new_AGEMA_signal_212, new_AGEMA_signal_210, new_AGEMA_signal_208}), .b ({new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, new_AGEMA_signal_89, T2}), .c ({new_AGEMA_signal_104, new_AGEMA_signal_103, new_AGEMA_signal_102, new_AGEMA_signal_101, Q7}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR11_U1 ( .a ({new_AGEMA_signal_226, new_AGEMA_signal_224, new_AGEMA_signal_222, new_AGEMA_signal_220, new_AGEMA_signal_218}), .b ({new_AGEMA_signal_88, new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, T0}), .c ({new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, new_AGEMA_signal_105, L3}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR12_U1 ( .a ({new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, new_AGEMA_signal_105, L3}), .b ({new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, new_AGEMA_signal_89, T2}), .c ({new_AGEMA_signal_124, new_AGEMA_signal_123, new_AGEMA_signal_122, new_AGEMA_signal_121, YY[1]}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR13_U1 ( .a ({new_AGEMA_signal_236, new_AGEMA_signal_234, new_AGEMA_signal_232, new_AGEMA_signal_230, new_AGEMA_signal_228}), .b ({new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, new_AGEMA_signal_89, T2}), .c ({new_AGEMA_signal_112, new_AGEMA_signal_111, new_AGEMA_signal_110, new_AGEMA_signal_109, YY[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C (clk), .D (new_AGEMA_signal_197), .Q (new_AGEMA_signal_198) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C (clk), .D (new_AGEMA_signal_199), .Q (new_AGEMA_signal_200) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C (clk), .D (new_AGEMA_signal_201), .Q (new_AGEMA_signal_202) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C (clk), .D (new_AGEMA_signal_203), .Q (new_AGEMA_signal_204) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C (clk), .D (new_AGEMA_signal_205), .Q (new_AGEMA_signal_206) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C (clk), .D (new_AGEMA_signal_207), .Q (new_AGEMA_signal_208) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C (clk), .D (new_AGEMA_signal_209), .Q (new_AGEMA_signal_210) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C (clk), .D (new_AGEMA_signal_211), .Q (new_AGEMA_signal_212) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C (clk), .D (new_AGEMA_signal_213), .Q (new_AGEMA_signal_214) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C (clk), .D (new_AGEMA_signal_215), .Q (new_AGEMA_signal_216) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C (clk), .D (new_AGEMA_signal_217), .Q (new_AGEMA_signal_218) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C (clk), .D (new_AGEMA_signal_219), .Q (new_AGEMA_signal_220) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C (clk), .D (new_AGEMA_signal_221), .Q (new_AGEMA_signal_222) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C (clk), .D (new_AGEMA_signal_223), .Q (new_AGEMA_signal_224) ) ;
    buf_clk new_AGEMA_reg_buffer_55 ( .C (clk), .D (new_AGEMA_signal_225), .Q (new_AGEMA_signal_226) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C (clk), .D (new_AGEMA_signal_227), .Q (new_AGEMA_signal_228) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C (clk), .D (new_AGEMA_signal_229), .Q (new_AGEMA_signal_230) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C (clk), .D (new_AGEMA_signal_231), .Q (new_AGEMA_signal_232) ) ;
    buf_clk new_AGEMA_reg_buffer_63 ( .C (clk), .D (new_AGEMA_signal_233), .Q (new_AGEMA_signal_234) ) ;
    buf_clk new_AGEMA_reg_buffer_65 ( .C (clk), .D (new_AGEMA_signal_235), .Q (new_AGEMA_signal_236) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C (clk), .D (new_AGEMA_signal_237), .Q (new_AGEMA_signal_238) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C (clk), .D (new_AGEMA_signal_239), .Q (new_AGEMA_signal_240) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C (clk), .D (new_AGEMA_signal_241), .Q (new_AGEMA_signal_242) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C (clk), .D (new_AGEMA_signal_243), .Q (new_AGEMA_signal_244) ) ;
    buf_clk new_AGEMA_reg_buffer_75 ( .C (clk), .D (new_AGEMA_signal_245), .Q (new_AGEMA_signal_246) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C (clk), .D (new_AGEMA_signal_257), .Q (new_AGEMA_signal_258) ) ;
    buf_clk new_AGEMA_reg_buffer_89 ( .C (clk), .D (new_AGEMA_signal_259), .Q (new_AGEMA_signal_260) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C (clk), .D (new_AGEMA_signal_261), .Q (new_AGEMA_signal_262) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C (clk), .D (new_AGEMA_signal_263), .Q (new_AGEMA_signal_264) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C (clk), .D (new_AGEMA_signal_265), .Q (new_AGEMA_signal_266) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C (clk), .D (new_AGEMA_signal_267), .Q (new_AGEMA_signal_268) ) ;
    buf_clk new_AGEMA_reg_buffer_101 ( .C (clk), .D (new_AGEMA_signal_271), .Q (new_AGEMA_signal_272) ) ;
    buf_clk new_AGEMA_reg_buffer_105 ( .C (clk), .D (new_AGEMA_signal_275), .Q (new_AGEMA_signal_276) ) ;
    buf_clk new_AGEMA_reg_buffer_109 ( .C (clk), .D (new_AGEMA_signal_279), .Q (new_AGEMA_signal_280) ) ;
    buf_clk new_AGEMA_reg_buffer_113 ( .C (clk), .D (new_AGEMA_signal_283), .Q (new_AGEMA_signal_284) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_76 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_247) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C (clk), .D (new_AGEMA_signal_89), .Q (new_AGEMA_signal_249) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C (clk), .D (new_AGEMA_signal_90), .Q (new_AGEMA_signal_251) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C (clk), .D (new_AGEMA_signal_91), .Q (new_AGEMA_signal_253) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C (clk), .D (new_AGEMA_signal_92), .Q (new_AGEMA_signal_255) ) ;
    buf_clk new_AGEMA_reg_buffer_98 ( .C (clk), .D (new_AGEMA_signal_268), .Q (new_AGEMA_signal_269) ) ;
    buf_clk new_AGEMA_reg_buffer_102 ( .C (clk), .D (new_AGEMA_signal_272), .Q (new_AGEMA_signal_273) ) ;
    buf_clk new_AGEMA_reg_buffer_106 ( .C (clk), .D (new_AGEMA_signal_276), .Q (new_AGEMA_signal_277) ) ;
    buf_clk new_AGEMA_reg_buffer_110 ( .C (clk), .D (new_AGEMA_signal_280), .Q (new_AGEMA_signal_281) ) ;
    buf_clk new_AGEMA_reg_buffer_114 ( .C (clk), .D (new_AGEMA_signal_284), .Q (new_AGEMA_signal_285) ) ;
    buf_clk new_AGEMA_reg_buffer_116 ( .C (clk), .D (L3), .Q (new_AGEMA_signal_287) ) ;
    buf_clk new_AGEMA_reg_buffer_118 ( .C (clk), .D (new_AGEMA_signal_105), .Q (new_AGEMA_signal_289) ) ;
    buf_clk new_AGEMA_reg_buffer_120 ( .C (clk), .D (new_AGEMA_signal_106), .Q (new_AGEMA_signal_291) ) ;
    buf_clk new_AGEMA_reg_buffer_122 ( .C (clk), .D (new_AGEMA_signal_107), .Q (new_AGEMA_signal_293) ) ;
    buf_clk new_AGEMA_reg_buffer_124 ( .C (clk), .D (new_AGEMA_signal_108), .Q (new_AGEMA_signal_295) ) ;
    buf_clk new_AGEMA_reg_buffer_126 ( .C (clk), .D (YY[1]), .Q (new_AGEMA_signal_297) ) ;
    buf_clk new_AGEMA_reg_buffer_128 ( .C (clk), .D (new_AGEMA_signal_121), .Q (new_AGEMA_signal_299) ) ;
    buf_clk new_AGEMA_reg_buffer_130 ( .C (clk), .D (new_AGEMA_signal_122), .Q (new_AGEMA_signal_301) ) ;
    buf_clk new_AGEMA_reg_buffer_132 ( .C (clk), .D (new_AGEMA_signal_123), .Q (new_AGEMA_signal_303) ) ;
    buf_clk new_AGEMA_reg_buffer_134 ( .C (clk), .D (new_AGEMA_signal_124), .Q (new_AGEMA_signal_305) ) ;
    buf_clk new_AGEMA_reg_buffer_136 ( .C (clk), .D (YY[0]), .Q (new_AGEMA_signal_307) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C (clk), .D (new_AGEMA_signal_109), .Q (new_AGEMA_signal_309) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C (clk), .D (new_AGEMA_signal_110), .Q (new_AGEMA_signal_311) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C (clk), .D (new_AGEMA_signal_111), .Q (new_AGEMA_signal_313) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C (clk), .D (new_AGEMA_signal_112), .Q (new_AGEMA_signal_315) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) AND2_U1 ( .a ({new_AGEMA_signal_246, new_AGEMA_signal_244, new_AGEMA_signal_242, new_AGEMA_signal_240, new_AGEMA_signal_238}), .b ({new_AGEMA_signal_100, new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, Q2}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_116, new_AGEMA_signal_115, new_AGEMA_signal_114, new_AGEMA_signal_113, T1}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR4_U1 ( .a ({new_AGEMA_signal_116, new_AGEMA_signal_115, new_AGEMA_signal_114, new_AGEMA_signal_113, T1}), .b ({new_AGEMA_signal_256, new_AGEMA_signal_254, new_AGEMA_signal_252, new_AGEMA_signal_250, new_AGEMA_signal_248}), .c ({new_AGEMA_signal_128, new_AGEMA_signal_127, new_AGEMA_signal_126, new_AGEMA_signal_125, L0}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) AND4_U1 ( .a ({new_AGEMA_signal_266, new_AGEMA_signal_264, new_AGEMA_signal_262, new_AGEMA_signal_260, new_AGEMA_signal_258}), .b ({new_AGEMA_signal_104, new_AGEMA_signal_103, new_AGEMA_signal_102, new_AGEMA_signal_101, Q7}), .clk (clk), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_120, new_AGEMA_signal_119, new_AGEMA_signal_118, new_AGEMA_signal_117, T3}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR81_U1 ( .a ({new_AGEMA_signal_286, new_AGEMA_signal_282, new_AGEMA_signal_278, new_AGEMA_signal_274, new_AGEMA_signal_270}), .b ({new_AGEMA_signal_116, new_AGEMA_signal_115, new_AGEMA_signal_114, new_AGEMA_signal_113, T1}), .c ({new_AGEMA_signal_132, new_AGEMA_signal_131, new_AGEMA_signal_130, new_AGEMA_signal_129, L2_T1}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) XOR9_U1 ( .a ({new_AGEMA_signal_132, new_AGEMA_signal_131, new_AGEMA_signal_130, new_AGEMA_signal_129, L2_T1}), .b ({new_AGEMA_signal_296, new_AGEMA_signal_294, new_AGEMA_signal_292, new_AGEMA_signal_290, new_AGEMA_signal_288}), .c ({new_AGEMA_signal_136, new_AGEMA_signal_135, new_AGEMA_signal_134, new_AGEMA_signal_133, YY[3]}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) XOR10_U1 ( .a ({new_AGEMA_signal_128, new_AGEMA_signal_127, new_AGEMA_signal_126, new_AGEMA_signal_125, L0}), .b ({new_AGEMA_signal_120, new_AGEMA_signal_119, new_AGEMA_signal_118, new_AGEMA_signal_117, T3}), .c ({new_AGEMA_signal_140, new_AGEMA_signal_139, new_AGEMA_signal_138, new_AGEMA_signal_137, YY[2]}) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C (clk), .D (new_AGEMA_signal_247), .Q (new_AGEMA_signal_248) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C (clk), .D (new_AGEMA_signal_249), .Q (new_AGEMA_signal_250) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C (clk), .D (new_AGEMA_signal_251), .Q (new_AGEMA_signal_252) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C (clk), .D (new_AGEMA_signal_253), .Q (new_AGEMA_signal_254) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C (clk), .D (new_AGEMA_signal_255), .Q (new_AGEMA_signal_256) ) ;
    buf_clk new_AGEMA_reg_buffer_99 ( .C (clk), .D (new_AGEMA_signal_269), .Q (new_AGEMA_signal_270) ) ;
    buf_clk new_AGEMA_reg_buffer_103 ( .C (clk), .D (new_AGEMA_signal_273), .Q (new_AGEMA_signal_274) ) ;
    buf_clk new_AGEMA_reg_buffer_107 ( .C (clk), .D (new_AGEMA_signal_277), .Q (new_AGEMA_signal_278) ) ;
    buf_clk new_AGEMA_reg_buffer_111 ( .C (clk), .D (new_AGEMA_signal_281), .Q (new_AGEMA_signal_282) ) ;
    buf_clk new_AGEMA_reg_buffer_115 ( .C (clk), .D (new_AGEMA_signal_285), .Q (new_AGEMA_signal_286) ) ;
    buf_clk new_AGEMA_reg_buffer_117 ( .C (clk), .D (new_AGEMA_signal_287), .Q (new_AGEMA_signal_288) ) ;
    buf_clk new_AGEMA_reg_buffer_119 ( .C (clk), .D (new_AGEMA_signal_289), .Q (new_AGEMA_signal_290) ) ;
    buf_clk new_AGEMA_reg_buffer_121 ( .C (clk), .D (new_AGEMA_signal_291), .Q (new_AGEMA_signal_292) ) ;
    buf_clk new_AGEMA_reg_buffer_123 ( .C (clk), .D (new_AGEMA_signal_293), .Q (new_AGEMA_signal_294) ) ;
    buf_clk new_AGEMA_reg_buffer_125 ( .C (clk), .D (new_AGEMA_signal_295), .Q (new_AGEMA_signal_296) ) ;
    buf_clk new_AGEMA_reg_buffer_127 ( .C (clk), .D (new_AGEMA_signal_297), .Q (new_AGEMA_signal_298) ) ;
    buf_clk new_AGEMA_reg_buffer_129 ( .C (clk), .D (new_AGEMA_signal_299), .Q (new_AGEMA_signal_300) ) ;
    buf_clk new_AGEMA_reg_buffer_131 ( .C (clk), .D (new_AGEMA_signal_301), .Q (new_AGEMA_signal_302) ) ;
    buf_clk new_AGEMA_reg_buffer_133 ( .C (clk), .D (new_AGEMA_signal_303), .Q (new_AGEMA_signal_304) ) ;
    buf_clk new_AGEMA_reg_buffer_135 ( .C (clk), .D (new_AGEMA_signal_305), .Q (new_AGEMA_signal_306) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C (clk), .D (new_AGEMA_signal_307), .Q (new_AGEMA_signal_308) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C (clk), .D (new_AGEMA_signal_309), .Q (new_AGEMA_signal_310) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C (clk), .D (new_AGEMA_signal_311), .Q (new_AGEMA_signal_312) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C (clk), .D (new_AGEMA_signal_313), .Q (new_AGEMA_signal_314) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C (clk), .D (new_AGEMA_signal_315), .Q (new_AGEMA_signal_316) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_306, new_AGEMA_signal_304, new_AGEMA_signal_302, new_AGEMA_signal_300, new_AGEMA_signal_298}), .Q ({Y_s4[3], Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_316, new_AGEMA_signal_314, new_AGEMA_signal_312, new_AGEMA_signal_310, new_AGEMA_signal_308}), .Q ({Y_s4[2], Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_136, new_AGEMA_signal_135, new_AGEMA_signal_134, new_AGEMA_signal_133, YY[3]}), .Q ({Y_s4[1], Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_140, new_AGEMA_signal_139, new_AGEMA_signal_138, new_AGEMA_signal_137, YY[2]}), .Q ({Y_s4[0], Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
