//
// taken from https://github.com/cassiersg/fullverif
//

`include "MSKref.vh"
localparam and_pini_mul_nrnd = d*(d-1)/2;
localparam and_pini_nrnd = ref_n_rnd + and_pini_mul_nrnd;