/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module AES_GHPC_ANF_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [159:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_423 ;
    wire signal_425 ;
    wire signal_427 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_443 ;
    wire signal_445 ;
    wire signal_447 ;
    wire signal_449 ;
    wire signal_451 ;
    wire signal_453 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_459 ;
    wire signal_461 ;
    wire signal_463 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_792 ;
    wire signal_912 ;
    wire signal_1032 ;
    wire signal_1152 ;
    wire signal_1272 ;
    wire signal_1392 ;
    wire signal_1512 ;
    wire signal_1632 ;
    wire signal_1752 ;
    wire signal_1872 ;
    wire signal_1992 ;
    wire signal_2112 ;
    wire signal_2232 ;
    wire signal_2352 ;
    wire signal_2472 ;
    wire signal_2592 ;
    wire signal_2597 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3874 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3882 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3890 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3898 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3906 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3914 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3922 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3930 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3938 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3946 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3954 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3962 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3970 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3978 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3986 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4394 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4402 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4410 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4474 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4482 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4490 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4498 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4506 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4514 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5403 ;
    wire signal_5405 ;
    wire signal_5407 ;
    wire signal_5409 ;
    wire signal_5411 ;
    wire signal_5413 ;
    wire signal_5415 ;
    wire signal_5417 ;
    wire signal_5419 ;
    wire signal_5421 ;
    wire signal_5423 ;
    wire signal_5425 ;
    wire signal_5427 ;
    wire signal_5429 ;
    wire signal_5431 ;
    wire signal_5433 ;
    wire signal_5435 ;
    wire signal_5437 ;
    wire signal_5439 ;
    wire signal_5441 ;
    wire signal_5443 ;
    wire signal_5445 ;
    wire signal_5447 ;
    wire signal_5449 ;
    wire signal_5451 ;
    wire signal_5453 ;
    wire signal_5455 ;
    wire signal_5457 ;
    wire signal_5459 ;
    wire signal_5461 ;
    wire signal_5463 ;
    wire signal_5465 ;
    wire signal_5467 ;
    wire signal_5469 ;
    wire signal_5471 ;
    wire signal_5473 ;
    wire signal_5475 ;
    wire signal_5477 ;
    wire signal_5479 ;
    wire signal_5481 ;
    wire signal_5483 ;
    wire signal_5485 ;
    wire signal_5487 ;
    wire signal_5489 ;
    wire signal_5491 ;
    wire signal_5493 ;
    wire signal_5495 ;
    wire signal_5497 ;
    wire signal_5499 ;
    wire signal_5501 ;
    wire signal_5503 ;
    wire signal_5505 ;
    wire signal_5507 ;
    wire signal_5509 ;
    wire signal_5511 ;
    wire signal_5513 ;
    wire signal_5515 ;
    wire signal_5517 ;
    wire signal_5519 ;
    wire signal_5521 ;
    wire signal_5523 ;
    wire signal_5525 ;
    wire signal_5527 ;
    wire signal_5529 ;
    wire signal_5531 ;
    wire signal_5533 ;
    wire signal_5535 ;
    wire signal_5537 ;
    wire signal_5539 ;
    wire signal_5541 ;
    wire signal_5543 ;
    wire signal_5545 ;
    wire signal_5547 ;
    wire signal_5549 ;
    wire signal_5551 ;
    wire signal_5553 ;
    wire signal_5555 ;
    wire signal_5557 ;
    wire signal_5559 ;
    wire signal_5561 ;
    wire signal_5563 ;
    wire signal_5565 ;
    wire signal_5567 ;
    wire signal_5569 ;
    wire signal_5571 ;
    wire signal_5573 ;
    wire signal_5575 ;
    wire signal_5577 ;
    wire signal_5579 ;
    wire signal_5581 ;
    wire signal_5583 ;
    wire signal_5585 ;
    wire signal_5587 ;
    wire signal_5589 ;
    wire signal_5591 ;
    wire signal_5593 ;
    wire signal_5595 ;
    wire signal_5597 ;
    wire signal_5599 ;
    wire signal_5601 ;
    wire signal_5603 ;
    wire signal_5605 ;
    wire signal_5607 ;
    wire signal_5609 ;
    wire signal_5611 ;
    wire signal_5613 ;
    wire signal_5615 ;
    wire signal_5617 ;
    wire signal_5619 ;
    wire signal_5621 ;
    wire signal_5623 ;
    wire signal_5625 ;
    wire signal_5627 ;
    wire signal_5629 ;
    wire signal_5631 ;
    wire signal_5633 ;
    wire signal_5635 ;
    wire signal_5637 ;
    wire signal_5639 ;
    wire signal_5641 ;
    wire signal_5643 ;
    wire signal_5645 ;
    wire signal_5647 ;
    wire signal_5649 ;
    wire signal_5651 ;
    wire signal_5653 ;
    wire signal_5655 ;
    wire signal_5657 ;
    wire signal_5659 ;
    wire signal_5661 ;
    wire signal_5663 ;
    wire signal_5665 ;
    wire signal_5667 ;
    wire signal_5669 ;
    wire signal_5671 ;
    wire signal_5673 ;
    wire signal_5675 ;
    wire signal_5677 ;
    wire signal_5679 ;
    wire signal_5681 ;
    wire signal_5683 ;
    wire signal_5685 ;
    wire signal_5687 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5723 ;
    wire signal_5725 ;
    wire signal_5727 ;
    wire signal_5729 ;
    wire signal_5731 ;
    wire signal_5733 ;
    wire signal_5735 ;
    wire signal_5737 ;
    wire signal_5739 ;
    wire signal_5741 ;
    wire signal_5743 ;
    wire signal_5745 ;
    wire signal_5747 ;
    wire signal_5749 ;
    wire signal_5751 ;
    wire signal_5753 ;
    wire signal_5755 ;
    wire signal_5757 ;
    wire signal_5759 ;
    wire signal_5761 ;
    wire signal_5763 ;
    wire signal_5765 ;
    wire signal_5767 ;
    wire signal_5769 ;
    wire signal_5771 ;
    wire signal_5773 ;
    wire signal_5775 ;
    wire signal_5777 ;
    wire signal_5779 ;
    wire signal_5781 ;
    wire signal_5783 ;
    wire signal_5785 ;
    wire signal_5787 ;
    wire signal_5789 ;
    wire signal_5791 ;
    wire signal_5793 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5829 ;
    wire signal_5831 ;
    wire signal_5833 ;
    wire signal_5835 ;
    wire signal_5837 ;
    wire signal_5839 ;
    wire signal_5841 ;
    wire signal_5843 ;
    wire signal_5845 ;
    wire signal_5847 ;
    wire signal_5849 ;
    wire signal_5851 ;
    wire signal_5853 ;
    wire signal_5855 ;
    wire signal_5857 ;
    wire signal_5859 ;
    wire signal_5861 ;
    wire signal_5863 ;
    wire signal_5865 ;
    wire signal_5867 ;
    wire signal_5869 ;
    wire signal_5871 ;
    wire signal_5873 ;
    wire signal_5875 ;
    wire signal_5877 ;
    wire signal_5879 ;
    wire signal_5881 ;
    wire signal_5883 ;
    wire signal_5885 ;
    wire signal_5887 ;
    wire signal_5889 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5925 ;
    wire signal_5927 ;
    wire signal_5929 ;
    wire signal_5931 ;
    wire signal_5933 ;
    wire signal_5935 ;
    wire signal_5937 ;
    wire signal_5939 ;
    wire signal_5941 ;
    wire signal_5943 ;
    wire signal_5945 ;
    wire signal_5947 ;
    wire signal_5949 ;
    wire signal_5951 ;
    wire signal_5953 ;
    wire signal_5955 ;
    wire signal_5957 ;
    wire signal_5959 ;
    wire signal_5961 ;
    wire signal_5963 ;
    wire signal_5965 ;
    wire signal_5967 ;
    wire signal_5969 ;
    wire signal_5971 ;
    wire signal_5973 ;
    wire signal_5975 ;
    wire signal_5977 ;
    wire signal_5979 ;
    wire signal_5981 ;
    wire signal_5983 ;
    wire signal_5985 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5997 ;
    wire signal_5999 ;
    wire signal_6001 ;
    wire signal_6003 ;
    wire signal_6005 ;
    wire signal_6007 ;
    wire signal_6009 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6016 ;
    wire signal_6018 ;
    wire signal_6020 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_400) ) ;
    INV_X1 cell_1 ( .A (signal_395), .ZN (signal_401) ) ;
    INV_X1 cell_2 ( .A (signal_395), .ZN (signal_398) ) ;
    INV_X1 cell_3 ( .A (signal_395), .ZN (signal_396) ) ;
    INV_X1 cell_4 ( .A (signal_395), .ZN (signal_397) ) ;
    INV_X1 cell_5 ( .A (signal_395), .ZN (signal_399) ) ;
    NOR2_X1 cell_6 ( .A1 (signal_406), .A2 (signal_411), .ZN (signal_395) ) ;
    INV_X1 cell_7 ( .A (signal_4388), .ZN (signal_406) ) ;
    INV_X1 cell_8 ( .A (signal_395), .ZN (signal_402) ) ;
    NOR2_X1 cell_9 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_404) ) ;
    INV_X1 cell_10 ( .A (signal_404), .ZN (signal_403) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_4388), .A2 (signal_403), .ZN (signal_4384) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_4388), .A2 (signal_4385), .ZN (signal_418) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_418), .A2 (signal_403), .ZN (signal_4383) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_4385), .A2 (signal_404), .ZN (signal_411) ) ;
    INV_X1 cell_15 ( .A (signal_4386), .ZN (signal_409) ) ;
    AND2_X1 cell_16 ( .A1 (signal_409), .A2 (signal_4387), .ZN (signal_414) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_418), .A2 (signal_414), .ZN (signal_405) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_402), .A2 (signal_405), .ZN (signal_4382) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_4385), .A2 (signal_406), .ZN (signal_416) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_414), .A2 (signal_416), .ZN (signal_408) ) ;
    NAND2_X1 cell_21 ( .A1 (signal_4385), .A2 (signal_4384), .ZN (signal_407) ) ;
    NAND2_X1 cell_22 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_4381) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_4387), .A2 (signal_409), .ZN (signal_412) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_418), .A2 (signal_412), .ZN (signal_410) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_411), .A2 (signal_410), .ZN (signal_4380) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_416), .A2 (signal_412), .ZN (signal_413) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_402), .A2 (signal_413), .ZN (signal_4379) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_156 ( .a ({signal_4549, signal_3870}), .b ({signal_4550, signal_4378}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_157 ( .a ({signal_4552, signal_3770}), .b ({signal_4553, signal_4278}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_158 ( .a ({signal_4555, signal_3769}), .b ({signal_4556, signal_4277}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_159 ( .a ({signal_4558, signal_3768}), .b ({signal_4559, signal_4276}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_160 ( .a ({signal_4561, signal_3767}), .b ({signal_4562, signal_4275}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_161 ( .a ({signal_4564, signal_3766}), .b ({signal_4565, signal_4274}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_162 ( .a ({signal_4567, signal_3765}), .b ({signal_4568, signal_4273}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_163 ( .a ({signal_4570, signal_3764}), .b ({signal_4571, signal_4272}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_164 ( .a ({signal_4573, signal_3763}), .b ({signal_4574, signal_4271}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_165 ( .a ({signal_4576, signal_3762}), .b ({signal_4577, signal_4270}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_166 ( .a ({signal_4579, signal_3761}), .b ({signal_4580, signal_4269}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_167 ( .a ({signal_4582, signal_3860}), .b ({signal_4583, signal_4368}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_168 ( .a ({signal_4585, signal_3760}), .b ({signal_4586, signal_4268}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_169 ( .a ({signal_4588, signal_3759}), .b ({signal_4589, signal_4267}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_170 ( .a ({signal_4591, signal_3758}), .b ({signal_4592, signal_4266}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_171 ( .a ({signal_4594, signal_3757}), .b ({signal_4595, signal_4265}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_172 ( .a ({signal_4597, signal_3756}), .b ({signal_4598, signal_4264}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_173 ( .a ({signal_4600, signal_3755}), .b ({signal_4601, signal_4263}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_174 ( .a ({signal_4603, signal_3754}), .b ({signal_4604, signal_4262}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_175 ( .a ({signal_4606, signal_3753}), .b ({signal_4607, signal_4261}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_176 ( .a ({signal_4609, signal_3752}), .b ({signal_4610, signal_4260}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_177 ( .a ({signal_4612, signal_3751}), .b ({signal_4613, signal_4259}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_178 ( .a ({signal_4615, signal_3859}), .b ({signal_4616, signal_4367}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_179 ( .a ({signal_4618, signal_3750}), .b ({signal_4619, signal_4258}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_180 ( .a ({signal_4621, signal_3749}), .b ({signal_4622, signal_4257}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_181 ( .a ({signal_4624, signal_3748}), .b ({signal_4625, signal_4256}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_182 ( .a ({signal_4627, signal_3747}), .b ({signal_4628, signal_4255}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_183 ( .a ({signal_4630, signal_3746}), .b ({signal_4631, signal_4254}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_184 ( .a ({signal_4633, signal_3745}), .b ({signal_4634, signal_4253}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_185 ( .a ({signal_4636, signal_3744}), .b ({signal_4637, signal_4252}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_186 ( .a ({signal_4639, signal_3743}), .b ({signal_4640, signal_4251}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_187 ( .a ({signal_4642, signal_3858}), .b ({signal_4643, signal_4366}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_188 ( .a ({signal_4645, signal_3857}), .b ({signal_4646, signal_4365}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_189 ( .a ({signal_4648, signal_3856}), .b ({signal_4649, signal_4364}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_190 ( .a ({signal_4651, signal_3855}), .b ({signal_4652, signal_4363}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_191 ( .a ({signal_4654, signal_3854}), .b ({signal_4655, signal_4362}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_192 ( .a ({signal_4657, signal_3853}), .b ({signal_4658, signal_4361}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_193 ( .a ({signal_4660, signal_3852}), .b ({signal_4661, signal_4360}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_194 ( .a ({signal_4663, signal_3851}), .b ({signal_4664, signal_4359}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_195 ( .a ({signal_4666, signal_3869}), .b ({signal_4667, signal_4377}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_196 ( .a ({signal_4669, signal_3850}), .b ({signal_4670, signal_4358}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_197 ( .a ({signal_4672, signal_3849}), .b ({signal_4673, signal_4357}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_198 ( .a ({signal_4675, signal_3848}), .b ({signal_4676, signal_4356}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_199 ( .a ({signal_4678, signal_3847}), .b ({signal_4679, signal_4355}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_200 ( .a ({signal_4681, signal_3846}), .b ({signal_4682, signal_4354}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_201 ( .a ({signal_4684, signal_3845}), .b ({signal_4685, signal_4353}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_202 ( .a ({signal_4687, signal_3844}), .b ({signal_4688, signal_4352}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_203 ( .a ({signal_4690, signal_3843}), .b ({signal_4691, signal_4351}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_204 ( .a ({signal_4693, signal_3842}), .b ({signal_4694, signal_4350}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_205 ( .a ({signal_4696, signal_3841}), .b ({signal_4697, signal_4349}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_206 ( .a ({signal_4699, signal_3868}), .b ({signal_4700, signal_4376}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_207 ( .a ({signal_4702, signal_3840}), .b ({signal_4703, signal_4348}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_208 ( .a ({signal_4705, signal_3839}), .b ({signal_4706, signal_4347}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_209 ( .a ({signal_4708, signal_3838}), .b ({signal_4709, signal_4346}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_210 ( .a ({signal_4711, signal_3837}), .b ({signal_4712, signal_4345}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_211 ( .a ({signal_4714, signal_3836}), .b ({signal_4715, signal_4344}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_212 ( .a ({signal_4717, signal_3835}), .b ({signal_4718, signal_4343}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_213 ( .a ({signal_4720, signal_3834}), .b ({signal_4721, signal_4342}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_214 ( .a ({signal_4723, signal_3833}), .b ({signal_4724, signal_4341}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_215 ( .a ({signal_4726, signal_3832}), .b ({signal_4727, signal_4340}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_216 ( .a ({signal_4729, signal_3831}), .b ({signal_4730, signal_4339}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_217 ( .a ({signal_4732, signal_3867}), .b ({signal_4733, signal_4375}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_218 ( .a ({signal_4735, signal_3830}), .b ({signal_4736, signal_4338}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_219 ( .a ({signal_4738, signal_3829}), .b ({signal_4739, signal_4337}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_220 ( .a ({signal_4741, signal_3828}), .b ({signal_4742, signal_4336}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_221 ( .a ({signal_4744, signal_3827}), .b ({signal_4745, signal_4335}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_222 ( .a ({signal_4747, signal_3826}), .b ({signal_4748, signal_4334}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_223 ( .a ({signal_4750, signal_3825}), .b ({signal_4751, signal_4333}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_224 ( .a ({signal_4753, signal_3824}), .b ({signal_4754, signal_4332}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_225 ( .a ({signal_4756, signal_3823}), .b ({signal_4757, signal_4331}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_226 ( .a ({signal_4759, signal_3822}), .b ({signal_4760, signal_4330}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_227 ( .a ({signal_4762, signal_3821}), .b ({signal_4763, signal_4329}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_228 ( .a ({signal_4765, signal_3866}), .b ({signal_4766, signal_4374}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_229 ( .a ({signal_4768, signal_3820}), .b ({signal_4769, signal_4328}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_230 ( .a ({signal_4771, signal_3819}), .b ({signal_4772, signal_4327}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_231 ( .a ({signal_4774, signal_3818}), .b ({signal_4775, signal_4326}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_232 ( .a ({signal_4777, signal_3817}), .b ({signal_4778, signal_4325}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_233 ( .a ({signal_4780, signal_3816}), .b ({signal_4781, signal_4324}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_234 ( .a ({signal_4783, signal_3815}), .b ({signal_4784, signal_4323}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_235 ( .a ({signal_4786, signal_3814}), .b ({signal_4787, signal_4322}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_236 ( .a ({signal_4789, signal_3813}), .b ({signal_4790, signal_4321}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_237 ( .a ({signal_4792, signal_3812}), .b ({signal_4793, signal_4320}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_238 ( .a ({signal_4795, signal_3811}), .b ({signal_4796, signal_4319}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_239 ( .a ({signal_4798, signal_3865}), .b ({signal_4799, signal_4373}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_240 ( .a ({signal_4801, signal_3810}), .b ({signal_4802, signal_4318}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_241 ( .a ({signal_4804, signal_3809}), .b ({signal_4805, signal_4317}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_242 ( .a ({signal_4807, signal_3808}), .b ({signal_4808, signal_4316}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_243 ( .a ({signal_4810, signal_3807}), .b ({signal_4811, signal_4315}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_244 ( .a ({signal_4813, signal_3806}), .b ({signal_4814, signal_4314}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_245 ( .a ({signal_4816, signal_3805}), .b ({signal_4817, signal_4313}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_246 ( .a ({signal_4819, signal_3804}), .b ({signal_4820, signal_4312}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_247 ( .a ({signal_4822, signal_3803}), .b ({signal_4823, signal_4311}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_248 ( .a ({signal_4825, signal_3802}), .b ({signal_4826, signal_4310}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_249 ( .a ({signal_4828, signal_3801}), .b ({signal_4829, signal_4309}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_250 ( .a ({signal_4831, signal_3864}), .b ({signal_4832, signal_4372}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_251 ( .a ({signal_4834, signal_3800}), .b ({signal_4835, signal_4308}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_252 ( .a ({signal_4837, signal_3799}), .b ({signal_4838, signal_4307}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_253 ( .a ({signal_4840, signal_3798}), .b ({signal_4841, signal_4306}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_254 ( .a ({signal_4843, signal_3797}), .b ({signal_4844, signal_4305}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_255 ( .a ({signal_4846, signal_3796}), .b ({signal_4847, signal_4304}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_256 ( .a ({signal_4849, signal_3795}), .b ({signal_4850, signal_4303}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_257 ( .a ({signal_4852, signal_3794}), .b ({signal_4853, signal_4302}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_258 ( .a ({signal_4855, signal_3793}), .b ({signal_4856, signal_4301}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_259 ( .a ({signal_4858, signal_3792}), .b ({signal_4859, signal_4300}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_260 ( .a ({signal_4861, signal_3791}), .b ({signal_4862, signal_4299}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_261 ( .a ({signal_4864, signal_3863}), .b ({signal_4865, signal_4371}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_262 ( .a ({signal_4867, signal_3790}), .b ({signal_4868, signal_4298}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_263 ( .a ({signal_4870, signal_3789}), .b ({signal_4871, signal_4297}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_264 ( .a ({signal_4873, signal_3788}), .b ({signal_4874, signal_4296}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_265 ( .a ({signal_4876, signal_3787}), .b ({signal_4877, signal_4295}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_266 ( .a ({signal_4879, signal_3786}), .b ({signal_4880, signal_4294}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_267 ( .a ({signal_4882, signal_3785}), .b ({signal_4883, signal_4293}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_268 ( .a ({signal_4885, signal_3784}), .b ({signal_4886, signal_4292}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_269 ( .a ({signal_4888, signal_3783}), .b ({signal_4889, signal_4291}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_270 ( .a ({signal_4891, signal_3782}), .b ({signal_4892, signal_4290}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_271 ( .a ({signal_4894, signal_3781}), .b ({signal_4895, signal_4289}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_272 ( .a ({signal_4897, signal_3862}), .b ({signal_4898, signal_4370}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_273 ( .a ({signal_4900, signal_3780}), .b ({signal_4901, signal_4288}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_274 ( .a ({signal_4903, signal_3779}), .b ({signal_4904, signal_4287}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_275 ( .a ({signal_4906, signal_3778}), .b ({signal_4907, signal_4286}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_276 ( .a ({signal_4909, signal_3777}), .b ({signal_4910, signal_4285}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_277 ( .a ({signal_4912, signal_3776}), .b ({signal_4913, signal_4284}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_278 ( .a ({signal_4915, signal_3775}), .b ({signal_4916, signal_4283}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_279 ( .a ({signal_4918, signal_3774}), .b ({signal_4919, signal_4282}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_280 ( .a ({signal_4921, signal_3773}), .b ({signal_4922, signal_4281}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_281 ( .a ({signal_4924, signal_3772}), .b ({signal_4925, signal_4280}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_282 ( .a ({signal_4927, signal_3771}), .b ({signal_4928, signal_4279}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_283 ( .a ({signal_4930, signal_3861}), .b ({signal_4931, signal_4369}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 cell_284 ( .A1 (signal_4385), .A2 (signal_414), .ZN (signal_415) ) ;
    NOR2_X1 cell_285 ( .A1 (signal_4388), .A2 (signal_415), .ZN (done) ) ;
    INV_X1 cell_286 ( .A (signal_416), .ZN (signal_417) ) ;
    NAND2_X1 cell_287 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_419) ) ;
    NOR2_X1 cell_288 ( .A1 (signal_417), .A2 (signal_419), .ZN (signal_393) ) ;
    INV_X1 cell_289 ( .A (signal_418), .ZN (signal_420) ) ;
    NOR2_X1 cell_290 ( .A1 (signal_420), .A2 (signal_419), .ZN (signal_394) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_679 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_4933, signal_792}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_807 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_4934, signal_912}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_935 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_4935, signal_1032}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1063 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_4936, signal_1152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1191 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_4937, signal_1272}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1319 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_4938, signal_1392}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1447 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_4939, signal_1512}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1575 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_4940, signal_1632}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1703 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_4941, signal_1752}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1831 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_4942, signal_1872}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1959 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_4943, signal_1992}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2087 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_4944, signal_2112}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2215 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_4945, signal_2232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2343 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_4946, signal_2352}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2471 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_4947, signal_2472}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2599 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_4948, signal_2592}) ) ;
    INV_X1 cell_4187 ( .A (signal_3597), .ZN (signal_3607) ) ;
    MUX2_X1 cell_4188 ( .S (signal_3609), .A (signal_3598), .B (signal_3599), .Z (signal_3597) ) ;
    NOR2_X1 cell_4189 ( .A1 (reset), .A2 (signal_3600), .ZN (signal_3610) ) ;
    XNOR2_X1 cell_4190 ( .A (signal_4388), .B (signal_4387), .ZN (signal_3600) ) ;
    MUX2_X1 cell_4191 ( .S (signal_4385), .A (signal_3601), .B (signal_3602), .Z (signal_3608) ) ;
    NAND2_X1 cell_4192 ( .A1 (signal_3598), .A2 (signal_3603), .ZN (signal_3602) ) ;
    NAND2_X1 cell_4193 ( .A1 (signal_3609), .A2 (signal_3606), .ZN (signal_3603) ) ;
    NOR2_X1 cell_4194 ( .A1 (signal_3604), .A2 (signal_3612), .ZN (signal_3598) ) ;
    NOR2_X1 cell_4195 ( .A1 (signal_4387), .A2 (reset), .ZN (signal_3604) ) ;
    NOR2_X1 cell_4196 ( .A1 (signal_3609), .A2 (signal_3599), .ZN (signal_3601) ) ;
    NAND2_X1 cell_4197 ( .A1 (signal_4387), .A2 (signal_3605), .ZN (signal_3599) ) ;
    NOR2_X1 cell_4198 ( .A1 (reset), .A2 (signal_3611), .ZN (signal_3605) ) ;
    NOR2_X1 cell_4199 ( .A1 (reset), .A2 (signal_4388), .ZN (signal_3612) ) ;
    INV_X1 cell_4200 ( .A (reset), .ZN (signal_3606) ) ;
    INV_X1 cell_4201 ( .A (signal_4388), .ZN (signal_3611) ) ;
    INV_X1 cell_4205 ( .A (signal_4386), .ZN (signal_3609) ) ;

    /* cells in depth 1 */
    buf_clk cell_4210 ( .C (clk), .D (signal_402), .Q (signal_6181) ) ;
    buf_clk cell_4212 ( .C (clk), .D (signal_396), .Q (signal_6183) ) ;
    buf_clk cell_4214 ( .C (clk), .D (signal_397), .Q (signal_6185) ) ;
    buf_clk cell_4216 ( .C (clk), .D (signal_398), .Q (signal_6187) ) ;
    buf_clk cell_4218 ( .C (clk), .D (signal_399), .Q (signal_6189) ) ;
    buf_clk cell_4220 ( .C (clk), .D (signal_400), .Q (signal_6191) ) ;
    buf_clk cell_4222 ( .C (clk), .D (signal_401), .Q (signal_6193) ) ;
    buf_clk cell_4224 ( .C (clk), .D (reset), .Q (signal_6195) ) ;
    buf_clk cell_4226 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_6197) ) ;
    buf_clk cell_4228 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_6199) ) ;
    buf_clk cell_4230 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_6201) ) ;
    buf_clk cell_4232 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_6203) ) ;
    buf_clk cell_4234 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_6205) ) ;
    buf_clk cell_4236 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_6207) ) ;
    buf_clk cell_4238 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_6209) ) ;
    buf_clk cell_4240 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_6211) ) ;
    buf_clk cell_4242 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_6213) ) ;
    buf_clk cell_4244 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_6215) ) ;
    buf_clk cell_4246 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_6217) ) ;
    buf_clk cell_4248 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_6219) ) ;
    buf_clk cell_4250 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_6221) ) ;
    buf_clk cell_4252 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_6223) ) ;
    buf_clk cell_4254 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_6225) ) ;
    buf_clk cell_4256 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_6227) ) ;
    buf_clk cell_4258 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_6229) ) ;
    buf_clk cell_4260 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_6231) ) ;
    buf_clk cell_4262 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_6233) ) ;
    buf_clk cell_4264 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_6235) ) ;
    buf_clk cell_4266 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_6237) ) ;
    buf_clk cell_4268 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_6239) ) ;
    buf_clk cell_4270 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_6241) ) ;
    buf_clk cell_4272 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_6243) ) ;
    buf_clk cell_4274 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_6245) ) ;
    buf_clk cell_4276 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_6247) ) ;
    buf_clk cell_4278 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_6249) ) ;
    buf_clk cell_4280 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_6251) ) ;
    buf_clk cell_4282 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_6253) ) ;
    buf_clk cell_4284 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_6255) ) ;
    buf_clk cell_4286 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_6257) ) ;
    buf_clk cell_4288 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_6259) ) ;
    buf_clk cell_4290 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_6261) ) ;
    buf_clk cell_4292 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_6263) ) ;
    buf_clk cell_4294 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_6265) ) ;
    buf_clk cell_4296 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_6267) ) ;
    buf_clk cell_4298 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_6269) ) ;
    buf_clk cell_4300 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_6271) ) ;
    buf_clk cell_4302 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_6273) ) ;
    buf_clk cell_4304 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_6275) ) ;
    buf_clk cell_4306 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_6277) ) ;
    buf_clk cell_4308 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_6279) ) ;
    buf_clk cell_4310 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_6281) ) ;
    buf_clk cell_4312 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_6283) ) ;
    buf_clk cell_4314 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_6285) ) ;
    buf_clk cell_4316 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_6287) ) ;
    buf_clk cell_4318 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_6289) ) ;
    buf_clk cell_4320 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_6291) ) ;
    buf_clk cell_4322 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_6293) ) ;
    buf_clk cell_4324 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_6295) ) ;
    buf_clk cell_4326 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_6297) ) ;
    buf_clk cell_4328 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_6299) ) ;
    buf_clk cell_4330 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_6301) ) ;
    buf_clk cell_4332 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_6303) ) ;
    buf_clk cell_4334 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_6305) ) ;
    buf_clk cell_4336 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_6307) ) ;
    buf_clk cell_4338 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_6309) ) ;
    buf_clk cell_4340 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_6311) ) ;
    buf_clk cell_4342 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_6313) ) ;
    buf_clk cell_4344 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_6315) ) ;
    buf_clk cell_4346 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_6317) ) ;
    buf_clk cell_4348 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_6319) ) ;
    buf_clk cell_4350 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_6321) ) ;
    buf_clk cell_4352 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_6323) ) ;
    buf_clk cell_4354 ( .C (clk), .D (plaintext_s0[32]), .Q (signal_6325) ) ;
    buf_clk cell_4356 ( .C (clk), .D (plaintext_s1[32]), .Q (signal_6327) ) ;
    buf_clk cell_4358 ( .C (clk), .D (plaintext_s0[33]), .Q (signal_6329) ) ;
    buf_clk cell_4360 ( .C (clk), .D (plaintext_s1[33]), .Q (signal_6331) ) ;
    buf_clk cell_4362 ( .C (clk), .D (plaintext_s0[34]), .Q (signal_6333) ) ;
    buf_clk cell_4364 ( .C (clk), .D (plaintext_s1[34]), .Q (signal_6335) ) ;
    buf_clk cell_4366 ( .C (clk), .D (plaintext_s0[35]), .Q (signal_6337) ) ;
    buf_clk cell_4368 ( .C (clk), .D (plaintext_s1[35]), .Q (signal_6339) ) ;
    buf_clk cell_4370 ( .C (clk), .D (plaintext_s0[36]), .Q (signal_6341) ) ;
    buf_clk cell_4372 ( .C (clk), .D (plaintext_s1[36]), .Q (signal_6343) ) ;
    buf_clk cell_4374 ( .C (clk), .D (plaintext_s0[37]), .Q (signal_6345) ) ;
    buf_clk cell_4376 ( .C (clk), .D (plaintext_s1[37]), .Q (signal_6347) ) ;
    buf_clk cell_4378 ( .C (clk), .D (plaintext_s0[38]), .Q (signal_6349) ) ;
    buf_clk cell_4380 ( .C (clk), .D (plaintext_s1[38]), .Q (signal_6351) ) ;
    buf_clk cell_4382 ( .C (clk), .D (plaintext_s0[39]), .Q (signal_6353) ) ;
    buf_clk cell_4384 ( .C (clk), .D (plaintext_s1[39]), .Q (signal_6355) ) ;
    buf_clk cell_4386 ( .C (clk), .D (plaintext_s0[40]), .Q (signal_6357) ) ;
    buf_clk cell_4388 ( .C (clk), .D (plaintext_s1[40]), .Q (signal_6359) ) ;
    buf_clk cell_4390 ( .C (clk), .D (plaintext_s0[41]), .Q (signal_6361) ) ;
    buf_clk cell_4392 ( .C (clk), .D (plaintext_s1[41]), .Q (signal_6363) ) ;
    buf_clk cell_4394 ( .C (clk), .D (plaintext_s0[42]), .Q (signal_6365) ) ;
    buf_clk cell_4396 ( .C (clk), .D (plaintext_s1[42]), .Q (signal_6367) ) ;
    buf_clk cell_4398 ( .C (clk), .D (plaintext_s0[43]), .Q (signal_6369) ) ;
    buf_clk cell_4400 ( .C (clk), .D (plaintext_s1[43]), .Q (signal_6371) ) ;
    buf_clk cell_4402 ( .C (clk), .D (plaintext_s0[44]), .Q (signal_6373) ) ;
    buf_clk cell_4404 ( .C (clk), .D (plaintext_s1[44]), .Q (signal_6375) ) ;
    buf_clk cell_4406 ( .C (clk), .D (plaintext_s0[45]), .Q (signal_6377) ) ;
    buf_clk cell_4408 ( .C (clk), .D (plaintext_s1[45]), .Q (signal_6379) ) ;
    buf_clk cell_4410 ( .C (clk), .D (plaintext_s0[46]), .Q (signal_6381) ) ;
    buf_clk cell_4412 ( .C (clk), .D (plaintext_s1[46]), .Q (signal_6383) ) ;
    buf_clk cell_4414 ( .C (clk), .D (plaintext_s0[47]), .Q (signal_6385) ) ;
    buf_clk cell_4416 ( .C (clk), .D (plaintext_s1[47]), .Q (signal_6387) ) ;
    buf_clk cell_4418 ( .C (clk), .D (plaintext_s0[48]), .Q (signal_6389) ) ;
    buf_clk cell_4420 ( .C (clk), .D (plaintext_s1[48]), .Q (signal_6391) ) ;
    buf_clk cell_4422 ( .C (clk), .D (plaintext_s0[49]), .Q (signal_6393) ) ;
    buf_clk cell_4424 ( .C (clk), .D (plaintext_s1[49]), .Q (signal_6395) ) ;
    buf_clk cell_4426 ( .C (clk), .D (plaintext_s0[50]), .Q (signal_6397) ) ;
    buf_clk cell_4428 ( .C (clk), .D (plaintext_s1[50]), .Q (signal_6399) ) ;
    buf_clk cell_4430 ( .C (clk), .D (plaintext_s0[51]), .Q (signal_6401) ) ;
    buf_clk cell_4432 ( .C (clk), .D (plaintext_s1[51]), .Q (signal_6403) ) ;
    buf_clk cell_4434 ( .C (clk), .D (plaintext_s0[52]), .Q (signal_6405) ) ;
    buf_clk cell_4436 ( .C (clk), .D (plaintext_s1[52]), .Q (signal_6407) ) ;
    buf_clk cell_4438 ( .C (clk), .D (plaintext_s0[53]), .Q (signal_6409) ) ;
    buf_clk cell_4440 ( .C (clk), .D (plaintext_s1[53]), .Q (signal_6411) ) ;
    buf_clk cell_4442 ( .C (clk), .D (plaintext_s0[54]), .Q (signal_6413) ) ;
    buf_clk cell_4444 ( .C (clk), .D (plaintext_s1[54]), .Q (signal_6415) ) ;
    buf_clk cell_4446 ( .C (clk), .D (plaintext_s0[55]), .Q (signal_6417) ) ;
    buf_clk cell_4448 ( .C (clk), .D (plaintext_s1[55]), .Q (signal_6419) ) ;
    buf_clk cell_4450 ( .C (clk), .D (plaintext_s0[56]), .Q (signal_6421) ) ;
    buf_clk cell_4452 ( .C (clk), .D (plaintext_s1[56]), .Q (signal_6423) ) ;
    buf_clk cell_4454 ( .C (clk), .D (plaintext_s0[57]), .Q (signal_6425) ) ;
    buf_clk cell_4456 ( .C (clk), .D (plaintext_s1[57]), .Q (signal_6427) ) ;
    buf_clk cell_4458 ( .C (clk), .D (plaintext_s0[58]), .Q (signal_6429) ) ;
    buf_clk cell_4460 ( .C (clk), .D (plaintext_s1[58]), .Q (signal_6431) ) ;
    buf_clk cell_4462 ( .C (clk), .D (plaintext_s0[59]), .Q (signal_6433) ) ;
    buf_clk cell_4464 ( .C (clk), .D (plaintext_s1[59]), .Q (signal_6435) ) ;
    buf_clk cell_4466 ( .C (clk), .D (plaintext_s0[60]), .Q (signal_6437) ) ;
    buf_clk cell_4468 ( .C (clk), .D (plaintext_s1[60]), .Q (signal_6439) ) ;
    buf_clk cell_4470 ( .C (clk), .D (plaintext_s0[61]), .Q (signal_6441) ) ;
    buf_clk cell_4472 ( .C (clk), .D (plaintext_s1[61]), .Q (signal_6443) ) ;
    buf_clk cell_4474 ( .C (clk), .D (plaintext_s0[62]), .Q (signal_6445) ) ;
    buf_clk cell_4476 ( .C (clk), .D (plaintext_s1[62]), .Q (signal_6447) ) ;
    buf_clk cell_4478 ( .C (clk), .D (plaintext_s0[63]), .Q (signal_6449) ) ;
    buf_clk cell_4480 ( .C (clk), .D (plaintext_s1[63]), .Q (signal_6451) ) ;
    buf_clk cell_4482 ( .C (clk), .D (plaintext_s0[64]), .Q (signal_6453) ) ;
    buf_clk cell_4484 ( .C (clk), .D (plaintext_s1[64]), .Q (signal_6455) ) ;
    buf_clk cell_4486 ( .C (clk), .D (plaintext_s0[65]), .Q (signal_6457) ) ;
    buf_clk cell_4488 ( .C (clk), .D (plaintext_s1[65]), .Q (signal_6459) ) ;
    buf_clk cell_4490 ( .C (clk), .D (plaintext_s0[66]), .Q (signal_6461) ) ;
    buf_clk cell_4492 ( .C (clk), .D (plaintext_s1[66]), .Q (signal_6463) ) ;
    buf_clk cell_4494 ( .C (clk), .D (plaintext_s0[67]), .Q (signal_6465) ) ;
    buf_clk cell_4496 ( .C (clk), .D (plaintext_s1[67]), .Q (signal_6467) ) ;
    buf_clk cell_4498 ( .C (clk), .D (plaintext_s0[68]), .Q (signal_6469) ) ;
    buf_clk cell_4500 ( .C (clk), .D (plaintext_s1[68]), .Q (signal_6471) ) ;
    buf_clk cell_4502 ( .C (clk), .D (plaintext_s0[69]), .Q (signal_6473) ) ;
    buf_clk cell_4504 ( .C (clk), .D (plaintext_s1[69]), .Q (signal_6475) ) ;
    buf_clk cell_4506 ( .C (clk), .D (plaintext_s0[70]), .Q (signal_6477) ) ;
    buf_clk cell_4508 ( .C (clk), .D (plaintext_s1[70]), .Q (signal_6479) ) ;
    buf_clk cell_4510 ( .C (clk), .D (plaintext_s0[71]), .Q (signal_6481) ) ;
    buf_clk cell_4512 ( .C (clk), .D (plaintext_s1[71]), .Q (signal_6483) ) ;
    buf_clk cell_4514 ( .C (clk), .D (plaintext_s0[72]), .Q (signal_6485) ) ;
    buf_clk cell_4516 ( .C (clk), .D (plaintext_s1[72]), .Q (signal_6487) ) ;
    buf_clk cell_4518 ( .C (clk), .D (plaintext_s0[73]), .Q (signal_6489) ) ;
    buf_clk cell_4520 ( .C (clk), .D (plaintext_s1[73]), .Q (signal_6491) ) ;
    buf_clk cell_4522 ( .C (clk), .D (plaintext_s0[74]), .Q (signal_6493) ) ;
    buf_clk cell_4524 ( .C (clk), .D (plaintext_s1[74]), .Q (signal_6495) ) ;
    buf_clk cell_4526 ( .C (clk), .D (plaintext_s0[75]), .Q (signal_6497) ) ;
    buf_clk cell_4528 ( .C (clk), .D (plaintext_s1[75]), .Q (signal_6499) ) ;
    buf_clk cell_4530 ( .C (clk), .D (plaintext_s0[76]), .Q (signal_6501) ) ;
    buf_clk cell_4532 ( .C (clk), .D (plaintext_s1[76]), .Q (signal_6503) ) ;
    buf_clk cell_4534 ( .C (clk), .D (plaintext_s0[77]), .Q (signal_6505) ) ;
    buf_clk cell_4536 ( .C (clk), .D (plaintext_s1[77]), .Q (signal_6507) ) ;
    buf_clk cell_4538 ( .C (clk), .D (plaintext_s0[78]), .Q (signal_6509) ) ;
    buf_clk cell_4540 ( .C (clk), .D (plaintext_s1[78]), .Q (signal_6511) ) ;
    buf_clk cell_4542 ( .C (clk), .D (plaintext_s0[79]), .Q (signal_6513) ) ;
    buf_clk cell_4544 ( .C (clk), .D (plaintext_s1[79]), .Q (signal_6515) ) ;
    buf_clk cell_4546 ( .C (clk), .D (plaintext_s0[80]), .Q (signal_6517) ) ;
    buf_clk cell_4548 ( .C (clk), .D (plaintext_s1[80]), .Q (signal_6519) ) ;
    buf_clk cell_4550 ( .C (clk), .D (plaintext_s0[81]), .Q (signal_6521) ) ;
    buf_clk cell_4552 ( .C (clk), .D (plaintext_s1[81]), .Q (signal_6523) ) ;
    buf_clk cell_4554 ( .C (clk), .D (plaintext_s0[82]), .Q (signal_6525) ) ;
    buf_clk cell_4556 ( .C (clk), .D (plaintext_s1[82]), .Q (signal_6527) ) ;
    buf_clk cell_4558 ( .C (clk), .D (plaintext_s0[83]), .Q (signal_6529) ) ;
    buf_clk cell_4560 ( .C (clk), .D (plaintext_s1[83]), .Q (signal_6531) ) ;
    buf_clk cell_4562 ( .C (clk), .D (plaintext_s0[84]), .Q (signal_6533) ) ;
    buf_clk cell_4564 ( .C (clk), .D (plaintext_s1[84]), .Q (signal_6535) ) ;
    buf_clk cell_4566 ( .C (clk), .D (plaintext_s0[85]), .Q (signal_6537) ) ;
    buf_clk cell_4568 ( .C (clk), .D (plaintext_s1[85]), .Q (signal_6539) ) ;
    buf_clk cell_4570 ( .C (clk), .D (plaintext_s0[86]), .Q (signal_6541) ) ;
    buf_clk cell_4572 ( .C (clk), .D (plaintext_s1[86]), .Q (signal_6543) ) ;
    buf_clk cell_4574 ( .C (clk), .D (plaintext_s0[87]), .Q (signal_6545) ) ;
    buf_clk cell_4576 ( .C (clk), .D (plaintext_s1[87]), .Q (signal_6547) ) ;
    buf_clk cell_4578 ( .C (clk), .D (plaintext_s0[88]), .Q (signal_6549) ) ;
    buf_clk cell_4580 ( .C (clk), .D (plaintext_s1[88]), .Q (signal_6551) ) ;
    buf_clk cell_4582 ( .C (clk), .D (plaintext_s0[89]), .Q (signal_6553) ) ;
    buf_clk cell_4584 ( .C (clk), .D (plaintext_s1[89]), .Q (signal_6555) ) ;
    buf_clk cell_4586 ( .C (clk), .D (plaintext_s0[90]), .Q (signal_6557) ) ;
    buf_clk cell_4588 ( .C (clk), .D (plaintext_s1[90]), .Q (signal_6559) ) ;
    buf_clk cell_4590 ( .C (clk), .D (plaintext_s0[91]), .Q (signal_6561) ) ;
    buf_clk cell_4592 ( .C (clk), .D (plaintext_s1[91]), .Q (signal_6563) ) ;
    buf_clk cell_4594 ( .C (clk), .D (plaintext_s0[92]), .Q (signal_6565) ) ;
    buf_clk cell_4596 ( .C (clk), .D (plaintext_s1[92]), .Q (signal_6567) ) ;
    buf_clk cell_4598 ( .C (clk), .D (plaintext_s0[93]), .Q (signal_6569) ) ;
    buf_clk cell_4600 ( .C (clk), .D (plaintext_s1[93]), .Q (signal_6571) ) ;
    buf_clk cell_4602 ( .C (clk), .D (plaintext_s0[94]), .Q (signal_6573) ) ;
    buf_clk cell_4604 ( .C (clk), .D (plaintext_s1[94]), .Q (signal_6575) ) ;
    buf_clk cell_4606 ( .C (clk), .D (plaintext_s0[95]), .Q (signal_6577) ) ;
    buf_clk cell_4608 ( .C (clk), .D (plaintext_s1[95]), .Q (signal_6579) ) ;
    buf_clk cell_4610 ( .C (clk), .D (plaintext_s0[96]), .Q (signal_6581) ) ;
    buf_clk cell_4612 ( .C (clk), .D (plaintext_s1[96]), .Q (signal_6583) ) ;
    buf_clk cell_4614 ( .C (clk), .D (plaintext_s0[97]), .Q (signal_6585) ) ;
    buf_clk cell_4616 ( .C (clk), .D (plaintext_s1[97]), .Q (signal_6587) ) ;
    buf_clk cell_4618 ( .C (clk), .D (plaintext_s0[98]), .Q (signal_6589) ) ;
    buf_clk cell_4620 ( .C (clk), .D (plaintext_s1[98]), .Q (signal_6591) ) ;
    buf_clk cell_4622 ( .C (clk), .D (plaintext_s0[99]), .Q (signal_6593) ) ;
    buf_clk cell_4624 ( .C (clk), .D (plaintext_s1[99]), .Q (signal_6595) ) ;
    buf_clk cell_4626 ( .C (clk), .D (plaintext_s0[100]), .Q (signal_6597) ) ;
    buf_clk cell_4628 ( .C (clk), .D (plaintext_s1[100]), .Q (signal_6599) ) ;
    buf_clk cell_4630 ( .C (clk), .D (plaintext_s0[101]), .Q (signal_6601) ) ;
    buf_clk cell_4632 ( .C (clk), .D (plaintext_s1[101]), .Q (signal_6603) ) ;
    buf_clk cell_4634 ( .C (clk), .D (plaintext_s0[102]), .Q (signal_6605) ) ;
    buf_clk cell_4636 ( .C (clk), .D (plaintext_s1[102]), .Q (signal_6607) ) ;
    buf_clk cell_4638 ( .C (clk), .D (plaintext_s0[103]), .Q (signal_6609) ) ;
    buf_clk cell_4640 ( .C (clk), .D (plaintext_s1[103]), .Q (signal_6611) ) ;
    buf_clk cell_4642 ( .C (clk), .D (plaintext_s0[104]), .Q (signal_6613) ) ;
    buf_clk cell_4644 ( .C (clk), .D (plaintext_s1[104]), .Q (signal_6615) ) ;
    buf_clk cell_4646 ( .C (clk), .D (plaintext_s0[105]), .Q (signal_6617) ) ;
    buf_clk cell_4648 ( .C (clk), .D (plaintext_s1[105]), .Q (signal_6619) ) ;
    buf_clk cell_4650 ( .C (clk), .D (plaintext_s0[106]), .Q (signal_6621) ) ;
    buf_clk cell_4652 ( .C (clk), .D (plaintext_s1[106]), .Q (signal_6623) ) ;
    buf_clk cell_4654 ( .C (clk), .D (plaintext_s0[107]), .Q (signal_6625) ) ;
    buf_clk cell_4656 ( .C (clk), .D (plaintext_s1[107]), .Q (signal_6627) ) ;
    buf_clk cell_4658 ( .C (clk), .D (plaintext_s0[108]), .Q (signal_6629) ) ;
    buf_clk cell_4660 ( .C (clk), .D (plaintext_s1[108]), .Q (signal_6631) ) ;
    buf_clk cell_4662 ( .C (clk), .D (plaintext_s0[109]), .Q (signal_6633) ) ;
    buf_clk cell_4664 ( .C (clk), .D (plaintext_s1[109]), .Q (signal_6635) ) ;
    buf_clk cell_4666 ( .C (clk), .D (plaintext_s0[110]), .Q (signal_6637) ) ;
    buf_clk cell_4668 ( .C (clk), .D (plaintext_s1[110]), .Q (signal_6639) ) ;
    buf_clk cell_4670 ( .C (clk), .D (plaintext_s0[111]), .Q (signal_6641) ) ;
    buf_clk cell_4672 ( .C (clk), .D (plaintext_s1[111]), .Q (signal_6643) ) ;
    buf_clk cell_4674 ( .C (clk), .D (plaintext_s0[112]), .Q (signal_6645) ) ;
    buf_clk cell_4676 ( .C (clk), .D (plaintext_s1[112]), .Q (signal_6647) ) ;
    buf_clk cell_4678 ( .C (clk), .D (plaintext_s0[113]), .Q (signal_6649) ) ;
    buf_clk cell_4680 ( .C (clk), .D (plaintext_s1[113]), .Q (signal_6651) ) ;
    buf_clk cell_4682 ( .C (clk), .D (plaintext_s0[114]), .Q (signal_6653) ) ;
    buf_clk cell_4684 ( .C (clk), .D (plaintext_s1[114]), .Q (signal_6655) ) ;
    buf_clk cell_4686 ( .C (clk), .D (plaintext_s0[115]), .Q (signal_6657) ) ;
    buf_clk cell_4688 ( .C (clk), .D (plaintext_s1[115]), .Q (signal_6659) ) ;
    buf_clk cell_4690 ( .C (clk), .D (plaintext_s0[116]), .Q (signal_6661) ) ;
    buf_clk cell_4692 ( .C (clk), .D (plaintext_s1[116]), .Q (signal_6663) ) ;
    buf_clk cell_4694 ( .C (clk), .D (plaintext_s0[117]), .Q (signal_6665) ) ;
    buf_clk cell_4696 ( .C (clk), .D (plaintext_s1[117]), .Q (signal_6667) ) ;
    buf_clk cell_4698 ( .C (clk), .D (plaintext_s0[118]), .Q (signal_6669) ) ;
    buf_clk cell_4700 ( .C (clk), .D (plaintext_s1[118]), .Q (signal_6671) ) ;
    buf_clk cell_4702 ( .C (clk), .D (plaintext_s0[119]), .Q (signal_6673) ) ;
    buf_clk cell_4704 ( .C (clk), .D (plaintext_s1[119]), .Q (signal_6675) ) ;
    buf_clk cell_4706 ( .C (clk), .D (plaintext_s0[120]), .Q (signal_6677) ) ;
    buf_clk cell_4708 ( .C (clk), .D (plaintext_s1[120]), .Q (signal_6679) ) ;
    buf_clk cell_4710 ( .C (clk), .D (plaintext_s0[121]), .Q (signal_6681) ) ;
    buf_clk cell_4712 ( .C (clk), .D (plaintext_s1[121]), .Q (signal_6683) ) ;
    buf_clk cell_4714 ( .C (clk), .D (plaintext_s0[122]), .Q (signal_6685) ) ;
    buf_clk cell_4716 ( .C (clk), .D (plaintext_s1[122]), .Q (signal_6687) ) ;
    buf_clk cell_4718 ( .C (clk), .D (plaintext_s0[123]), .Q (signal_6689) ) ;
    buf_clk cell_4720 ( .C (clk), .D (plaintext_s1[123]), .Q (signal_6691) ) ;
    buf_clk cell_4722 ( .C (clk), .D (plaintext_s0[124]), .Q (signal_6693) ) ;
    buf_clk cell_4724 ( .C (clk), .D (plaintext_s1[124]), .Q (signal_6695) ) ;
    buf_clk cell_4726 ( .C (clk), .D (plaintext_s0[125]), .Q (signal_6697) ) ;
    buf_clk cell_4728 ( .C (clk), .D (plaintext_s1[125]), .Q (signal_6699) ) ;
    buf_clk cell_4730 ( .C (clk), .D (plaintext_s0[126]), .Q (signal_6701) ) ;
    buf_clk cell_4732 ( .C (clk), .D (plaintext_s1[126]), .Q (signal_6703) ) ;
    buf_clk cell_4734 ( .C (clk), .D (plaintext_s0[127]), .Q (signal_6705) ) ;
    buf_clk cell_4736 ( .C (clk), .D (plaintext_s1[127]), .Q (signal_6707) ) ;
    buf_clk cell_4738 ( .C (clk), .D (key_s0[0]), .Q (signal_6709) ) ;
    buf_clk cell_4740 ( .C (clk), .D (key_s1[0]), .Q (signal_6711) ) ;
    buf_clk cell_4742 ( .C (clk), .D (key_s0[1]), .Q (signal_6713) ) ;
    buf_clk cell_4744 ( .C (clk), .D (key_s1[1]), .Q (signal_6715) ) ;
    buf_clk cell_4746 ( .C (clk), .D (key_s0[2]), .Q (signal_6717) ) ;
    buf_clk cell_4748 ( .C (clk), .D (key_s1[2]), .Q (signal_6719) ) ;
    buf_clk cell_4750 ( .C (clk), .D (key_s0[3]), .Q (signal_6721) ) ;
    buf_clk cell_4752 ( .C (clk), .D (key_s1[3]), .Q (signal_6723) ) ;
    buf_clk cell_4754 ( .C (clk), .D (key_s0[4]), .Q (signal_6725) ) ;
    buf_clk cell_4756 ( .C (clk), .D (key_s1[4]), .Q (signal_6727) ) ;
    buf_clk cell_4758 ( .C (clk), .D (key_s0[5]), .Q (signal_6729) ) ;
    buf_clk cell_4760 ( .C (clk), .D (key_s1[5]), .Q (signal_6731) ) ;
    buf_clk cell_4762 ( .C (clk), .D (key_s0[6]), .Q (signal_6733) ) ;
    buf_clk cell_4764 ( .C (clk), .D (key_s1[6]), .Q (signal_6735) ) ;
    buf_clk cell_4766 ( .C (clk), .D (key_s0[7]), .Q (signal_6737) ) ;
    buf_clk cell_4768 ( .C (clk), .D (key_s1[7]), .Q (signal_6739) ) ;
    buf_clk cell_4770 ( .C (clk), .D (key_s0[8]), .Q (signal_6741) ) ;
    buf_clk cell_4772 ( .C (clk), .D (key_s1[8]), .Q (signal_6743) ) ;
    buf_clk cell_4774 ( .C (clk), .D (key_s0[9]), .Q (signal_6745) ) ;
    buf_clk cell_4776 ( .C (clk), .D (key_s1[9]), .Q (signal_6747) ) ;
    buf_clk cell_4778 ( .C (clk), .D (key_s0[10]), .Q (signal_6749) ) ;
    buf_clk cell_4780 ( .C (clk), .D (key_s1[10]), .Q (signal_6751) ) ;
    buf_clk cell_4782 ( .C (clk), .D (key_s0[11]), .Q (signal_6753) ) ;
    buf_clk cell_4784 ( .C (clk), .D (key_s1[11]), .Q (signal_6755) ) ;
    buf_clk cell_4786 ( .C (clk), .D (key_s0[12]), .Q (signal_6757) ) ;
    buf_clk cell_4788 ( .C (clk), .D (key_s1[12]), .Q (signal_6759) ) ;
    buf_clk cell_4790 ( .C (clk), .D (key_s0[13]), .Q (signal_6761) ) ;
    buf_clk cell_4792 ( .C (clk), .D (key_s1[13]), .Q (signal_6763) ) ;
    buf_clk cell_4794 ( .C (clk), .D (key_s0[14]), .Q (signal_6765) ) ;
    buf_clk cell_4796 ( .C (clk), .D (key_s1[14]), .Q (signal_6767) ) ;
    buf_clk cell_4798 ( .C (clk), .D (key_s0[15]), .Q (signal_6769) ) ;
    buf_clk cell_4800 ( .C (clk), .D (key_s1[15]), .Q (signal_6771) ) ;
    buf_clk cell_4802 ( .C (clk), .D (key_s0[16]), .Q (signal_6773) ) ;
    buf_clk cell_4804 ( .C (clk), .D (key_s1[16]), .Q (signal_6775) ) ;
    buf_clk cell_4806 ( .C (clk), .D (key_s0[17]), .Q (signal_6777) ) ;
    buf_clk cell_4808 ( .C (clk), .D (key_s1[17]), .Q (signal_6779) ) ;
    buf_clk cell_4810 ( .C (clk), .D (key_s0[18]), .Q (signal_6781) ) ;
    buf_clk cell_4812 ( .C (clk), .D (key_s1[18]), .Q (signal_6783) ) ;
    buf_clk cell_4814 ( .C (clk), .D (key_s0[19]), .Q (signal_6785) ) ;
    buf_clk cell_4816 ( .C (clk), .D (key_s1[19]), .Q (signal_6787) ) ;
    buf_clk cell_4818 ( .C (clk), .D (key_s0[20]), .Q (signal_6789) ) ;
    buf_clk cell_4820 ( .C (clk), .D (key_s1[20]), .Q (signal_6791) ) ;
    buf_clk cell_4822 ( .C (clk), .D (key_s0[21]), .Q (signal_6793) ) ;
    buf_clk cell_4824 ( .C (clk), .D (key_s1[21]), .Q (signal_6795) ) ;
    buf_clk cell_4826 ( .C (clk), .D (key_s0[22]), .Q (signal_6797) ) ;
    buf_clk cell_4828 ( .C (clk), .D (key_s1[22]), .Q (signal_6799) ) ;
    buf_clk cell_4830 ( .C (clk), .D (key_s0[23]), .Q (signal_6801) ) ;
    buf_clk cell_4832 ( .C (clk), .D (key_s1[23]), .Q (signal_6803) ) ;
    buf_clk cell_4834 ( .C (clk), .D (key_s0[24]), .Q (signal_6805) ) ;
    buf_clk cell_4836 ( .C (clk), .D (key_s1[24]), .Q (signal_6807) ) ;
    buf_clk cell_4838 ( .C (clk), .D (key_s0[25]), .Q (signal_6809) ) ;
    buf_clk cell_4840 ( .C (clk), .D (key_s1[25]), .Q (signal_6811) ) ;
    buf_clk cell_4842 ( .C (clk), .D (key_s0[26]), .Q (signal_6813) ) ;
    buf_clk cell_4844 ( .C (clk), .D (key_s1[26]), .Q (signal_6815) ) ;
    buf_clk cell_4846 ( .C (clk), .D (key_s0[27]), .Q (signal_6817) ) ;
    buf_clk cell_4848 ( .C (clk), .D (key_s1[27]), .Q (signal_6819) ) ;
    buf_clk cell_4850 ( .C (clk), .D (key_s0[28]), .Q (signal_6821) ) ;
    buf_clk cell_4852 ( .C (clk), .D (key_s1[28]), .Q (signal_6823) ) ;
    buf_clk cell_4854 ( .C (clk), .D (key_s0[29]), .Q (signal_6825) ) ;
    buf_clk cell_4856 ( .C (clk), .D (key_s1[29]), .Q (signal_6827) ) ;
    buf_clk cell_4858 ( .C (clk), .D (key_s0[30]), .Q (signal_6829) ) ;
    buf_clk cell_4860 ( .C (clk), .D (key_s1[30]), .Q (signal_6831) ) ;
    buf_clk cell_4862 ( .C (clk), .D (key_s0[31]), .Q (signal_6833) ) ;
    buf_clk cell_4864 ( .C (clk), .D (key_s1[31]), .Q (signal_6835) ) ;
    buf_clk cell_4866 ( .C (clk), .D (key_s0[32]), .Q (signal_6837) ) ;
    buf_clk cell_4868 ( .C (clk), .D (key_s1[32]), .Q (signal_6839) ) ;
    buf_clk cell_4870 ( .C (clk), .D (key_s0[33]), .Q (signal_6841) ) ;
    buf_clk cell_4872 ( .C (clk), .D (key_s1[33]), .Q (signal_6843) ) ;
    buf_clk cell_4874 ( .C (clk), .D (key_s0[34]), .Q (signal_6845) ) ;
    buf_clk cell_4876 ( .C (clk), .D (key_s1[34]), .Q (signal_6847) ) ;
    buf_clk cell_4878 ( .C (clk), .D (key_s0[35]), .Q (signal_6849) ) ;
    buf_clk cell_4880 ( .C (clk), .D (key_s1[35]), .Q (signal_6851) ) ;
    buf_clk cell_4882 ( .C (clk), .D (key_s0[36]), .Q (signal_6853) ) ;
    buf_clk cell_4884 ( .C (clk), .D (key_s1[36]), .Q (signal_6855) ) ;
    buf_clk cell_4886 ( .C (clk), .D (key_s0[37]), .Q (signal_6857) ) ;
    buf_clk cell_4888 ( .C (clk), .D (key_s1[37]), .Q (signal_6859) ) ;
    buf_clk cell_4890 ( .C (clk), .D (key_s0[38]), .Q (signal_6861) ) ;
    buf_clk cell_4892 ( .C (clk), .D (key_s1[38]), .Q (signal_6863) ) ;
    buf_clk cell_4894 ( .C (clk), .D (key_s0[39]), .Q (signal_6865) ) ;
    buf_clk cell_4896 ( .C (clk), .D (key_s1[39]), .Q (signal_6867) ) ;
    buf_clk cell_4898 ( .C (clk), .D (key_s0[40]), .Q (signal_6869) ) ;
    buf_clk cell_4900 ( .C (clk), .D (key_s1[40]), .Q (signal_6871) ) ;
    buf_clk cell_4902 ( .C (clk), .D (key_s0[41]), .Q (signal_6873) ) ;
    buf_clk cell_4904 ( .C (clk), .D (key_s1[41]), .Q (signal_6875) ) ;
    buf_clk cell_4906 ( .C (clk), .D (key_s0[42]), .Q (signal_6877) ) ;
    buf_clk cell_4908 ( .C (clk), .D (key_s1[42]), .Q (signal_6879) ) ;
    buf_clk cell_4910 ( .C (clk), .D (key_s0[43]), .Q (signal_6881) ) ;
    buf_clk cell_4912 ( .C (clk), .D (key_s1[43]), .Q (signal_6883) ) ;
    buf_clk cell_4914 ( .C (clk), .D (key_s0[44]), .Q (signal_6885) ) ;
    buf_clk cell_4916 ( .C (clk), .D (key_s1[44]), .Q (signal_6887) ) ;
    buf_clk cell_4918 ( .C (clk), .D (key_s0[45]), .Q (signal_6889) ) ;
    buf_clk cell_4920 ( .C (clk), .D (key_s1[45]), .Q (signal_6891) ) ;
    buf_clk cell_4922 ( .C (clk), .D (key_s0[46]), .Q (signal_6893) ) ;
    buf_clk cell_4924 ( .C (clk), .D (key_s1[46]), .Q (signal_6895) ) ;
    buf_clk cell_4926 ( .C (clk), .D (key_s0[47]), .Q (signal_6897) ) ;
    buf_clk cell_4928 ( .C (clk), .D (key_s1[47]), .Q (signal_6899) ) ;
    buf_clk cell_4930 ( .C (clk), .D (key_s0[48]), .Q (signal_6901) ) ;
    buf_clk cell_4932 ( .C (clk), .D (key_s1[48]), .Q (signal_6903) ) ;
    buf_clk cell_4934 ( .C (clk), .D (key_s0[49]), .Q (signal_6905) ) ;
    buf_clk cell_4936 ( .C (clk), .D (key_s1[49]), .Q (signal_6907) ) ;
    buf_clk cell_4938 ( .C (clk), .D (key_s0[50]), .Q (signal_6909) ) ;
    buf_clk cell_4940 ( .C (clk), .D (key_s1[50]), .Q (signal_6911) ) ;
    buf_clk cell_4942 ( .C (clk), .D (key_s0[51]), .Q (signal_6913) ) ;
    buf_clk cell_4944 ( .C (clk), .D (key_s1[51]), .Q (signal_6915) ) ;
    buf_clk cell_4946 ( .C (clk), .D (key_s0[52]), .Q (signal_6917) ) ;
    buf_clk cell_4948 ( .C (clk), .D (key_s1[52]), .Q (signal_6919) ) ;
    buf_clk cell_4950 ( .C (clk), .D (key_s0[53]), .Q (signal_6921) ) ;
    buf_clk cell_4952 ( .C (clk), .D (key_s1[53]), .Q (signal_6923) ) ;
    buf_clk cell_4954 ( .C (clk), .D (key_s0[54]), .Q (signal_6925) ) ;
    buf_clk cell_4956 ( .C (clk), .D (key_s1[54]), .Q (signal_6927) ) ;
    buf_clk cell_4958 ( .C (clk), .D (key_s0[55]), .Q (signal_6929) ) ;
    buf_clk cell_4960 ( .C (clk), .D (key_s1[55]), .Q (signal_6931) ) ;
    buf_clk cell_4962 ( .C (clk), .D (key_s0[56]), .Q (signal_6933) ) ;
    buf_clk cell_4964 ( .C (clk), .D (key_s1[56]), .Q (signal_6935) ) ;
    buf_clk cell_4966 ( .C (clk), .D (key_s0[57]), .Q (signal_6937) ) ;
    buf_clk cell_4968 ( .C (clk), .D (key_s1[57]), .Q (signal_6939) ) ;
    buf_clk cell_4970 ( .C (clk), .D (key_s0[58]), .Q (signal_6941) ) ;
    buf_clk cell_4972 ( .C (clk), .D (key_s1[58]), .Q (signal_6943) ) ;
    buf_clk cell_4974 ( .C (clk), .D (key_s0[59]), .Q (signal_6945) ) ;
    buf_clk cell_4976 ( .C (clk), .D (key_s1[59]), .Q (signal_6947) ) ;
    buf_clk cell_4978 ( .C (clk), .D (key_s0[60]), .Q (signal_6949) ) ;
    buf_clk cell_4980 ( .C (clk), .D (key_s1[60]), .Q (signal_6951) ) ;
    buf_clk cell_4982 ( .C (clk), .D (key_s0[61]), .Q (signal_6953) ) ;
    buf_clk cell_4984 ( .C (clk), .D (key_s1[61]), .Q (signal_6955) ) ;
    buf_clk cell_4986 ( .C (clk), .D (key_s0[62]), .Q (signal_6957) ) ;
    buf_clk cell_4988 ( .C (clk), .D (key_s1[62]), .Q (signal_6959) ) ;
    buf_clk cell_4990 ( .C (clk), .D (key_s0[63]), .Q (signal_6961) ) ;
    buf_clk cell_4992 ( .C (clk), .D (key_s1[63]), .Q (signal_6963) ) ;
    buf_clk cell_4994 ( .C (clk), .D (key_s0[64]), .Q (signal_6965) ) ;
    buf_clk cell_4996 ( .C (clk), .D (key_s1[64]), .Q (signal_6967) ) ;
    buf_clk cell_4998 ( .C (clk), .D (key_s0[65]), .Q (signal_6969) ) ;
    buf_clk cell_5000 ( .C (clk), .D (key_s1[65]), .Q (signal_6971) ) ;
    buf_clk cell_5002 ( .C (clk), .D (key_s0[66]), .Q (signal_6973) ) ;
    buf_clk cell_5004 ( .C (clk), .D (key_s1[66]), .Q (signal_6975) ) ;
    buf_clk cell_5006 ( .C (clk), .D (key_s0[67]), .Q (signal_6977) ) ;
    buf_clk cell_5008 ( .C (clk), .D (key_s1[67]), .Q (signal_6979) ) ;
    buf_clk cell_5010 ( .C (clk), .D (key_s0[68]), .Q (signal_6981) ) ;
    buf_clk cell_5012 ( .C (clk), .D (key_s1[68]), .Q (signal_6983) ) ;
    buf_clk cell_5014 ( .C (clk), .D (key_s0[69]), .Q (signal_6985) ) ;
    buf_clk cell_5016 ( .C (clk), .D (key_s1[69]), .Q (signal_6987) ) ;
    buf_clk cell_5018 ( .C (clk), .D (key_s0[70]), .Q (signal_6989) ) ;
    buf_clk cell_5020 ( .C (clk), .D (key_s1[70]), .Q (signal_6991) ) ;
    buf_clk cell_5022 ( .C (clk), .D (key_s0[71]), .Q (signal_6993) ) ;
    buf_clk cell_5024 ( .C (clk), .D (key_s1[71]), .Q (signal_6995) ) ;
    buf_clk cell_5026 ( .C (clk), .D (key_s0[72]), .Q (signal_6997) ) ;
    buf_clk cell_5028 ( .C (clk), .D (key_s1[72]), .Q (signal_6999) ) ;
    buf_clk cell_5030 ( .C (clk), .D (key_s0[73]), .Q (signal_7001) ) ;
    buf_clk cell_5032 ( .C (clk), .D (key_s1[73]), .Q (signal_7003) ) ;
    buf_clk cell_5034 ( .C (clk), .D (key_s0[74]), .Q (signal_7005) ) ;
    buf_clk cell_5036 ( .C (clk), .D (key_s1[74]), .Q (signal_7007) ) ;
    buf_clk cell_5038 ( .C (clk), .D (key_s0[75]), .Q (signal_7009) ) ;
    buf_clk cell_5040 ( .C (clk), .D (key_s1[75]), .Q (signal_7011) ) ;
    buf_clk cell_5042 ( .C (clk), .D (key_s0[76]), .Q (signal_7013) ) ;
    buf_clk cell_5044 ( .C (clk), .D (key_s1[76]), .Q (signal_7015) ) ;
    buf_clk cell_5046 ( .C (clk), .D (key_s0[77]), .Q (signal_7017) ) ;
    buf_clk cell_5048 ( .C (clk), .D (key_s1[77]), .Q (signal_7019) ) ;
    buf_clk cell_5050 ( .C (clk), .D (key_s0[78]), .Q (signal_7021) ) ;
    buf_clk cell_5052 ( .C (clk), .D (key_s1[78]), .Q (signal_7023) ) ;
    buf_clk cell_5054 ( .C (clk), .D (key_s0[79]), .Q (signal_7025) ) ;
    buf_clk cell_5056 ( .C (clk), .D (key_s1[79]), .Q (signal_7027) ) ;
    buf_clk cell_5058 ( .C (clk), .D (key_s0[80]), .Q (signal_7029) ) ;
    buf_clk cell_5060 ( .C (clk), .D (key_s1[80]), .Q (signal_7031) ) ;
    buf_clk cell_5062 ( .C (clk), .D (key_s0[81]), .Q (signal_7033) ) ;
    buf_clk cell_5064 ( .C (clk), .D (key_s1[81]), .Q (signal_7035) ) ;
    buf_clk cell_5066 ( .C (clk), .D (key_s0[82]), .Q (signal_7037) ) ;
    buf_clk cell_5068 ( .C (clk), .D (key_s1[82]), .Q (signal_7039) ) ;
    buf_clk cell_5070 ( .C (clk), .D (key_s0[83]), .Q (signal_7041) ) ;
    buf_clk cell_5072 ( .C (clk), .D (key_s1[83]), .Q (signal_7043) ) ;
    buf_clk cell_5074 ( .C (clk), .D (key_s0[84]), .Q (signal_7045) ) ;
    buf_clk cell_5076 ( .C (clk), .D (key_s1[84]), .Q (signal_7047) ) ;
    buf_clk cell_5078 ( .C (clk), .D (key_s0[85]), .Q (signal_7049) ) ;
    buf_clk cell_5080 ( .C (clk), .D (key_s1[85]), .Q (signal_7051) ) ;
    buf_clk cell_5082 ( .C (clk), .D (key_s0[86]), .Q (signal_7053) ) ;
    buf_clk cell_5084 ( .C (clk), .D (key_s1[86]), .Q (signal_7055) ) ;
    buf_clk cell_5086 ( .C (clk), .D (key_s0[87]), .Q (signal_7057) ) ;
    buf_clk cell_5088 ( .C (clk), .D (key_s1[87]), .Q (signal_7059) ) ;
    buf_clk cell_5090 ( .C (clk), .D (key_s0[88]), .Q (signal_7061) ) ;
    buf_clk cell_5092 ( .C (clk), .D (key_s1[88]), .Q (signal_7063) ) ;
    buf_clk cell_5094 ( .C (clk), .D (key_s0[89]), .Q (signal_7065) ) ;
    buf_clk cell_5096 ( .C (clk), .D (key_s1[89]), .Q (signal_7067) ) ;
    buf_clk cell_5098 ( .C (clk), .D (key_s0[90]), .Q (signal_7069) ) ;
    buf_clk cell_5100 ( .C (clk), .D (key_s1[90]), .Q (signal_7071) ) ;
    buf_clk cell_5102 ( .C (clk), .D (key_s0[91]), .Q (signal_7073) ) ;
    buf_clk cell_5104 ( .C (clk), .D (key_s1[91]), .Q (signal_7075) ) ;
    buf_clk cell_5106 ( .C (clk), .D (key_s0[92]), .Q (signal_7077) ) ;
    buf_clk cell_5108 ( .C (clk), .D (key_s1[92]), .Q (signal_7079) ) ;
    buf_clk cell_5110 ( .C (clk), .D (key_s0[93]), .Q (signal_7081) ) ;
    buf_clk cell_5112 ( .C (clk), .D (key_s1[93]), .Q (signal_7083) ) ;
    buf_clk cell_5114 ( .C (clk), .D (key_s0[94]), .Q (signal_7085) ) ;
    buf_clk cell_5116 ( .C (clk), .D (key_s1[94]), .Q (signal_7087) ) ;
    buf_clk cell_5118 ( .C (clk), .D (key_s0[95]), .Q (signal_7089) ) ;
    buf_clk cell_5120 ( .C (clk), .D (key_s1[95]), .Q (signal_7091) ) ;
    buf_clk cell_5122 ( .C (clk), .D (key_s0[96]), .Q (signal_7093) ) ;
    buf_clk cell_5124 ( .C (clk), .D (key_s1[96]), .Q (signal_7095) ) ;
    buf_clk cell_5126 ( .C (clk), .D (key_s0[97]), .Q (signal_7097) ) ;
    buf_clk cell_5128 ( .C (clk), .D (key_s1[97]), .Q (signal_7099) ) ;
    buf_clk cell_5130 ( .C (clk), .D (key_s0[98]), .Q (signal_7101) ) ;
    buf_clk cell_5132 ( .C (clk), .D (key_s1[98]), .Q (signal_7103) ) ;
    buf_clk cell_5134 ( .C (clk), .D (key_s0[99]), .Q (signal_7105) ) ;
    buf_clk cell_5136 ( .C (clk), .D (key_s1[99]), .Q (signal_7107) ) ;
    buf_clk cell_5138 ( .C (clk), .D (key_s0[100]), .Q (signal_7109) ) ;
    buf_clk cell_5140 ( .C (clk), .D (key_s1[100]), .Q (signal_7111) ) ;
    buf_clk cell_5142 ( .C (clk), .D (key_s0[101]), .Q (signal_7113) ) ;
    buf_clk cell_5144 ( .C (clk), .D (key_s1[101]), .Q (signal_7115) ) ;
    buf_clk cell_5146 ( .C (clk), .D (key_s0[102]), .Q (signal_7117) ) ;
    buf_clk cell_5148 ( .C (clk), .D (key_s1[102]), .Q (signal_7119) ) ;
    buf_clk cell_5150 ( .C (clk), .D (key_s0[103]), .Q (signal_7121) ) ;
    buf_clk cell_5152 ( .C (clk), .D (key_s1[103]), .Q (signal_7123) ) ;
    buf_clk cell_5154 ( .C (clk), .D (key_s0[104]), .Q (signal_7125) ) ;
    buf_clk cell_5156 ( .C (clk), .D (key_s1[104]), .Q (signal_7127) ) ;
    buf_clk cell_5158 ( .C (clk), .D (key_s0[105]), .Q (signal_7129) ) ;
    buf_clk cell_5160 ( .C (clk), .D (key_s1[105]), .Q (signal_7131) ) ;
    buf_clk cell_5162 ( .C (clk), .D (key_s0[106]), .Q (signal_7133) ) ;
    buf_clk cell_5164 ( .C (clk), .D (key_s1[106]), .Q (signal_7135) ) ;
    buf_clk cell_5166 ( .C (clk), .D (key_s0[107]), .Q (signal_7137) ) ;
    buf_clk cell_5168 ( .C (clk), .D (key_s1[107]), .Q (signal_7139) ) ;
    buf_clk cell_5170 ( .C (clk), .D (key_s0[108]), .Q (signal_7141) ) ;
    buf_clk cell_5172 ( .C (clk), .D (key_s1[108]), .Q (signal_7143) ) ;
    buf_clk cell_5174 ( .C (clk), .D (key_s0[109]), .Q (signal_7145) ) ;
    buf_clk cell_5176 ( .C (clk), .D (key_s1[109]), .Q (signal_7147) ) ;
    buf_clk cell_5178 ( .C (clk), .D (key_s0[110]), .Q (signal_7149) ) ;
    buf_clk cell_5180 ( .C (clk), .D (key_s1[110]), .Q (signal_7151) ) ;
    buf_clk cell_5182 ( .C (clk), .D (key_s0[111]), .Q (signal_7153) ) ;
    buf_clk cell_5184 ( .C (clk), .D (key_s1[111]), .Q (signal_7155) ) ;
    buf_clk cell_5186 ( .C (clk), .D (key_s0[112]), .Q (signal_7157) ) ;
    buf_clk cell_5188 ( .C (clk), .D (key_s1[112]), .Q (signal_7159) ) ;
    buf_clk cell_5190 ( .C (clk), .D (key_s0[113]), .Q (signal_7161) ) ;
    buf_clk cell_5192 ( .C (clk), .D (key_s1[113]), .Q (signal_7163) ) ;
    buf_clk cell_5194 ( .C (clk), .D (key_s0[114]), .Q (signal_7165) ) ;
    buf_clk cell_5196 ( .C (clk), .D (key_s1[114]), .Q (signal_7167) ) ;
    buf_clk cell_5198 ( .C (clk), .D (key_s0[115]), .Q (signal_7169) ) ;
    buf_clk cell_5200 ( .C (clk), .D (key_s1[115]), .Q (signal_7171) ) ;
    buf_clk cell_5202 ( .C (clk), .D (key_s0[116]), .Q (signal_7173) ) ;
    buf_clk cell_5204 ( .C (clk), .D (key_s1[116]), .Q (signal_7175) ) ;
    buf_clk cell_5206 ( .C (clk), .D (key_s0[117]), .Q (signal_7177) ) ;
    buf_clk cell_5208 ( .C (clk), .D (key_s1[117]), .Q (signal_7179) ) ;
    buf_clk cell_5210 ( .C (clk), .D (key_s0[118]), .Q (signal_7181) ) ;
    buf_clk cell_5212 ( .C (clk), .D (key_s1[118]), .Q (signal_7183) ) ;
    buf_clk cell_5214 ( .C (clk), .D (key_s0[119]), .Q (signal_7185) ) ;
    buf_clk cell_5216 ( .C (clk), .D (key_s1[119]), .Q (signal_7187) ) ;
    buf_clk cell_5218 ( .C (clk), .D (key_s0[120]), .Q (signal_7189) ) ;
    buf_clk cell_5220 ( .C (clk), .D (key_s1[120]), .Q (signal_7191) ) ;
    buf_clk cell_5222 ( .C (clk), .D (key_s0[121]), .Q (signal_7193) ) ;
    buf_clk cell_5224 ( .C (clk), .D (key_s1[121]), .Q (signal_7195) ) ;
    buf_clk cell_5226 ( .C (clk), .D (key_s0[122]), .Q (signal_7197) ) ;
    buf_clk cell_5228 ( .C (clk), .D (key_s1[122]), .Q (signal_7199) ) ;
    buf_clk cell_5230 ( .C (clk), .D (key_s0[123]), .Q (signal_7201) ) ;
    buf_clk cell_5232 ( .C (clk), .D (key_s1[123]), .Q (signal_7203) ) ;
    buf_clk cell_5234 ( .C (clk), .D (key_s0[124]), .Q (signal_7205) ) ;
    buf_clk cell_5236 ( .C (clk), .D (key_s1[124]), .Q (signal_7207) ) ;
    buf_clk cell_5238 ( .C (clk), .D (key_s0[125]), .Q (signal_7209) ) ;
    buf_clk cell_5240 ( .C (clk), .D (key_s1[125]), .Q (signal_7211) ) ;
    buf_clk cell_5242 ( .C (clk), .D (key_s0[126]), .Q (signal_7213) ) ;
    buf_clk cell_5244 ( .C (clk), .D (key_s1[126]), .Q (signal_7215) ) ;
    buf_clk cell_5246 ( .C (clk), .D (key_s0[127]), .Q (signal_7217) ) ;
    buf_clk cell_5248 ( .C (clk), .D (key_s1[127]), .Q (signal_7219) ) ;
    buf_clk cell_5250 ( .C (clk), .D (signal_4369), .Q (signal_7221) ) ;
    buf_clk cell_5252 ( .C (clk), .D (signal_4931), .Q (signal_7223) ) ;
    buf_clk cell_5254 ( .C (clk), .D (signal_4370), .Q (signal_7225) ) ;
    buf_clk cell_5256 ( .C (clk), .D (signal_4898), .Q (signal_7227) ) ;
    buf_clk cell_5258 ( .C (clk), .D (signal_4371), .Q (signal_7229) ) ;
    buf_clk cell_5260 ( .C (clk), .D (signal_4865), .Q (signal_7231) ) ;
    buf_clk cell_5262 ( .C (clk), .D (signal_4372), .Q (signal_7233) ) ;
    buf_clk cell_5264 ( .C (clk), .D (signal_4832), .Q (signal_7235) ) ;
    buf_clk cell_5266 ( .C (clk), .D (signal_4373), .Q (signal_7237) ) ;
    buf_clk cell_5268 ( .C (clk), .D (signal_4799), .Q (signal_7239) ) ;
    buf_clk cell_5270 ( .C (clk), .D (signal_4374), .Q (signal_7241) ) ;
    buf_clk cell_5272 ( .C (clk), .D (signal_4766), .Q (signal_7243) ) ;
    buf_clk cell_5274 ( .C (clk), .D (signal_4337), .Q (signal_7245) ) ;
    buf_clk cell_5276 ( .C (clk), .D (signal_4739), .Q (signal_7247) ) ;
    buf_clk cell_5278 ( .C (clk), .D (signal_4305), .Q (signal_7249) ) ;
    buf_clk cell_5280 ( .C (clk), .D (signal_4844), .Q (signal_7251) ) ;
    buf_clk cell_5282 ( .C (clk), .D (signal_4338), .Q (signal_7253) ) ;
    buf_clk cell_5284 ( .C (clk), .D (signal_4736), .Q (signal_7255) ) ;
    buf_clk cell_5286 ( .C (clk), .D (signal_4306), .Q (signal_7257) ) ;
    buf_clk cell_5288 ( .C (clk), .D (signal_4841), .Q (signal_7259) ) ;
    buf_clk cell_5290 ( .C (clk), .D (signal_4375), .Q (signal_7261) ) ;
    buf_clk cell_5292 ( .C (clk), .D (signal_4733), .Q (signal_7263) ) ;
    buf_clk cell_5294 ( .C (clk), .D (signal_4339), .Q (signal_7265) ) ;
    buf_clk cell_5296 ( .C (clk), .D (signal_4730), .Q (signal_7267) ) ;
    buf_clk cell_5298 ( .C (clk), .D (signal_4307), .Q (signal_7269) ) ;
    buf_clk cell_5300 ( .C (clk), .D (signal_4838), .Q (signal_7271) ) ;
    buf_clk cell_5302 ( .C (clk), .D (signal_4340), .Q (signal_7273) ) ;
    buf_clk cell_5304 ( .C (clk), .D (signal_4727), .Q (signal_7275) ) ;
    buf_clk cell_5306 ( .C (clk), .D (signal_4308), .Q (signal_7277) ) ;
    buf_clk cell_5308 ( .C (clk), .D (signal_4835), .Q (signal_7279) ) ;
    buf_clk cell_5310 ( .C (clk), .D (signal_4341), .Q (signal_7281) ) ;
    buf_clk cell_5312 ( .C (clk), .D (signal_4724), .Q (signal_7283) ) ;
    buf_clk cell_5314 ( .C (clk), .D (signal_4309), .Q (signal_7285) ) ;
    buf_clk cell_5316 ( .C (clk), .D (signal_4829), .Q (signal_7287) ) ;
    buf_clk cell_5318 ( .C (clk), .D (signal_4342), .Q (signal_7289) ) ;
    buf_clk cell_5320 ( .C (clk), .D (signal_4721), .Q (signal_7291) ) ;
    buf_clk cell_5322 ( .C (clk), .D (signal_4310), .Q (signal_7293) ) ;
    buf_clk cell_5324 ( .C (clk), .D (signal_4826), .Q (signal_7295) ) ;
    buf_clk cell_5326 ( .C (clk), .D (signal_4343), .Q (signal_7297) ) ;
    buf_clk cell_5328 ( .C (clk), .D (signal_4718), .Q (signal_7299) ) ;
    buf_clk cell_5330 ( .C (clk), .D (signal_4311), .Q (signal_7301) ) ;
    buf_clk cell_5332 ( .C (clk), .D (signal_4823), .Q (signal_7303) ) ;
    buf_clk cell_5334 ( .C (clk), .D (signal_4279), .Q (signal_7305) ) ;
    buf_clk cell_5336 ( .C (clk), .D (signal_4928), .Q (signal_7307) ) ;
    buf_clk cell_5338 ( .C (clk), .D (signal_4347), .Q (signal_7309) ) ;
    buf_clk cell_5340 ( .C (clk), .D (signal_4706), .Q (signal_7311) ) ;
    buf_clk cell_5342 ( .C (clk), .D (signal_4315), .Q (signal_7313) ) ;
    buf_clk cell_5344 ( .C (clk), .D (signal_4811), .Q (signal_7315) ) ;
    buf_clk cell_5346 ( .C (clk), .D (signal_4283), .Q (signal_7317) ) ;
    buf_clk cell_5348 ( .C (clk), .D (signal_4916), .Q (signal_7319) ) ;
    buf_clk cell_5350 ( .C (clk), .D (signal_4348), .Q (signal_7321) ) ;
    buf_clk cell_5352 ( .C (clk), .D (signal_4703), .Q (signal_7323) ) ;
    buf_clk cell_5354 ( .C (clk), .D (signal_4316), .Q (signal_7325) ) ;
    buf_clk cell_5356 ( .C (clk), .D (signal_4808), .Q (signal_7327) ) ;
    buf_clk cell_5358 ( .C (clk), .D (signal_4284), .Q (signal_7329) ) ;
    buf_clk cell_5360 ( .C (clk), .D (signal_4913), .Q (signal_7331) ) ;
    buf_clk cell_5362 ( .C (clk), .D (signal_4376), .Q (signal_7333) ) ;
    buf_clk cell_5364 ( .C (clk), .D (signal_4700), .Q (signal_7335) ) ;
    buf_clk cell_5366 ( .C (clk), .D (signal_4344), .Q (signal_7337) ) ;
    buf_clk cell_5368 ( .C (clk), .D (signal_4715), .Q (signal_7339) ) ;
    buf_clk cell_5370 ( .C (clk), .D (signal_4312), .Q (signal_7341) ) ;
    buf_clk cell_5372 ( .C (clk), .D (signal_4820), .Q (signal_7343) ) ;
    buf_clk cell_5374 ( .C (clk), .D (signal_4280), .Q (signal_7345) ) ;
    buf_clk cell_5376 ( .C (clk), .D (signal_4925), .Q (signal_7347) ) ;
    buf_clk cell_5378 ( .C (clk), .D (signal_4349), .Q (signal_7349) ) ;
    buf_clk cell_5380 ( .C (clk), .D (signal_4697), .Q (signal_7351) ) ;
    buf_clk cell_5382 ( .C (clk), .D (signal_4317), .Q (signal_7353) ) ;
    buf_clk cell_5384 ( .C (clk), .D (signal_4805), .Q (signal_7355) ) ;
    buf_clk cell_5386 ( .C (clk), .D (signal_4285), .Q (signal_7357) ) ;
    buf_clk cell_5388 ( .C (clk), .D (signal_4910), .Q (signal_7359) ) ;
    buf_clk cell_5390 ( .C (clk), .D (signal_4350), .Q (signal_7361) ) ;
    buf_clk cell_5392 ( .C (clk), .D (signal_4694), .Q (signal_7363) ) ;
    buf_clk cell_5394 ( .C (clk), .D (signal_4318), .Q (signal_7365) ) ;
    buf_clk cell_5396 ( .C (clk), .D (signal_4802), .Q (signal_7367) ) ;
    buf_clk cell_5398 ( .C (clk), .D (signal_4286), .Q (signal_7369) ) ;
    buf_clk cell_5400 ( .C (clk), .D (signal_4907), .Q (signal_7371) ) ;
    buf_clk cell_5402 ( .C (clk), .D (signal_4351), .Q (signal_7373) ) ;
    buf_clk cell_5404 ( .C (clk), .D (signal_4691), .Q (signal_7375) ) ;
    buf_clk cell_5406 ( .C (clk), .D (signal_4319), .Q (signal_7377) ) ;
    buf_clk cell_5408 ( .C (clk), .D (signal_4796), .Q (signal_7379) ) ;
    buf_clk cell_5410 ( .C (clk), .D (signal_4287), .Q (signal_7381) ) ;
    buf_clk cell_5412 ( .C (clk), .D (signal_4904), .Q (signal_7383) ) ;
    buf_clk cell_5414 ( .C (clk), .D (signal_4352), .Q (signal_7385) ) ;
    buf_clk cell_5416 ( .C (clk), .D (signal_4688), .Q (signal_7387) ) ;
    buf_clk cell_5418 ( .C (clk), .D (signal_4320), .Q (signal_7389) ) ;
    buf_clk cell_5420 ( .C (clk), .D (signal_4793), .Q (signal_7391) ) ;
    buf_clk cell_5422 ( .C (clk), .D (signal_4288), .Q (signal_7393) ) ;
    buf_clk cell_5424 ( .C (clk), .D (signal_4901), .Q (signal_7395) ) ;
    buf_clk cell_5426 ( .C (clk), .D (signal_4353), .Q (signal_7397) ) ;
    buf_clk cell_5428 ( .C (clk), .D (signal_4685), .Q (signal_7399) ) ;
    buf_clk cell_5430 ( .C (clk), .D (signal_4321), .Q (signal_7401) ) ;
    buf_clk cell_5432 ( .C (clk), .D (signal_4790), .Q (signal_7403) ) ;
    buf_clk cell_5434 ( .C (clk), .D (signal_4289), .Q (signal_7405) ) ;
    buf_clk cell_5436 ( .C (clk), .D (signal_4895), .Q (signal_7407) ) ;
    buf_clk cell_5438 ( .C (clk), .D (signal_4354), .Q (signal_7409) ) ;
    buf_clk cell_5440 ( .C (clk), .D (signal_4682), .Q (signal_7411) ) ;
    buf_clk cell_5442 ( .C (clk), .D (signal_4322), .Q (signal_7413) ) ;
    buf_clk cell_5444 ( .C (clk), .D (signal_4787), .Q (signal_7415) ) ;
    buf_clk cell_5446 ( .C (clk), .D (signal_4290), .Q (signal_7417) ) ;
    buf_clk cell_5448 ( .C (clk), .D (signal_4892), .Q (signal_7419) ) ;
    buf_clk cell_5450 ( .C (clk), .D (signal_4355), .Q (signal_7421) ) ;
    buf_clk cell_5452 ( .C (clk), .D (signal_4679), .Q (signal_7423) ) ;
    buf_clk cell_5454 ( .C (clk), .D (signal_4323), .Q (signal_7425) ) ;
    buf_clk cell_5456 ( .C (clk), .D (signal_4784), .Q (signal_7427) ) ;
    buf_clk cell_5458 ( .C (clk), .D (signal_4291), .Q (signal_7429) ) ;
    buf_clk cell_5460 ( .C (clk), .D (signal_4889), .Q (signal_7431) ) ;
    buf_clk cell_5462 ( .C (clk), .D (signal_4356), .Q (signal_7433) ) ;
    buf_clk cell_5464 ( .C (clk), .D (signal_4676), .Q (signal_7435) ) ;
    buf_clk cell_5466 ( .C (clk), .D (signal_4324), .Q (signal_7437) ) ;
    buf_clk cell_5468 ( .C (clk), .D (signal_4781), .Q (signal_7439) ) ;
    buf_clk cell_5470 ( .C (clk), .D (signal_4292), .Q (signal_7441) ) ;
    buf_clk cell_5472 ( .C (clk), .D (signal_4886), .Q (signal_7443) ) ;
    buf_clk cell_5474 ( .C (clk), .D (signal_4357), .Q (signal_7445) ) ;
    buf_clk cell_5476 ( .C (clk), .D (signal_4673), .Q (signal_7447) ) ;
    buf_clk cell_5478 ( .C (clk), .D (signal_4325), .Q (signal_7449) ) ;
    buf_clk cell_5480 ( .C (clk), .D (signal_4778), .Q (signal_7451) ) ;
    buf_clk cell_5482 ( .C (clk), .D (signal_4293), .Q (signal_7453) ) ;
    buf_clk cell_5484 ( .C (clk), .D (signal_4883), .Q (signal_7455) ) ;
    buf_clk cell_5486 ( .C (clk), .D (signal_4358), .Q (signal_7457) ) ;
    buf_clk cell_5488 ( .C (clk), .D (signal_4670), .Q (signal_7459) ) ;
    buf_clk cell_5490 ( .C (clk), .D (signal_4326), .Q (signal_7461) ) ;
    buf_clk cell_5492 ( .C (clk), .D (signal_4775), .Q (signal_7463) ) ;
    buf_clk cell_5494 ( .C (clk), .D (signal_4294), .Q (signal_7465) ) ;
    buf_clk cell_5496 ( .C (clk), .D (signal_4880), .Q (signal_7467) ) ;
    buf_clk cell_5498 ( .C (clk), .D (signal_4377), .Q (signal_7469) ) ;
    buf_clk cell_5500 ( .C (clk), .D (signal_4667), .Q (signal_7471) ) ;
    buf_clk cell_5502 ( .C (clk), .D (signal_4345), .Q (signal_7473) ) ;
    buf_clk cell_5504 ( .C (clk), .D (signal_4712), .Q (signal_7475) ) ;
    buf_clk cell_5506 ( .C (clk), .D (signal_4313), .Q (signal_7477) ) ;
    buf_clk cell_5508 ( .C (clk), .D (signal_4817), .Q (signal_7479) ) ;
    buf_clk cell_5510 ( .C (clk), .D (signal_4281), .Q (signal_7481) ) ;
    buf_clk cell_5512 ( .C (clk), .D (signal_4922), .Q (signal_7483) ) ;
    buf_clk cell_5514 ( .C (clk), .D (signal_4359), .Q (signal_7485) ) ;
    buf_clk cell_5516 ( .C (clk), .D (signal_4664), .Q (signal_7487) ) ;
    buf_clk cell_5518 ( .C (clk), .D (signal_4327), .Q (signal_7489) ) ;
    buf_clk cell_5520 ( .C (clk), .D (signal_4772), .Q (signal_7491) ) ;
    buf_clk cell_5522 ( .C (clk), .D (signal_4295), .Q (signal_7493) ) ;
    buf_clk cell_5524 ( .C (clk), .D (signal_4877), .Q (signal_7495) ) ;
    buf_clk cell_5526 ( .C (clk), .D (signal_4360), .Q (signal_7497) ) ;
    buf_clk cell_5528 ( .C (clk), .D (signal_4661), .Q (signal_7499) ) ;
    buf_clk cell_5530 ( .C (clk), .D (signal_4328), .Q (signal_7501) ) ;
    buf_clk cell_5532 ( .C (clk), .D (signal_4769), .Q (signal_7503) ) ;
    buf_clk cell_5534 ( .C (clk), .D (signal_4296), .Q (signal_7505) ) ;
    buf_clk cell_5536 ( .C (clk), .D (signal_4874), .Q (signal_7507) ) ;
    buf_clk cell_5538 ( .C (clk), .D (signal_4361), .Q (signal_7509) ) ;
    buf_clk cell_5540 ( .C (clk), .D (signal_4658), .Q (signal_7511) ) ;
    buf_clk cell_5542 ( .C (clk), .D (signal_4329), .Q (signal_7513) ) ;
    buf_clk cell_5544 ( .C (clk), .D (signal_4763), .Q (signal_7515) ) ;
    buf_clk cell_5546 ( .C (clk), .D (signal_4297), .Q (signal_7517) ) ;
    buf_clk cell_5548 ( .C (clk), .D (signal_4871), .Q (signal_7519) ) ;
    buf_clk cell_5550 ( .C (clk), .D (signal_4362), .Q (signal_7521) ) ;
    buf_clk cell_5552 ( .C (clk), .D (signal_4655), .Q (signal_7523) ) ;
    buf_clk cell_5554 ( .C (clk), .D (signal_4330), .Q (signal_7525) ) ;
    buf_clk cell_5556 ( .C (clk), .D (signal_4760), .Q (signal_7527) ) ;
    buf_clk cell_5558 ( .C (clk), .D (signal_4298), .Q (signal_7529) ) ;
    buf_clk cell_5560 ( .C (clk), .D (signal_4868), .Q (signal_7531) ) ;
    buf_clk cell_5562 ( .C (clk), .D (signal_4363), .Q (signal_7533) ) ;
    buf_clk cell_5564 ( .C (clk), .D (signal_4652), .Q (signal_7535) ) ;
    buf_clk cell_5566 ( .C (clk), .D (signal_4331), .Q (signal_7537) ) ;
    buf_clk cell_5568 ( .C (clk), .D (signal_4757), .Q (signal_7539) ) ;
    buf_clk cell_5570 ( .C (clk), .D (signal_4299), .Q (signal_7541) ) ;
    buf_clk cell_5572 ( .C (clk), .D (signal_4862), .Q (signal_7543) ) ;
    buf_clk cell_5574 ( .C (clk), .D (signal_4364), .Q (signal_7545) ) ;
    buf_clk cell_5576 ( .C (clk), .D (signal_4649), .Q (signal_7547) ) ;
    buf_clk cell_5578 ( .C (clk), .D (signal_4332), .Q (signal_7549) ) ;
    buf_clk cell_5580 ( .C (clk), .D (signal_4754), .Q (signal_7551) ) ;
    buf_clk cell_5582 ( .C (clk), .D (signal_4300), .Q (signal_7553) ) ;
    buf_clk cell_5584 ( .C (clk), .D (signal_4859), .Q (signal_7555) ) ;
    buf_clk cell_5586 ( .C (clk), .D (signal_4365), .Q (signal_7557) ) ;
    buf_clk cell_5588 ( .C (clk), .D (signal_4646), .Q (signal_7559) ) ;
    buf_clk cell_5590 ( .C (clk), .D (signal_4333), .Q (signal_7561) ) ;
    buf_clk cell_5592 ( .C (clk), .D (signal_4751), .Q (signal_7563) ) ;
    buf_clk cell_5594 ( .C (clk), .D (signal_4301), .Q (signal_7565) ) ;
    buf_clk cell_5596 ( .C (clk), .D (signal_4856), .Q (signal_7567) ) ;
    buf_clk cell_5598 ( .C (clk), .D (signal_4366), .Q (signal_7569) ) ;
    buf_clk cell_5600 ( .C (clk), .D (signal_4643), .Q (signal_7571) ) ;
    buf_clk cell_5602 ( .C (clk), .D (signal_4334), .Q (signal_7573) ) ;
    buf_clk cell_5604 ( .C (clk), .D (signal_4748), .Q (signal_7575) ) ;
    buf_clk cell_5606 ( .C (clk), .D (signal_4302), .Q (signal_7577) ) ;
    buf_clk cell_5608 ( .C (clk), .D (signal_4853), .Q (signal_7579) ) ;
    buf_clk cell_5610 ( .C (clk), .D (signal_4251), .Q (signal_7581) ) ;
    buf_clk cell_5612 ( .C (clk), .D (signal_4640), .Q (signal_7583) ) ;
    buf_clk cell_5614 ( .C (clk), .D (signal_4252), .Q (signal_7585) ) ;
    buf_clk cell_5616 ( .C (clk), .D (signal_4637), .Q (signal_7587) ) ;
    buf_clk cell_5618 ( .C (clk), .D (signal_4253), .Q (signal_7589) ) ;
    buf_clk cell_5620 ( .C (clk), .D (signal_4634), .Q (signal_7591) ) ;
    buf_clk cell_5622 ( .C (clk), .D (signal_4254), .Q (signal_7593) ) ;
    buf_clk cell_5624 ( .C (clk), .D (signal_4631), .Q (signal_7595) ) ;
    buf_clk cell_5626 ( .C (clk), .D (signal_4255), .Q (signal_7597) ) ;
    buf_clk cell_5628 ( .C (clk), .D (signal_4628), .Q (signal_7599) ) ;
    buf_clk cell_5630 ( .C (clk), .D (signal_4256), .Q (signal_7601) ) ;
    buf_clk cell_5632 ( .C (clk), .D (signal_4625), .Q (signal_7603) ) ;
    buf_clk cell_5634 ( .C (clk), .D (signal_4257), .Q (signal_7605) ) ;
    buf_clk cell_5636 ( .C (clk), .D (signal_4622), .Q (signal_7607) ) ;
    buf_clk cell_5638 ( .C (clk), .D (signal_4258), .Q (signal_7609) ) ;
    buf_clk cell_5640 ( .C (clk), .D (signal_4619), .Q (signal_7611) ) ;
    buf_clk cell_5642 ( .C (clk), .D (signal_4367), .Q (signal_7613) ) ;
    buf_clk cell_5644 ( .C (clk), .D (signal_4616), .Q (signal_7615) ) ;
    buf_clk cell_5646 ( .C (clk), .D (signal_4335), .Q (signal_7617) ) ;
    buf_clk cell_5648 ( .C (clk), .D (signal_4745), .Q (signal_7619) ) ;
    buf_clk cell_5650 ( .C (clk), .D (signal_4303), .Q (signal_7621) ) ;
    buf_clk cell_5652 ( .C (clk), .D (signal_4850), .Q (signal_7623) ) ;
    buf_clk cell_5654 ( .C (clk), .D (signal_4259), .Q (signal_7625) ) ;
    buf_clk cell_5656 ( .C (clk), .D (signal_4613), .Q (signal_7627) ) ;
    buf_clk cell_5658 ( .C (clk), .D (signal_4260), .Q (signal_7629) ) ;
    buf_clk cell_5660 ( .C (clk), .D (signal_4610), .Q (signal_7631) ) ;
    buf_clk cell_5662 ( .C (clk), .D (signal_4261), .Q (signal_7633) ) ;
    buf_clk cell_5664 ( .C (clk), .D (signal_4607), .Q (signal_7635) ) ;
    buf_clk cell_5666 ( .C (clk), .D (signal_4262), .Q (signal_7637) ) ;
    buf_clk cell_5668 ( .C (clk), .D (signal_4604), .Q (signal_7639) ) ;
    buf_clk cell_5670 ( .C (clk), .D (signal_4263), .Q (signal_7641) ) ;
    buf_clk cell_5672 ( .C (clk), .D (signal_4601), .Q (signal_7643) ) ;
    buf_clk cell_5674 ( .C (clk), .D (signal_4264), .Q (signal_7645) ) ;
    buf_clk cell_5676 ( .C (clk), .D (signal_4598), .Q (signal_7647) ) ;
    buf_clk cell_5678 ( .C (clk), .D (signal_4265), .Q (signal_7649) ) ;
    buf_clk cell_5680 ( .C (clk), .D (signal_4595), .Q (signal_7651) ) ;
    buf_clk cell_5682 ( .C (clk), .D (signal_4266), .Q (signal_7653) ) ;
    buf_clk cell_5684 ( .C (clk), .D (signal_4592), .Q (signal_7655) ) ;
    buf_clk cell_5686 ( .C (clk), .D (signal_4267), .Q (signal_7657) ) ;
    buf_clk cell_5688 ( .C (clk), .D (signal_4589), .Q (signal_7659) ) ;
    buf_clk cell_5690 ( .C (clk), .D (signal_4268), .Q (signal_7661) ) ;
    buf_clk cell_5692 ( .C (clk), .D (signal_4586), .Q (signal_7663) ) ;
    buf_clk cell_5694 ( .C (clk), .D (signal_4368), .Q (signal_7665) ) ;
    buf_clk cell_5696 ( .C (clk), .D (signal_4583), .Q (signal_7667) ) ;
    buf_clk cell_5698 ( .C (clk), .D (signal_4336), .Q (signal_7669) ) ;
    buf_clk cell_5700 ( .C (clk), .D (signal_4742), .Q (signal_7671) ) ;
    buf_clk cell_5702 ( .C (clk), .D (signal_4304), .Q (signal_7673) ) ;
    buf_clk cell_5704 ( .C (clk), .D (signal_4847), .Q (signal_7675) ) ;
    buf_clk cell_5706 ( .C (clk), .D (signal_4269), .Q (signal_7677) ) ;
    buf_clk cell_5708 ( .C (clk), .D (signal_4580), .Q (signal_7679) ) ;
    buf_clk cell_5710 ( .C (clk), .D (signal_4270), .Q (signal_7681) ) ;
    buf_clk cell_5712 ( .C (clk), .D (signal_4577), .Q (signal_7683) ) ;
    buf_clk cell_5714 ( .C (clk), .D (signal_4271), .Q (signal_7685) ) ;
    buf_clk cell_5716 ( .C (clk), .D (signal_4574), .Q (signal_7687) ) ;
    buf_clk cell_5718 ( .C (clk), .D (signal_4272), .Q (signal_7689) ) ;
    buf_clk cell_5720 ( .C (clk), .D (signal_4571), .Q (signal_7691) ) ;
    buf_clk cell_5722 ( .C (clk), .D (signal_4273), .Q (signal_7693) ) ;
    buf_clk cell_5724 ( .C (clk), .D (signal_4568), .Q (signal_7695) ) ;
    buf_clk cell_5726 ( .C (clk), .D (signal_4274), .Q (signal_7697) ) ;
    buf_clk cell_5728 ( .C (clk), .D (signal_4565), .Q (signal_7699) ) ;
    buf_clk cell_5730 ( .C (clk), .D (signal_4275), .Q (signal_7701) ) ;
    buf_clk cell_5732 ( .C (clk), .D (signal_4562), .Q (signal_7703) ) ;
    buf_clk cell_5734 ( .C (clk), .D (signal_4276), .Q (signal_7705) ) ;
    buf_clk cell_5736 ( .C (clk), .D (signal_4559), .Q (signal_7707) ) ;
    buf_clk cell_5738 ( .C (clk), .D (signal_4277), .Q (signal_7709) ) ;
    buf_clk cell_5740 ( .C (clk), .D (signal_4556), .Q (signal_7711) ) ;
    buf_clk cell_5742 ( .C (clk), .D (signal_4278), .Q (signal_7713) ) ;
    buf_clk cell_5744 ( .C (clk), .D (signal_4553), .Q (signal_7715) ) ;
    buf_clk cell_5746 ( .C (clk), .D (signal_4378), .Q (signal_7717) ) ;
    buf_clk cell_5748 ( .C (clk), .D (signal_4550), .Q (signal_7719) ) ;
    buf_clk cell_5750 ( .C (clk), .D (signal_4346), .Q (signal_7721) ) ;
    buf_clk cell_5752 ( .C (clk), .D (signal_4709), .Q (signal_7723) ) ;
    buf_clk cell_5754 ( .C (clk), .D (signal_4314), .Q (signal_7725) ) ;
    buf_clk cell_5756 ( .C (clk), .D (signal_4814), .Q (signal_7727) ) ;
    buf_clk cell_5758 ( .C (clk), .D (signal_4282), .Q (signal_7729) ) ;
    buf_clk cell_5760 ( .C (clk), .D (signal_4919), .Q (signal_7731) ) ;
    buf_clk cell_5762 ( .C (clk), .D (signal_393), .Q (signal_7733) ) ;
    buf_clk cell_5764 ( .C (clk), .D (signal_394), .Q (signal_7735) ) ;
    buf_clk cell_5766 ( .C (clk), .D (signal_4379), .Q (signal_7737) ) ;
    buf_clk cell_5768 ( .C (clk), .D (signal_4380), .Q (signal_7739) ) ;
    buf_clk cell_5770 ( .C (clk), .D (signal_4381), .Q (signal_7741) ) ;
    buf_clk cell_5772 ( .C (clk), .D (signal_4382), .Q (signal_7743) ) ;
    buf_clk cell_5774 ( .C (clk), .D (signal_4383), .Q (signal_7745) ) ;
    buf_clk cell_5776 ( .C (clk), .D (signal_4384), .Q (signal_7747) ) ;
    buf_clk cell_5778 ( .C (clk), .D (signal_3612), .Q (signal_7749) ) ;
    buf_clk cell_5780 ( .C (clk), .D (signal_3610), .Q (signal_7751) ) ;
    buf_clk cell_5782 ( .C (clk), .D (signal_3607), .Q (signal_7753) ) ;
    buf_clk cell_5784 ( .C (clk), .D (signal_3608), .Q (signal_7755) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_28 ( .s (signal_6182), .b ({signal_5012, signal_3994}), .a ({signal_5364, signal_4122}), .c ({signal_5394, signal_3742}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_29 ( .s (signal_6182), .b ({signal_5150, signal_4415}), .a ({signal_5039, signal_4022}), .c ({signal_5237, signal_3642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_30 ( .s (signal_6182), .b ({signal_5149, signal_4414}), .a ({signal_5038, signal_4021}), .c ({signal_5238, signal_3641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_31 ( .s (signal_6182), .b ({signal_5148, signal_4413}), .a ({signal_5037, signal_4020}), .c ({signal_5239, signal_3640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_32 ( .s (signal_6182), .b ({signal_5152, signal_4420}), .a ({signal_5036, signal_4019}), .c ({signal_5240, signal_3639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_33 ( .s (signal_6182), .b ({signal_4973, signal_3890}), .a ({signal_5035, signal_4018}), .c ({signal_5241, signal_3638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_34 ( .s (signal_6182), .b ({signal_5146, signal_4410}), .a ({signal_5357, signal_4017}), .c ({signal_5395, signal_3637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_35 ( .s (signal_6182), .b ({signal_4972, signal_3888}), .a ({signal_5034, signal_4016}), .c ({signal_5242, signal_3636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_36 ( .s (signal_6184), .b ({signal_4971, signal_3887}), .a ({signal_5033, signal_4015}), .c ({signal_5243, signal_3635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_37 ( .s (signal_6186), .b ({signal_5145, signal_4407}), .a ({signal_5032, signal_4014}), .c ({signal_5244, signal_3634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_38 ( .s (signal_6188), .b ({signal_5144, signal_4406}), .a ({signal_5031, signal_4013}), .c ({signal_5245, signal_3633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_39 ( .s (signal_6190), .b ({signal_5008, signal_3984}), .a ({signal_5124, signal_4112}), .c ({signal_5246, signal_3732}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_40 ( .s (signal_6192), .b ({signal_5143, signal_4405}), .a ({signal_5030, signal_4012}), .c ({signal_5247, signal_3632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_41 ( .s (signal_6194), .b ({signal_5147, signal_4412}), .a ({signal_5029, signal_4011}), .c ({signal_5248, signal_3631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_42 ( .s (signal_6192), .b ({signal_4970, signal_3882}), .a ({signal_5028, signal_4010}), .c ({signal_5249, signal_3630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_43 ( .s (signal_6190), .b ({signal_5141, signal_4402}), .a ({signal_5027, signal_4009}), .c ({signal_5250, signal_3629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_44 ( .s (signal_6190), .b ({signal_4969, signal_3880}), .a ({signal_5026, signal_4008}), .c ({signal_5251, signal_3628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_45 ( .s (signal_6184), .b ({signal_4968, signal_3879}), .a ({signal_5025, signal_4007}), .c ({signal_5252, signal_3627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_46 ( .s (signal_6186), .b ({signal_5140, signal_4399}), .a ({signal_5024, signal_4006}), .c ({signal_5253, signal_3626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_47 ( .s (signal_6188), .b ({signal_5139, signal_4398}), .a ({signal_5023, signal_4005}), .c ({signal_5254, signal_3625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_48 ( .s (signal_6192), .b ({signal_5138, signal_4397}), .a ({signal_5022, signal_4004}), .c ({signal_5255, signal_3624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_49 ( .s (signal_6194), .b ({signal_5142, signal_4404}), .a ({signal_5021, signal_4003}), .c ({signal_5256, signal_3623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_50 ( .s (signal_6194), .b ({signal_5007, signal_3983}), .a ({signal_5123, signal_4111}), .c ({signal_5257, signal_3731}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_51 ( .s (signal_6192), .b ({signal_4967, signal_3874}), .a ({signal_5020, signal_4002}), .c ({signal_5258, signal_3622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_52 ( .s (signal_6190), .b ({signal_5136, signal_4394}), .a ({signal_5019, signal_4001}), .c ({signal_5259, signal_3621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_53 ( .s (signal_6192), .b ({signal_4966, signal_3872}), .a ({signal_5018, signal_4000}), .c ({signal_5260, signal_3620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_54 ( .s (signal_6194), .b ({signal_4965, signal_3871}), .a ({signal_5017, signal_3999}), .c ({signal_5261, signal_3619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_55 ( .s (signal_6186), .b ({signal_5135, signal_4391}), .a ({signal_5016, signal_3998}), .c ({signal_5262, signal_3618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_56 ( .s (signal_6194), .b ({signal_5134, signal_4390}), .a ({signal_5015, signal_3997}), .c ({signal_5263, signal_3617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_57 ( .s (signal_6186), .b ({signal_5133, signal_4389}), .a ({signal_5014, signal_3996}), .c ({signal_5264, signal_3616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_58 ( .s (signal_6188), .b ({signal_5137, signal_4396}), .a ({signal_5013, signal_3995}), .c ({signal_5265, signal_3615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_59 ( .s (signal_6184), .b ({signal_5205, signal_4503}), .a ({signal_5122, signal_4110}), .c ({signal_5266, signal_3730}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_60 ( .s (signal_6188), .b ({signal_5204, signal_4502}), .a ({signal_5121, signal_4109}), .c ({signal_5267, signal_3729}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_61 ( .s (signal_6186), .b ({signal_5203, signal_4501}), .a ({signal_5120, signal_4108}), .c ({signal_5268, signal_3728}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_62 ( .s (signal_6188), .b ({signal_5207, signal_4508}), .a ({signal_5119, signal_4107}), .c ({signal_5269, signal_3727}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_63 ( .s (signal_6184), .b ({signal_5006, signal_3978}), .a ({signal_5118, signal_4106}), .c ({signal_5270, signal_3726}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_64 ( .s (signal_6190), .b ({signal_5201, signal_4498}), .a ({signal_5117, signal_4105}), .c ({signal_5271, signal_3725}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_65 ( .s (signal_6192), .b ({signal_5005, signal_3976}), .a ({signal_5116, signal_4104}), .c ({signal_5272, signal_3724}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_66 ( .s (signal_6194), .b ({signal_5004, signal_3975}), .a ({signal_5115, signal_4103}), .c ({signal_5273, signal_3723}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_67 ( .s (signal_6190), .b ({signal_5211, signal_4514}), .a ({signal_5132, signal_4121}), .c ({signal_5274, signal_3741}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_68 ( .s (signal_6192), .b ({signal_5200, signal_4495}), .a ({signal_5114, signal_4102}), .c ({signal_5275, signal_3722}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_69 ( .s (signal_6186), .b ({signal_5199, signal_4494}), .a ({signal_5113, signal_4101}), .c ({signal_5276, signal_3721}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_70 ( .s (signal_6188), .b ({signal_5198, signal_4493}), .a ({signal_5112, signal_4100}), .c ({signal_5277, signal_3720}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_71 ( .s (signal_6184), .b ({signal_5202, signal_4500}), .a ({signal_5111, signal_4099}), .c ({signal_5278, signal_3719}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_72 ( .s (signal_6194), .b ({signal_5003, signal_3970}), .a ({signal_5110, signal_4098}), .c ({signal_5279, signal_3718}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_73 ( .s (signal_6190), .b ({signal_5196, signal_4490}), .a ({signal_5109, signal_4097}), .c ({signal_5280, signal_3717}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_74 ( .s (signal_6186), .b ({signal_5002, signal_3968}), .a ({signal_5108, signal_4096}), .c ({signal_5281, signal_3716}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_75 ( .s (signal_6188), .b ({signal_5001, signal_3967}), .a ({signal_5107, signal_4095}), .c ({signal_5282, signal_3715}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_76 ( .s (signal_6184), .b ({signal_5195, signal_4487}), .a ({signal_5106, signal_4094}), .c ({signal_5283, signal_3714}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_77 ( .s (signal_6192), .b ({signal_5194, signal_4486}), .a ({signal_5105, signal_4093}), .c ({signal_5284, signal_3713}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_78 ( .s (signal_6184), .b ({signal_5011, signal_3992}), .a ({signal_5131, signal_4120}), .c ({signal_5285, signal_3740}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_79 ( .s (signal_6194), .b ({signal_5193, signal_4485}), .a ({signal_5104, signal_4092}), .c ({signal_5286, signal_3712}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_80 ( .s (signal_6190), .b ({signal_5197, signal_4492}), .a ({signal_5103, signal_4091}), .c ({signal_5287, signal_3711}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_81 ( .s (signal_6186), .b ({signal_5000, signal_3962}), .a ({signal_5362, signal_4090}), .c ({signal_5396, signal_3710}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_82 ( .s (signal_6188), .b ({signal_5191, signal_4482}), .a ({signal_5102, signal_4089}), .c ({signal_5288, signal_3709}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_83 ( .s (signal_6184), .b ({signal_4999, signal_3960}), .a ({signal_5101, signal_4088}), .c ({signal_5289, signal_3708}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_84 ( .s (signal_6194), .b ({signal_4998, signal_3959}), .a ({signal_5100, signal_4087}), .c ({signal_5290, signal_3707}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_85 ( .s (signal_6194), .b ({signal_5190, signal_4479}), .a ({signal_5099, signal_4086}), .c ({signal_5291, signal_3706}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_86 ( .s (signal_6194), .b ({signal_5189, signal_4478}), .a ({signal_5098, signal_4085}), .c ({signal_5292, signal_3705}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_87 ( .s (signal_6194), .b ({signal_5188, signal_4477}), .a ({signal_5097, signal_4084}), .c ({signal_5293, signal_3704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_88 ( .s (signal_6194), .b ({signal_5192, signal_4484}), .a ({signal_5096, signal_4083}), .c ({signal_5294, signal_3703}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_89 ( .s (signal_6194), .b ({signal_5010, signal_3991}), .a ({signal_5130, signal_4119}), .c ({signal_5295, signal_3739}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_90 ( .s (signal_6194), .b ({signal_4997, signal_3954}), .a ({signal_5095, signal_4082}), .c ({signal_5296, signal_3702}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_91 ( .s (signal_6194), .b ({signal_5186, signal_4474}), .a ({signal_5361, signal_4081}), .c ({signal_5397, signal_3701}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_92 ( .s (signal_6194), .b ({signal_4996, signal_3952}), .a ({signal_5094, signal_4080}), .c ({signal_5297, signal_3700}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_93 ( .s (signal_6194), .b ({signal_4995, signal_3951}), .a ({signal_5093, signal_4079}), .c ({signal_5298, signal_3699}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_94 ( .s (signal_6194), .b ({signal_5185, signal_4471}), .a ({signal_5092, signal_4078}), .c ({signal_5299, signal_3698}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_95 ( .s (signal_6194), .b ({signal_5184, signal_4470}), .a ({signal_5091, signal_4077}), .c ({signal_5300, signal_3697}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_96 ( .s (signal_6192), .b ({signal_5183, signal_4469}), .a ({signal_5090, signal_4076}), .c ({signal_5301, signal_3696}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_97 ( .s (signal_6192), .b ({signal_5187, signal_4476}), .a ({signal_5089, signal_4075}), .c ({signal_5302, signal_3695}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_98 ( .s (signal_6192), .b ({signal_4994, signal_3946}), .a ({signal_5088, signal_4074}), .c ({signal_5303, signal_3694}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_99 ( .s (signal_6192), .b ({signal_5181, signal_4466}), .a ({signal_5087, signal_4073}), .c ({signal_5304, signal_3693}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_100 ( .s (signal_6192), .b ({signal_5210, signal_4511}), .a ({signal_5129, signal_4118}), .c ({signal_5305, signal_3738}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_101 ( .s (signal_6192), .b ({signal_4993, signal_3944}), .a ({signal_5086, signal_4072}), .c ({signal_5306, signal_3692}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_102 ( .s (signal_6192), .b ({signal_4992, signal_3943}), .a ({signal_5085, signal_4071}), .c ({signal_5307, signal_3691}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_103 ( .s (signal_6192), .b ({signal_5180, signal_4463}), .a ({signal_5084, signal_4070}), .c ({signal_5308, signal_3690}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_104 ( .s (signal_6192), .b ({signal_5179, signal_4462}), .a ({signal_5083, signal_4069}), .c ({signal_5309, signal_3689}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_105 ( .s (signal_6192), .b ({signal_5178, signal_4461}), .a ({signal_5082, signal_4068}), .c ({signal_5310, signal_3688}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_106 ( .s (signal_6192), .b ({signal_5182, signal_4468}), .a ({signal_5081, signal_4067}), .c ({signal_5311, signal_3687}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_107 ( .s (signal_6192), .b ({signal_4991, signal_3938}), .a ({signal_5080, signal_4066}), .c ({signal_5312, signal_3686}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_108 ( .s (signal_6190), .b ({signal_5176, signal_4458}), .a ({signal_5079, signal_4065}), .c ({signal_5313, signal_3685}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_109 ( .s (signal_6190), .b ({signal_4990, signal_3936}), .a ({signal_5078, signal_4064}), .c ({signal_5314, signal_3684}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_110 ( .s (signal_6190), .b ({signal_4989, signal_3935}), .a ({signal_5077, signal_4063}), .c ({signal_5315, signal_3683}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_111 ( .s (signal_6190), .b ({signal_5209, signal_4510}), .a ({signal_5128, signal_4117}), .c ({signal_5316, signal_3737}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_112 ( .s (signal_6190), .b ({signal_5175, signal_4455}), .a ({signal_5076, signal_4062}), .c ({signal_5317, signal_3682}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_113 ( .s (signal_6190), .b ({signal_5174, signal_4454}), .a ({signal_5075, signal_4061}), .c ({signal_5318, signal_3681}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_114 ( .s (signal_6190), .b ({signal_5173, signal_4453}), .a ({signal_5074, signal_4060}), .c ({signal_5319, signal_3680}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_115 ( .s (signal_6190), .b ({signal_5177, signal_4460}), .a ({signal_5073, signal_4059}), .c ({signal_5320, signal_3679}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_116 ( .s (signal_6190), .b ({signal_4988, signal_3930}), .a ({signal_5360, signal_4058}), .c ({signal_5398, signal_3678}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_117 ( .s (signal_6190), .b ({signal_5171, signal_4450}), .a ({signal_5072, signal_4057}), .c ({signal_5321, signal_3677}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_118 ( .s (signal_6190), .b ({signal_4987, signal_3928}), .a ({signal_5071, signal_4056}), .c ({signal_5322, signal_3676}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_119 ( .s (signal_6190), .b ({signal_4986, signal_3927}), .a ({signal_5070, signal_4055}), .c ({signal_5323, signal_3675}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_120 ( .s (signal_6188), .b ({signal_5170, signal_4447}), .a ({signal_5069, signal_4054}), .c ({signal_5324, signal_3674}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_121 ( .s (signal_6188), .b ({signal_5169, signal_4446}), .a ({signal_5068, signal_4053}), .c ({signal_5325, signal_3673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_122 ( .s (signal_6188), .b ({signal_5208, signal_4509}), .a ({signal_5127, signal_4116}), .c ({signal_5326, signal_3736}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_123 ( .s (signal_6188), .b ({signal_5168, signal_4445}), .a ({signal_5067, signal_4052}), .c ({signal_5327, signal_3672}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_124 ( .s (signal_6188), .b ({signal_5172, signal_4452}), .a ({signal_5066, signal_4051}), .c ({signal_5328, signal_3671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_125 ( .s (signal_6188), .b ({signal_4985, signal_3922}), .a ({signal_5065, signal_4050}), .c ({signal_5329, signal_3670}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_126 ( .s (signal_6188), .b ({signal_5166, signal_4442}), .a ({signal_5359, signal_4049}), .c ({signal_5399, signal_3669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_127 ( .s (signal_6188), .b ({signal_4984, signal_3920}), .a ({signal_5064, signal_4048}), .c ({signal_5330, signal_3668}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_128 ( .s (signal_6188), .b ({signal_4983, signal_3919}), .a ({signal_5063, signal_4047}), .c ({signal_5331, signal_3667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_129 ( .s (signal_6188), .b ({signal_5165, signal_4439}), .a ({signal_5062, signal_4046}), .c ({signal_5332, signal_3666}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_130 ( .s (signal_6188), .b ({signal_5164, signal_4438}), .a ({signal_5061, signal_4045}), .c ({signal_5333, signal_3665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_131 ( .s (signal_6188), .b ({signal_5163, signal_4437}), .a ({signal_5060, signal_4044}), .c ({signal_5334, signal_3664}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_132 ( .s (signal_6186), .b ({signal_5167, signal_4444}), .a ({signal_5059, signal_4043}), .c ({signal_5335, signal_3663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_133 ( .s (signal_6186), .b ({signal_5212, signal_4516}), .a ({signal_5126, signal_4115}), .c ({signal_5336, signal_3735}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_134 ( .s (signal_6186), .b ({signal_4982, signal_3914}), .a ({signal_5058, signal_4042}), .c ({signal_5337, signal_3662}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_135 ( .s (signal_6186), .b ({signal_5161, signal_4434}), .a ({signal_5057, signal_4041}), .c ({signal_5338, signal_3661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_136 ( .s (signal_6186), .b ({signal_4981, signal_3912}), .a ({signal_5056, signal_4040}), .c ({signal_5339, signal_3660}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_137 ( .s (signal_6186), .b ({signal_4980, signal_3911}), .a ({signal_5055, signal_4039}), .c ({signal_5340, signal_3659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_138 ( .s (signal_6186), .b ({signal_5160, signal_4431}), .a ({signal_5054, signal_4038}), .c ({signal_5341, signal_3658}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_139 ( .s (signal_6186), .b ({signal_5159, signal_4430}), .a ({signal_5053, signal_4037}), .c ({signal_5342, signal_3657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_140 ( .s (signal_6186), .b ({signal_5158, signal_4429}), .a ({signal_5052, signal_4036}), .c ({signal_5343, signal_3656}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_141 ( .s (signal_6186), .b ({signal_5162, signal_4436}), .a ({signal_5051, signal_4035}), .c ({signal_5344, signal_3655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_142 ( .s (signal_6186), .b ({signal_4979, signal_3906}), .a ({signal_5050, signal_4034}), .c ({signal_5345, signal_3654}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_143 ( .s (signal_6186), .b ({signal_5156, signal_4426}), .a ({signal_5049, signal_4033}), .c ({signal_5346, signal_3653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_144 ( .s (signal_6184), .b ({signal_5009, signal_3986}), .a ({signal_5125, signal_4114}), .c ({signal_5347, signal_3734}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_145 ( .s (signal_6184), .b ({signal_4978, signal_3904}), .a ({signal_5048, signal_4032}), .c ({signal_5348, signal_3652}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_146 ( .s (signal_6184), .b ({signal_4977, signal_3903}), .a ({signal_5047, signal_4031}), .c ({signal_5349, signal_3651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_147 ( .s (signal_6184), .b ({signal_5155, signal_4423}), .a ({signal_5046, signal_4030}), .c ({signal_5350, signal_3650}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_148 ( .s (signal_6184), .b ({signal_5154, signal_4422}), .a ({signal_5045, signal_4029}), .c ({signal_5351, signal_3649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_149 ( .s (signal_6184), .b ({signal_5153, signal_4421}), .a ({signal_5044, signal_4028}), .c ({signal_5352, signal_3648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_150 ( .s (signal_6184), .b ({signal_5157, signal_4428}), .a ({signal_5043, signal_4027}), .c ({signal_5353, signal_3647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_151 ( .s (signal_6184), .b ({signal_4976, signal_3898}), .a ({signal_5358, signal_4026}), .c ({signal_5400, signal_3646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_152 ( .s (signal_6184), .b ({signal_5151, signal_4418}), .a ({signal_5042, signal_4025}), .c ({signal_5354, signal_3645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_153 ( .s (signal_6184), .b ({signal_4975, signal_3896}), .a ({signal_5041, signal_4024}), .c ({signal_5355, signal_3644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_154 ( .s (signal_6184), .b ({signal_4974, signal_3895}), .a ({signal_5040, signal_4023}), .c ({signal_5356, signal_3643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_155 ( .s (signal_6184), .b ({signal_5206, signal_4506}), .a ({signal_5363, signal_4113}), .c ({signal_5401, signal_3733}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_291 ( .s (signal_6196), .b ({signal_5394, signal_3742}), .a ({signal_6200, signal_6198}), .c ({signal_5723, signal_421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_294 ( .s (signal_6196), .b ({signal_5274, signal_3741}), .a ({signal_6204, signal_6202}), .c ({signal_5403, signal_423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_297 ( .s (signal_6196), .b ({signal_5285, signal_3740}), .a ({signal_6208, signal_6206}), .c ({signal_5405, signal_425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_300 ( .s (signal_6196), .b ({signal_5295, signal_3739}), .a ({signal_6212, signal_6210}), .c ({signal_5407, signal_427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_303 ( .s (signal_6196), .b ({signal_5305, signal_3738}), .a ({signal_6216, signal_6214}), .c ({signal_5409, signal_429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_306 ( .s (signal_6196), .b ({signal_5316, signal_3737}), .a ({signal_6220, signal_6218}), .c ({signal_5411, signal_431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_309 ( .s (signal_6196), .b ({signal_5326, signal_3736}), .a ({signal_6224, signal_6222}), .c ({signal_5413, signal_433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_312 ( .s (signal_6196), .b ({signal_5336, signal_3735}), .a ({signal_6228, signal_6226}), .c ({signal_5415, signal_435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_315 ( .s (signal_6196), .b ({signal_5347, signal_3734}), .a ({signal_6232, signal_6230}), .c ({signal_5417, signal_437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_318 ( .s (signal_6196), .b ({signal_5401, signal_3733}), .a ({signal_6236, signal_6234}), .c ({signal_5725, signal_439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_321 ( .s (signal_6196), .b ({signal_5246, signal_3732}), .a ({signal_6240, signal_6238}), .c ({signal_5419, signal_441}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_324 ( .s (signal_6196), .b ({signal_5257, signal_3731}), .a ({signal_6244, signal_6242}), .c ({signal_5421, signal_443}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_327 ( .s (signal_6196), .b ({signal_5266, signal_3730}), .a ({signal_6248, signal_6246}), .c ({signal_5423, signal_445}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_330 ( .s (signal_6196), .b ({signal_5267, signal_3729}), .a ({signal_6252, signal_6250}), .c ({signal_5425, signal_447}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_333 ( .s (signal_6196), .b ({signal_5268, signal_3728}), .a ({signal_6256, signal_6254}), .c ({signal_5427, signal_449}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_336 ( .s (signal_6196), .b ({signal_5269, signal_3727}), .a ({signal_6260, signal_6258}), .c ({signal_5429, signal_451}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_339 ( .s (signal_6196), .b ({signal_5270, signal_3726}), .a ({signal_6264, signal_6262}), .c ({signal_5431, signal_453}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_342 ( .s (signal_6196), .b ({signal_5271, signal_3725}), .a ({signal_6268, signal_6266}), .c ({signal_5433, signal_455}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_345 ( .s (signal_6196), .b ({signal_5272, signal_3724}), .a ({signal_6272, signal_6270}), .c ({signal_5435, signal_457}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_348 ( .s (signal_6196), .b ({signal_5273, signal_3723}), .a ({signal_6276, signal_6274}), .c ({signal_5437, signal_459}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_351 ( .s (signal_6196), .b ({signal_5275, signal_3722}), .a ({signal_6280, signal_6278}), .c ({signal_5439, signal_461}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_354 ( .s (signal_6196), .b ({signal_5276, signal_3721}), .a ({signal_6284, signal_6282}), .c ({signal_5441, signal_463}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_357 ( .s (signal_6196), .b ({signal_5277, signal_3720}), .a ({signal_6288, signal_6286}), .c ({signal_5443, signal_465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_360 ( .s (signal_6196), .b ({signal_5278, signal_3719}), .a ({signal_6292, signal_6290}), .c ({signal_5445, signal_467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_363 ( .s (signal_6196), .b ({signal_5279, signal_3718}), .a ({signal_6296, signal_6294}), .c ({signal_5447, signal_469}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_366 ( .s (signal_6196), .b ({signal_5280, signal_3717}), .a ({signal_6300, signal_6298}), .c ({signal_5449, signal_471}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_369 ( .s (signal_6196), .b ({signal_5281, signal_3716}), .a ({signal_6304, signal_6302}), .c ({signal_5451, signal_473}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_372 ( .s (signal_6196), .b ({signal_5282, signal_3715}), .a ({signal_6308, signal_6306}), .c ({signal_5453, signal_475}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_375 ( .s (signal_6196), .b ({signal_5283, signal_3714}), .a ({signal_6312, signal_6310}), .c ({signal_5455, signal_477}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_378 ( .s (signal_6196), .b ({signal_5284, signal_3713}), .a ({signal_6316, signal_6314}), .c ({signal_5457, signal_479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_381 ( .s (signal_6196), .b ({signal_5286, signal_3712}), .a ({signal_6320, signal_6318}), .c ({signal_5459, signal_481}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_384 ( .s (signal_6196), .b ({signal_5287, signal_3711}), .a ({signal_6324, signal_6322}), .c ({signal_5461, signal_483}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_387 ( .s (signal_6196), .b ({signal_5396, signal_3710}), .a ({signal_6328, signal_6326}), .c ({signal_5727, signal_485}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_390 ( .s (signal_6196), .b ({signal_5288, signal_3709}), .a ({signal_6332, signal_6330}), .c ({signal_5463, signal_487}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_393 ( .s (signal_6196), .b ({signal_5289, signal_3708}), .a ({signal_6336, signal_6334}), .c ({signal_5465, signal_489}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_396 ( .s (signal_6196), .b ({signal_5290, signal_3707}), .a ({signal_6340, signal_6338}), .c ({signal_5467, signal_491}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_399 ( .s (signal_6196), .b ({signal_5291, signal_3706}), .a ({signal_6344, signal_6342}), .c ({signal_5469, signal_493}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_402 ( .s (signal_6196), .b ({signal_5292, signal_3705}), .a ({signal_6348, signal_6346}), .c ({signal_5471, signal_495}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_405 ( .s (signal_6196), .b ({signal_5293, signal_3704}), .a ({signal_6352, signal_6350}), .c ({signal_5473, signal_497}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_408 ( .s (signal_6196), .b ({signal_5294, signal_3703}), .a ({signal_6356, signal_6354}), .c ({signal_5475, signal_499}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_411 ( .s (signal_6196), .b ({signal_5296, signal_3702}), .a ({signal_6360, signal_6358}), .c ({signal_5477, signal_501}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_414 ( .s (signal_6196), .b ({signal_5397, signal_3701}), .a ({signal_6364, signal_6362}), .c ({signal_5729, signal_503}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_417 ( .s (signal_6196), .b ({signal_5297, signal_3700}), .a ({signal_6368, signal_6366}), .c ({signal_5479, signal_505}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_420 ( .s (signal_6196), .b ({signal_5298, signal_3699}), .a ({signal_6372, signal_6370}), .c ({signal_5481, signal_507}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_423 ( .s (signal_6196), .b ({signal_5299, signal_3698}), .a ({signal_6376, signal_6374}), .c ({signal_5483, signal_509}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_426 ( .s (signal_6196), .b ({signal_5300, signal_3697}), .a ({signal_6380, signal_6378}), .c ({signal_5485, signal_511}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_429 ( .s (signal_6196), .b ({signal_5301, signal_3696}), .a ({signal_6384, signal_6382}), .c ({signal_5487, signal_513}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_432 ( .s (signal_6196), .b ({signal_5302, signal_3695}), .a ({signal_6388, signal_6386}), .c ({signal_5489, signal_515}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_435 ( .s (signal_6196), .b ({signal_5303, signal_3694}), .a ({signal_6392, signal_6390}), .c ({signal_5491, signal_517}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_438 ( .s (signal_6196), .b ({signal_5304, signal_3693}), .a ({signal_6396, signal_6394}), .c ({signal_5493, signal_519}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_441 ( .s (signal_6196), .b ({signal_5306, signal_3692}), .a ({signal_6400, signal_6398}), .c ({signal_5495, signal_521}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_444 ( .s (signal_6196), .b ({signal_5307, signal_3691}), .a ({signal_6404, signal_6402}), .c ({signal_5497, signal_523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_447 ( .s (signal_6196), .b ({signal_5308, signal_3690}), .a ({signal_6408, signal_6406}), .c ({signal_5499, signal_525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_450 ( .s (signal_6196), .b ({signal_5309, signal_3689}), .a ({signal_6412, signal_6410}), .c ({signal_5501, signal_527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_453 ( .s (signal_6196), .b ({signal_5310, signal_3688}), .a ({signal_6416, signal_6414}), .c ({signal_5503, signal_529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_456 ( .s (signal_6196), .b ({signal_5311, signal_3687}), .a ({signal_6420, signal_6418}), .c ({signal_5505, signal_531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_459 ( .s (signal_6196), .b ({signal_5312, signal_3686}), .a ({signal_6424, signal_6422}), .c ({signal_5507, signal_533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_462 ( .s (signal_6196), .b ({signal_5313, signal_3685}), .a ({signal_6428, signal_6426}), .c ({signal_5509, signal_535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_465 ( .s (signal_6196), .b ({signal_5314, signal_3684}), .a ({signal_6432, signal_6430}), .c ({signal_5511, signal_537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_468 ( .s (signal_6196), .b ({signal_5315, signal_3683}), .a ({signal_6436, signal_6434}), .c ({signal_5513, signal_539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_471 ( .s (signal_6196), .b ({signal_5317, signal_3682}), .a ({signal_6440, signal_6438}), .c ({signal_5515, signal_541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_474 ( .s (signal_6196), .b ({signal_5318, signal_3681}), .a ({signal_6444, signal_6442}), .c ({signal_5517, signal_543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_477 ( .s (signal_6196), .b ({signal_5319, signal_3680}), .a ({signal_6448, signal_6446}), .c ({signal_5519, signal_545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_480 ( .s (signal_6196), .b ({signal_5320, signal_3679}), .a ({signal_6452, signal_6450}), .c ({signal_5521, signal_547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_483 ( .s (signal_6196), .b ({signal_5398, signal_3678}), .a ({signal_6456, signal_6454}), .c ({signal_5731, signal_549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_486 ( .s (signal_6196), .b ({signal_5321, signal_3677}), .a ({signal_6460, signal_6458}), .c ({signal_5523, signal_551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_489 ( .s (signal_6196), .b ({signal_5322, signal_3676}), .a ({signal_6464, signal_6462}), .c ({signal_5525, signal_553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_492 ( .s (signal_6196), .b ({signal_5323, signal_3675}), .a ({signal_6468, signal_6466}), .c ({signal_5527, signal_555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_495 ( .s (signal_6196), .b ({signal_5324, signal_3674}), .a ({signal_6472, signal_6470}), .c ({signal_5529, signal_557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_498 ( .s (signal_6196), .b ({signal_5325, signal_3673}), .a ({signal_6476, signal_6474}), .c ({signal_5531, signal_559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_501 ( .s (signal_6196), .b ({signal_5327, signal_3672}), .a ({signal_6480, signal_6478}), .c ({signal_5533, signal_561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_504 ( .s (signal_6196), .b ({signal_5328, signal_3671}), .a ({signal_6484, signal_6482}), .c ({signal_5535, signal_563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_507 ( .s (signal_6196), .b ({signal_5329, signal_3670}), .a ({signal_6488, signal_6486}), .c ({signal_5537, signal_565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_510 ( .s (signal_6196), .b ({signal_5399, signal_3669}), .a ({signal_6492, signal_6490}), .c ({signal_5733, signal_567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_513 ( .s (signal_6196), .b ({signal_5330, signal_3668}), .a ({signal_6496, signal_6494}), .c ({signal_5539, signal_569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_516 ( .s (signal_6196), .b ({signal_5331, signal_3667}), .a ({signal_6500, signal_6498}), .c ({signal_5541, signal_571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_519 ( .s (signal_6196), .b ({signal_5332, signal_3666}), .a ({signal_6504, signal_6502}), .c ({signal_5543, signal_573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_522 ( .s (signal_6196), .b ({signal_5333, signal_3665}), .a ({signal_6508, signal_6506}), .c ({signal_5545, signal_575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_525 ( .s (signal_6196), .b ({signal_5334, signal_3664}), .a ({signal_6512, signal_6510}), .c ({signal_5547, signal_577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_528 ( .s (signal_6196), .b ({signal_5335, signal_3663}), .a ({signal_6516, signal_6514}), .c ({signal_5549, signal_579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_531 ( .s (signal_6196), .b ({signal_5337, signal_3662}), .a ({signal_6520, signal_6518}), .c ({signal_5551, signal_581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_534 ( .s (signal_6196), .b ({signal_5338, signal_3661}), .a ({signal_6524, signal_6522}), .c ({signal_5553, signal_583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_537 ( .s (signal_6196), .b ({signal_5339, signal_3660}), .a ({signal_6528, signal_6526}), .c ({signal_5555, signal_585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_540 ( .s (signal_6196), .b ({signal_5340, signal_3659}), .a ({signal_6532, signal_6530}), .c ({signal_5557, signal_587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_543 ( .s (signal_6196), .b ({signal_5341, signal_3658}), .a ({signal_6536, signal_6534}), .c ({signal_5559, signal_589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_546 ( .s (signal_6196), .b ({signal_5342, signal_3657}), .a ({signal_6540, signal_6538}), .c ({signal_5561, signal_591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_549 ( .s (signal_6196), .b ({signal_5343, signal_3656}), .a ({signal_6544, signal_6542}), .c ({signal_5563, signal_593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_552 ( .s (signal_6196), .b ({signal_5344, signal_3655}), .a ({signal_6548, signal_6546}), .c ({signal_5565, signal_595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_555 ( .s (signal_6196), .b ({signal_5345, signal_3654}), .a ({signal_6552, signal_6550}), .c ({signal_5567, signal_597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_558 ( .s (signal_6196), .b ({signal_5346, signal_3653}), .a ({signal_6556, signal_6554}), .c ({signal_5569, signal_599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_561 ( .s (signal_6196), .b ({signal_5348, signal_3652}), .a ({signal_6560, signal_6558}), .c ({signal_5571, signal_601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_564 ( .s (signal_6196), .b ({signal_5349, signal_3651}), .a ({signal_6564, signal_6562}), .c ({signal_5573, signal_603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_567 ( .s (signal_6196), .b ({signal_5350, signal_3650}), .a ({signal_6568, signal_6566}), .c ({signal_5575, signal_605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_570 ( .s (signal_6196), .b ({signal_5351, signal_3649}), .a ({signal_6572, signal_6570}), .c ({signal_5577, signal_607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_573 ( .s (signal_6196), .b ({signal_5352, signal_3648}), .a ({signal_6576, signal_6574}), .c ({signal_5579, signal_609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_576 ( .s (signal_6196), .b ({signal_5353, signal_3647}), .a ({signal_6580, signal_6578}), .c ({signal_5581, signal_611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_579 ( .s (signal_6196), .b ({signal_5400, signal_3646}), .a ({signal_6584, signal_6582}), .c ({signal_5735, signal_613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_582 ( .s (signal_6196), .b ({signal_5354, signal_3645}), .a ({signal_6588, signal_6586}), .c ({signal_5583, signal_615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_585 ( .s (signal_6196), .b ({signal_5355, signal_3644}), .a ({signal_6592, signal_6590}), .c ({signal_5585, signal_617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_588 ( .s (signal_6196), .b ({signal_5356, signal_3643}), .a ({signal_6596, signal_6594}), .c ({signal_5587, signal_619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_591 ( .s (signal_6196), .b ({signal_5237, signal_3642}), .a ({signal_6600, signal_6598}), .c ({signal_5589, signal_621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_594 ( .s (signal_6196), .b ({signal_5238, signal_3641}), .a ({signal_6604, signal_6602}), .c ({signal_5591, signal_623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_597 ( .s (signal_6196), .b ({signal_5239, signal_3640}), .a ({signal_6608, signal_6606}), .c ({signal_5593, signal_625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_600 ( .s (signal_6196), .b ({signal_5240, signal_3639}), .a ({signal_6612, signal_6610}), .c ({signal_5595, signal_627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_603 ( .s (signal_6196), .b ({signal_5241, signal_3638}), .a ({signal_6616, signal_6614}), .c ({signal_5597, signal_629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_606 ( .s (signal_6196), .b ({signal_5395, signal_3637}), .a ({signal_6620, signal_6618}), .c ({signal_5737, signal_631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_609 ( .s (signal_6196), .b ({signal_5242, signal_3636}), .a ({signal_6624, signal_6622}), .c ({signal_5599, signal_633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_612 ( .s (signal_6196), .b ({signal_5243, signal_3635}), .a ({signal_6628, signal_6626}), .c ({signal_5601, signal_635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_615 ( .s (signal_6196), .b ({signal_5244, signal_3634}), .a ({signal_6632, signal_6630}), .c ({signal_5603, signal_637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_618 ( .s (signal_6196), .b ({signal_5245, signal_3633}), .a ({signal_6636, signal_6634}), .c ({signal_5605, signal_639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_621 ( .s (signal_6196), .b ({signal_5247, signal_3632}), .a ({signal_6640, signal_6638}), .c ({signal_5607, signal_641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_624 ( .s (signal_6196), .b ({signal_5248, signal_3631}), .a ({signal_6644, signal_6642}), .c ({signal_5609, signal_643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_627 ( .s (signal_6196), .b ({signal_5249, signal_3630}), .a ({signal_6648, signal_6646}), .c ({signal_5611, signal_645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_630 ( .s (signal_6196), .b ({signal_5250, signal_3629}), .a ({signal_6652, signal_6650}), .c ({signal_5613, signal_647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_633 ( .s (signal_6196), .b ({signal_5251, signal_3628}), .a ({signal_6656, signal_6654}), .c ({signal_5615, signal_649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_636 ( .s (signal_6196), .b ({signal_5252, signal_3627}), .a ({signal_6660, signal_6658}), .c ({signal_5617, signal_651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_639 ( .s (signal_6196), .b ({signal_5253, signal_3626}), .a ({signal_6664, signal_6662}), .c ({signal_5619, signal_653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_642 ( .s (signal_6196), .b ({signal_5254, signal_3625}), .a ({signal_6668, signal_6666}), .c ({signal_5621, signal_655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_645 ( .s (signal_6196), .b ({signal_5255, signal_3624}), .a ({signal_6672, signal_6670}), .c ({signal_5623, signal_657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_648 ( .s (signal_6196), .b ({signal_5256, signal_3623}), .a ({signal_6676, signal_6674}), .c ({signal_5625, signal_659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_651 ( .s (signal_6196), .b ({signal_5258, signal_3622}), .a ({signal_6680, signal_6678}), .c ({signal_5627, signal_661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_654 ( .s (signal_6196), .b ({signal_5259, signal_3621}), .a ({signal_6684, signal_6682}), .c ({signal_5629, signal_663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_657 ( .s (signal_6196), .b ({signal_5260, signal_3620}), .a ({signal_6688, signal_6686}), .c ({signal_5631, signal_665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_660 ( .s (signal_6196), .b ({signal_5261, signal_3619}), .a ({signal_6692, signal_6690}), .c ({signal_5633, signal_667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_663 ( .s (signal_6196), .b ({signal_5262, signal_3618}), .a ({signal_6696, signal_6694}), .c ({signal_5635, signal_669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_666 ( .s (signal_6196), .b ({signal_5263, signal_3617}), .a ({signal_6700, signal_6698}), .c ({signal_5637, signal_671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_669 ( .s (signal_6196), .b ({signal_5264, signal_3616}), .a ({signal_6704, signal_6702}), .c ({signal_5639, signal_673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_672 ( .s (signal_6196), .b ({signal_5265, signal_3615}), .a ({signal_6708, signal_6706}), .c ({signal_5641, signal_675}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_2723 ( .a ({signal_4949, signal_2597}), .b ({signal_5141, signal_4402}), .c ({signal_5357, signal_4017}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_2815 ( .a ({signal_4950, signal_2660}), .b ({signal_4973, signal_3890}), .c ({signal_5358, signal_4026}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_2831 ( .a ({signal_4951, signal_2661}), .b ({signal_5161, signal_4434}), .c ({signal_5359, signal_4049}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_2923 ( .a ({signal_4952, signal_2724}), .b ({signal_4985, signal_3922}), .c ({signal_5360, signal_4058}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_2939 ( .a ({signal_4953, signal_2725}), .b ({signal_5181, signal_4466}), .c ({signal_5361, signal_4081}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_3031 ( .a ({signal_4954, signal_2788}), .b ({signal_4997, signal_3954}), .c ({signal_5362, signal_4090}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_3047 ( .a ({signal_4955, signal_2789}), .b ({signal_5201, signal_4498}), .c ({signal_5363, signal_4113}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_3139 ( .a ({signal_4956, signal_2852}), .b ({signal_5009, signal_3986}), .c ({signal_5364, signal_4122}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3155 ( .s (signal_6196), .b ({signal_5923, signal_4250}), .a ({signal_6712, signal_6710}), .c ({signal_5925, signal_2853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3158 ( .s (signal_6196), .b ({signal_5912, signal_4249}), .a ({signal_6716, signal_6714}), .c ({signal_5927, signal_2855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3161 ( .s (signal_6196), .b ({signal_5901, signal_4248}), .a ({signal_6720, signal_6718}), .c ({signal_5929, signal_2857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3164 ( .s (signal_6196), .b ({signal_5898, signal_4247}), .a ({signal_6724, signal_6722}), .c ({signal_5931, signal_2859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3167 ( .s (signal_6196), .b ({signal_5897, signal_4246}), .a ({signal_6728, signal_6726}), .c ({signal_5933, signal_2861}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3170 ( .s (signal_6196), .b ({signal_5896, signal_4245}), .a ({signal_6732, signal_6730}), .c ({signal_5935, signal_2863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3173 ( .s (signal_6196), .b ({signal_5895, signal_4244}), .a ({signal_6736, signal_6734}), .c ({signal_5937, signal_2865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3176 ( .s (signal_6196), .b ({signal_5894, signal_4243}), .a ({signal_6740, signal_6738}), .c ({signal_5939, signal_2867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3179 ( .s (signal_6196), .b ({signal_5893, signal_4242}), .a ({signal_6744, signal_6742}), .c ({signal_5941, signal_2869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3182 ( .s (signal_6196), .b ({signal_5892, signal_4241}), .a ({signal_6748, signal_6746}), .c ({signal_5943, signal_2871}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3185 ( .s (signal_6196), .b ({signal_5922, signal_4240}), .a ({signal_6752, signal_6750}), .c ({signal_5945, signal_2873}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3188 ( .s (signal_6196), .b ({signal_5921, signal_4239}), .a ({signal_6756, signal_6754}), .c ({signal_5947, signal_2875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3191 ( .s (signal_6196), .b ({signal_5920, signal_4238}), .a ({signal_6760, signal_6758}), .c ({signal_5949, signal_2877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3194 ( .s (signal_6196), .b ({signal_5919, signal_4237}), .a ({signal_6764, signal_6762}), .c ({signal_5951, signal_2879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3197 ( .s (signal_6196), .b ({signal_5918, signal_4236}), .a ({signal_6768, signal_6766}), .c ({signal_5953, signal_2881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3200 ( .s (signal_6196), .b ({signal_5917, signal_4235}), .a ({signal_6772, signal_6770}), .c ({signal_5955, signal_2883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3203 ( .s (signal_6196), .b ({signal_5916, signal_4234}), .a ({signal_6776, signal_6774}), .c ({signal_5957, signal_2885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3206 ( .s (signal_6196), .b ({signal_5915, signal_4233}), .a ({signal_6780, signal_6778}), .c ({signal_5959, signal_2887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3209 ( .s (signal_6196), .b ({signal_5914, signal_4232}), .a ({signal_6784, signal_6782}), .c ({signal_5961, signal_2889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3212 ( .s (signal_6196), .b ({signal_5913, signal_4231}), .a ({signal_6788, signal_6786}), .c ({signal_5963, signal_2891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3215 ( .s (signal_6196), .b ({signal_5911, signal_4230}), .a ({signal_6792, signal_6790}), .c ({signal_5965, signal_2893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3218 ( .s (signal_6196), .b ({signal_5910, signal_4229}), .a ({signal_6796, signal_6794}), .c ({signal_5967, signal_2895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3221 ( .s (signal_6196), .b ({signal_5909, signal_4228}), .a ({signal_6800, signal_6798}), .c ({signal_5969, signal_2897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3224 ( .s (signal_6196), .b ({signal_5908, signal_4227}), .a ({signal_6804, signal_6802}), .c ({signal_5971, signal_2899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3227 ( .s (signal_6196), .b ({signal_5995, signal_4226}), .a ({signal_6808, signal_6806}), .c ({signal_5997, signal_2901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3230 ( .s (signal_6196), .b ({signal_5994, signal_4225}), .a ({signal_6812, signal_6810}), .c ({signal_5999, signal_2903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3233 ( .s (signal_6196), .b ({signal_6014, signal_4224}), .a ({signal_6816, signal_6814}), .c ({signal_6016, signal_2905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3236 ( .s (signal_6196), .b ({signal_6013, signal_4223}), .a ({signal_6820, signal_6818}), .c ({signal_6018, signal_2907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3239 ( .s (signal_6196), .b ({signal_5991, signal_4222}), .a ({signal_6824, signal_6822}), .c ({signal_6001, signal_2909}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3242 ( .s (signal_6196), .b ({signal_6012, signal_4221}), .a ({signal_6828, signal_6826}), .c ({signal_6020, signal_2911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3245 ( .s (signal_6196), .b ({signal_5989, signal_4220}), .a ({signal_6832, signal_6830}), .c ({signal_6003, signal_2913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3248 ( .s (signal_6196), .b ({signal_5988, signal_4219}), .a ({signal_6836, signal_6834}), .c ({signal_6005, signal_2915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3251 ( .s (signal_6196), .b ({signal_5827, signal_4218}), .a ({signal_6840, signal_6838}), .c ({signal_5829, signal_2917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3254 ( .s (signal_6196), .b ({signal_5813, signal_4217}), .a ({signal_6844, signal_6842}), .c ({signal_5831, signal_2919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3257 ( .s (signal_6196), .b ({signal_5805, signal_4216}), .a ({signal_6848, signal_6846}), .c ({signal_5833, signal_2921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3260 ( .s (signal_6196), .b ({signal_5802, signal_4215}), .a ({signal_6852, signal_6850}), .c ({signal_5835, signal_2923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3263 ( .s (signal_6196), .b ({signal_5801, signal_4214}), .a ({signal_6856, signal_6854}), .c ({signal_5837, signal_2925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3266 ( .s (signal_6196), .b ({signal_5800, signal_4213}), .a ({signal_6860, signal_6858}), .c ({signal_5839, signal_2927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3269 ( .s (signal_6196), .b ({signal_5799, signal_4212}), .a ({signal_6864, signal_6862}), .c ({signal_5841, signal_2929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3272 ( .s (signal_6196), .b ({signal_5798, signal_4211}), .a ({signal_6868, signal_6866}), .c ({signal_5843, signal_2931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3275 ( .s (signal_6196), .b ({signal_5797, signal_4210}), .a ({signal_6872, signal_6870}), .c ({signal_5845, signal_2933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3278 ( .s (signal_6196), .b ({signal_5796, signal_4209}), .a ({signal_6876, signal_6874}), .c ({signal_5847, signal_2935}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3281 ( .s (signal_6196), .b ({signal_5826, signal_4208}), .a ({signal_6880, signal_6878}), .c ({signal_5849, signal_2937}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3284 ( .s (signal_6196), .b ({signal_5825, signal_4207}), .a ({signal_6884, signal_6882}), .c ({signal_5851, signal_2939}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3287 ( .s (signal_6196), .b ({signal_5821, signal_4206}), .a ({signal_6888, signal_6886}), .c ({signal_5853, signal_2941}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3290 ( .s (signal_6196), .b ({signal_5820, signal_4205}), .a ({signal_6892, signal_6890}), .c ({signal_5855, signal_2943}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3293 ( .s (signal_6196), .b ({signal_5819, signal_4204}), .a ({signal_6896, signal_6894}), .c ({signal_5857, signal_2945}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3296 ( .s (signal_6196), .b ({signal_5818, signal_4203}), .a ({signal_6900, signal_6898}), .c ({signal_5859, signal_2947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3299 ( .s (signal_6196), .b ({signal_5817, signal_4202}), .a ({signal_6904, signal_6902}), .c ({signal_5861, signal_2949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3302 ( .s (signal_6196), .b ({signal_5816, signal_4201}), .a ({signal_6908, signal_6906}), .c ({signal_5863, signal_2951}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3305 ( .s (signal_6196), .b ({signal_5815, signal_4200}), .a ({signal_6912, signal_6910}), .c ({signal_5865, signal_2953}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3308 ( .s (signal_6196), .b ({signal_5814, signal_4199}), .a ({signal_6916, signal_6914}), .c ({signal_5867, signal_2955}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3311 ( .s (signal_6196), .b ({signal_5812, signal_4198}), .a ({signal_6920, signal_6918}), .c ({signal_5869, signal_2957}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3314 ( .s (signal_6196), .b ({signal_5811, signal_4197}), .a ({signal_6924, signal_6922}), .c ({signal_5871, signal_2959}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3317 ( .s (signal_6196), .b ({signal_5810, signal_4196}), .a ({signal_6928, signal_6926}), .c ({signal_5873, signal_2961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3320 ( .s (signal_6196), .b ({signal_5809, signal_4195}), .a ({signal_6932, signal_6930}), .c ({signal_5875, signal_2963}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3323 ( .s (signal_6196), .b ({signal_5907, signal_4194}), .a ({signal_6936, signal_6934}), .c ({signal_5973, signal_2965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3326 ( .s (signal_6196), .b ({signal_5906, signal_4193}), .a ({signal_6940, signal_6938}), .c ({signal_5975, signal_2967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3329 ( .s (signal_6196), .b ({signal_5993, signal_4192}), .a ({signal_6944, signal_6942}), .c ({signal_6007, signal_2969}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3332 ( .s (signal_6196), .b ({signal_5992, signal_4191}), .a ({signal_6948, signal_6946}), .c ({signal_6009, signal_2971}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3335 ( .s (signal_6196), .b ({signal_5903, signal_4190}), .a ({signal_6952, signal_6950}), .c ({signal_5977, signal_2973}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3338 ( .s (signal_6196), .b ({signal_5990, signal_4189}), .a ({signal_6956, signal_6954}), .c ({signal_6011, signal_2975}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3341 ( .s (signal_6196), .b ({signal_5900, signal_4188}), .a ({signal_6960, signal_6958}), .c ({signal_5979, signal_2977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3344 ( .s (signal_6196), .b ({signal_5899, signal_4187}), .a ({signal_6964, signal_6962}), .c ({signal_5981, signal_2979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3347 ( .s (signal_6196), .b ({signal_5718, signal_4186}), .a ({signal_6968, signal_6966}), .c ({signal_5739, signal_2981}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3350 ( .s (signal_6196), .b ({signal_5702, signal_4185}), .a ({signal_6972, signal_6970}), .c ({signal_5741, signal_2983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3353 ( .s (signal_6196), .b ({signal_5697, signal_4184}), .a ({signal_6976, signal_6974}), .c ({signal_5743, signal_2985}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3356 ( .s (signal_6196), .b ({signal_5696, signal_4183}), .a ({signal_6980, signal_6978}), .c ({signal_5745, signal_2987}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3359 ( .s (signal_6196), .b ({signal_5695, signal_4182}), .a ({signal_6984, signal_6982}), .c ({signal_5747, signal_2989}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3362 ( .s (signal_6196), .b ({signal_5694, signal_4181}), .a ({signal_6988, signal_6986}), .c ({signal_5749, signal_2991}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3365 ( .s (signal_6196), .b ({signal_5693, signal_4180}), .a ({signal_6992, signal_6990}), .c ({signal_5751, signal_2993}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3368 ( .s (signal_6196), .b ({signal_5692, signal_4179}), .a ({signal_6996, signal_6994}), .c ({signal_5753, signal_2995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3371 ( .s (signal_6196), .b ({signal_5691, signal_4178}), .a ({signal_7000, signal_6998}), .c ({signal_5755, signal_2997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3374 ( .s (signal_6196), .b ({signal_5690, signal_4177}), .a ({signal_7004, signal_7002}), .c ({signal_5757, signal_2999}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3377 ( .s (signal_6196), .b ({signal_5717, signal_4176}), .a ({signal_7008, signal_7006}), .c ({signal_5759, signal_3001}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3380 ( .s (signal_6196), .b ({signal_5716, signal_4175}), .a ({signal_7012, signal_7010}), .c ({signal_5761, signal_3003}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3383 ( .s (signal_6196), .b ({signal_5710, signal_4174}), .a ({signal_7016, signal_7014}), .c ({signal_5763, signal_3005}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3386 ( .s (signal_6196), .b ({signal_5709, signal_4173}), .a ({signal_7020, signal_7018}), .c ({signal_5765, signal_3007}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3389 ( .s (signal_6196), .b ({signal_5708, signal_4172}), .a ({signal_7024, signal_7022}), .c ({signal_5767, signal_3009}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3392 ( .s (signal_6196), .b ({signal_5707, signal_4171}), .a ({signal_7028, signal_7026}), .c ({signal_5769, signal_3011}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3395 ( .s (signal_6196), .b ({signal_5706, signal_4170}), .a ({signal_7032, signal_7030}), .c ({signal_5771, signal_3013}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3398 ( .s (signal_6196), .b ({signal_5705, signal_4169}), .a ({signal_7036, signal_7034}), .c ({signal_5773, signal_3015}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3401 ( .s (signal_6196), .b ({signal_5704, signal_4168}), .a ({signal_7040, signal_7038}), .c ({signal_5775, signal_3017}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3404 ( .s (signal_6196), .b ({signal_5703, signal_4167}), .a ({signal_7044, signal_7042}), .c ({signal_5777, signal_3019}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3407 ( .s (signal_6196), .b ({signal_5701, signal_4166}), .a ({signal_7048, signal_7046}), .c ({signal_5779, signal_3021}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3410 ( .s (signal_6196), .b ({signal_5700, signal_4165}), .a ({signal_7052, signal_7050}), .c ({signal_5781, signal_3023}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3413 ( .s (signal_6196), .b ({signal_5699, signal_4164}), .a ({signal_7056, signal_7054}), .c ({signal_5783, signal_3025}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3416 ( .s (signal_6196), .b ({signal_5698, signal_4163}), .a ({signal_7060, signal_7058}), .c ({signal_5785, signal_3027}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3419 ( .s (signal_6196), .b ({signal_5808, signal_4162}), .a ({signal_7064, signal_7062}), .c ({signal_5877, signal_3029}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3422 ( .s (signal_6196), .b ({signal_5807, signal_4161}), .a ({signal_7068, signal_7066}), .c ({signal_5879, signal_3031}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3425 ( .s (signal_6196), .b ({signal_5905, signal_4160}), .a ({signal_7072, signal_7070}), .c ({signal_5983, signal_3033}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3428 ( .s (signal_6196), .b ({signal_5904, signal_4159}), .a ({signal_7076, signal_7074}), .c ({signal_5985, signal_3035}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3431 ( .s (signal_6196), .b ({signal_5806, signal_4158}), .a ({signal_7080, signal_7078}), .c ({signal_5881, signal_3037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3434 ( .s (signal_6196), .b ({signal_5902, signal_4157}), .a ({signal_7084, signal_7082}), .c ({signal_5987, signal_3039}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3437 ( .s (signal_6196), .b ({signal_5804, signal_4156}), .a ({signal_7088, signal_7086}), .c ({signal_5883, signal_3041}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3440 ( .s (signal_6196), .b ({signal_5803, signal_4155}), .a ({signal_7092, signal_7090}), .c ({signal_5885, signal_3043}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3443 ( .s (signal_6196), .b ({signal_5388, signal_4154}), .a ({signal_7096, signal_7094}), .c ({signal_5643, signal_3045}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3446 ( .s (signal_6196), .b ({signal_5367, signal_4153}), .a ({signal_7100, signal_7098}), .c ({signal_5645, signal_3047}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3449 ( .s (signal_6196), .b ({signal_5366, signal_4152}), .a ({signal_7104, signal_7102}), .c ({signal_5647, signal_3049}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3452 ( .s (signal_6196), .b ({signal_5365, signal_4151}), .a ({signal_7108, signal_7106}), .c ({signal_5649, signal_3051}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3455 ( .s (signal_6196), .b ({signal_5387, signal_4150}), .a ({signal_7112, signal_7110}), .c ({signal_5651, signal_3053}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3458 ( .s (signal_6196), .b ({signal_5386, signal_4149}), .a ({signal_7116, signal_7114}), .c ({signal_5653, signal_3055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3461 ( .s (signal_6196), .b ({signal_5385, signal_4148}), .a ({signal_7120, signal_7118}), .c ({signal_5655, signal_3057}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3464 ( .s (signal_6196), .b ({signal_5384, signal_4147}), .a ({signal_7124, signal_7122}), .c ({signal_5657, signal_3059}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3467 ( .s (signal_6196), .b ({signal_5383, signal_4146}), .a ({signal_7128, signal_7126}), .c ({signal_5659, signal_3061}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3470 ( .s (signal_6196), .b ({signal_5382, signal_4145}), .a ({signal_7132, signal_7130}), .c ({signal_5661, signal_3063}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3473 ( .s (signal_6196), .b ({signal_5381, signal_4144}), .a ({signal_7136, signal_7134}), .c ({signal_5663, signal_3065}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3476 ( .s (signal_6196), .b ({signal_5380, signal_4143}), .a ({signal_7140, signal_7138}), .c ({signal_5665, signal_3067}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3479 ( .s (signal_6196), .b ({signal_5379, signal_4142}), .a ({signal_7144, signal_7142}), .c ({signal_5667, signal_3069}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3482 ( .s (signal_6196), .b ({signal_5378, signal_4141}), .a ({signal_7148, signal_7146}), .c ({signal_5669, signal_3071}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3485 ( .s (signal_6196), .b ({signal_5377, signal_4140}), .a ({signal_7152, signal_7150}), .c ({signal_5671, signal_3073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3488 ( .s (signal_6196), .b ({signal_5376, signal_4139}), .a ({signal_7156, signal_7154}), .c ({signal_5673, signal_3075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3491 ( .s (signal_6196), .b ({signal_5375, signal_4138}), .a ({signal_7160, signal_7158}), .c ({signal_5675, signal_3077}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3494 ( .s (signal_6196), .b ({signal_5374, signal_4137}), .a ({signal_7164, signal_7162}), .c ({signal_5677, signal_3079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3497 ( .s (signal_6196), .b ({signal_5373, signal_4136}), .a ({signal_7168, signal_7166}), .c ({signal_5679, signal_3081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3500 ( .s (signal_6196), .b ({signal_5372, signal_4135}), .a ({signal_7172, signal_7170}), .c ({signal_5681, signal_3083}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3503 ( .s (signal_6196), .b ({signal_5371, signal_4134}), .a ({signal_7176, signal_7174}), .c ({signal_5683, signal_3085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3506 ( .s (signal_6196), .b ({signal_5370, signal_4133}), .a ({signal_7180, signal_7178}), .c ({signal_5685, signal_3087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3509 ( .s (signal_6196), .b ({signal_5369, signal_4132}), .a ({signal_7184, signal_7182}), .c ({signal_5687, signal_3089}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3512 ( .s (signal_6196), .b ({signal_5368, signal_4131}), .a ({signal_7188, signal_7186}), .c ({signal_5689, signal_3091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3515 ( .s (signal_6196), .b ({signal_5715, signal_4130}), .a ({signal_7192, signal_7190}), .c ({signal_5787, signal_3093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3518 ( .s (signal_6196), .b ({signal_5714, signal_4129}), .a ({signal_7196, signal_7194}), .c ({signal_5789, signal_3095}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3521 ( .s (signal_6196), .b ({signal_5824, signal_4128}), .a ({signal_7200, signal_7198}), .c ({signal_5887, signal_3097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3524 ( .s (signal_6196), .b ({signal_5823, signal_4127}), .a ({signal_7204, signal_7202}), .c ({signal_5889, signal_3099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3527 ( .s (signal_6196), .b ({signal_5713, signal_4126}), .a ({signal_7208, signal_7206}), .c ({signal_5791, signal_3101}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3530 ( .s (signal_6196), .b ({signal_5822, signal_4125}), .a ({signal_7212, signal_7210}), .c ({signal_5891, signal_3103}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3533 ( .s (signal_6196), .b ({signal_5712, signal_4124}), .a ({signal_7216, signal_7214}), .c ({signal_5793, signal_3105}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_3536 ( .s (signal_6196), .b ({signal_5711, signal_4123}), .a ({signal_7220, signal_7218}), .c ({signal_5795, signal_3107}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3539 ( .a ({signal_7224, signal_7222}), .b ({signal_5796, signal_4209}), .c ({signal_5892, signal_4241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3540 ( .a ({signal_7228, signal_7226}), .b ({signal_5797, signal_4210}), .c ({signal_5893, signal_4242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3541 ( .a ({signal_7232, signal_7230}), .b ({signal_5798, signal_4211}), .c ({signal_5894, signal_4243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3542 ( .a ({signal_7236, signal_7234}), .b ({signal_5799, signal_4212}), .c ({signal_5895, signal_4244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3543 ( .a ({signal_7240, signal_7238}), .b ({signal_5800, signal_4213}), .c ({signal_5896, signal_4245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3544 ( .a ({signal_7244, signal_7242}), .b ({signal_5801, signal_4214}), .c ({signal_5897, signal_4246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3545 ( .a ({signal_7248, signal_7246}), .b ({signal_5690, signal_4177}), .c ({signal_5796, signal_4209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3546 ( .a ({signal_7252, signal_7250}), .b ({signal_5382, signal_4145}), .c ({signal_5690, signal_4177}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3547 ( .a ({signal_7256, signal_7254}), .b ({signal_5691, signal_4178}), .c ({signal_5797, signal_4210}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3548 ( .a ({signal_7260, signal_7258}), .b ({signal_5383, signal_4146}), .c ({signal_5691, signal_4178}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3549 ( .a ({signal_7264, signal_7262}), .b ({signal_5802, signal_4215}), .c ({signal_5898, signal_4247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3550 ( .a ({signal_7268, signal_7266}), .b ({signal_5692, signal_4179}), .c ({signal_5798, signal_4211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3551 ( .a ({signal_7272, signal_7270}), .b ({signal_5384, signal_4147}), .c ({signal_5692, signal_4179}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3552 ( .a ({signal_7276, signal_7274}), .b ({signal_5693, signal_4180}), .c ({signal_5799, signal_4212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3553 ( .a ({signal_7280, signal_7278}), .b ({signal_5385, signal_4148}), .c ({signal_5693, signal_4180}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3554 ( .a ({signal_7284, signal_7282}), .b ({signal_5694, signal_4181}), .c ({signal_5800, signal_4213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3555 ( .a ({signal_7288, signal_7286}), .b ({signal_5386, signal_4149}), .c ({signal_5694, signal_4181}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3556 ( .a ({signal_7292, signal_7290}), .b ({signal_5695, signal_4182}), .c ({signal_5801, signal_4214}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3557 ( .a ({signal_7296, signal_7294}), .b ({signal_5387, signal_4150}), .c ({signal_5695, signal_4182}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3558 ( .a ({signal_7300, signal_7298}), .b ({signal_5696, signal_4183}), .c ({signal_5802, signal_4215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3559 ( .a ({signal_7304, signal_7302}), .b ({signal_5365, signal_4151}), .c ({signal_5696, signal_4183}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3560 ( .a ({signal_7308, signal_7306}), .b ({signal_5233, signal_4545}), .c ({signal_5365, signal_4151}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3561 ( .a ({signal_7312, signal_7310}), .b ({signal_5899, signal_4187}), .c ({signal_5988, signal_4219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3562 ( .a ({signal_7316, signal_7314}), .b ({signal_5803, signal_4155}), .c ({signal_5899, signal_4187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3563 ( .a ({signal_7320, signal_7318}), .b ({signal_5711, signal_4123}), .c ({signal_5803, signal_4155}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3564 ( .a ({signal_7324, signal_7322}), .b ({signal_5900, signal_4188}), .c ({signal_5989, signal_4220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3565 ( .a ({signal_7328, signal_7326}), .b ({signal_5804, signal_4156}), .c ({signal_5900, signal_4188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3566 ( .a ({signal_7332, signal_7330}), .b ({signal_5712, signal_4124}), .c ({signal_5804, signal_4156}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3567 ( .a ({signal_7336, signal_7334}), .b ({signal_5805, signal_4216}), .c ({signal_5901, signal_4248}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3568 ( .a ({signal_7340, signal_7338}), .b ({signal_5697, signal_4184}), .c ({signal_5805, signal_4216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3569 ( .a ({signal_7344, signal_7342}), .b ({signal_5366, signal_4152}), .c ({signal_5697, signal_4184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3570 ( .a ({signal_7348, signal_7346}), .b ({signal_5234, signal_4546}), .c ({signal_5366, signal_4152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3571 ( .a ({signal_7352, signal_7350}), .b ({signal_5990, signal_4189}), .c ({signal_6012, signal_4221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3572 ( .a ({signal_7356, signal_7354}), .b ({signal_5902, signal_4157}), .c ({signal_5990, signal_4189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3573 ( .a ({signal_7360, signal_7358}), .b ({signal_5822, signal_4125}), .c ({signal_5902, signal_4157}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3574 ( .a ({signal_7364, signal_7362}), .b ({signal_5903, signal_4190}), .c ({signal_5991, signal_4222}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3575 ( .a ({signal_7368, signal_7366}), .b ({signal_5806, signal_4158}), .c ({signal_5903, signal_4190}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3576 ( .a ({signal_7372, signal_7370}), .b ({signal_5713, signal_4126}), .c ({signal_5806, signal_4158}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3577 ( .a ({signal_7376, signal_7374}), .b ({signal_5992, signal_4191}), .c ({signal_6013, signal_4223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3578 ( .a ({signal_7380, signal_7378}), .b ({signal_5904, signal_4159}), .c ({signal_5992, signal_4191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3579 ( .a ({signal_7384, signal_7382}), .b ({signal_5823, signal_4127}), .c ({signal_5904, signal_4159}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3580 ( .a ({signal_7388, signal_7386}), .b ({signal_5993, signal_4192}), .c ({signal_6014, signal_4224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3581 ( .a ({signal_7392, signal_7390}), .b ({signal_5905, signal_4160}), .c ({signal_5993, signal_4192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3582 ( .a ({signal_7396, signal_7394}), .b ({signal_5824, signal_4128}), .c ({signal_5905, signal_4160}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3583 ( .a ({signal_7400, signal_7398}), .b ({signal_5906, signal_4193}), .c ({signal_5994, signal_4225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3584 ( .a ({signal_7404, signal_7402}), .b ({signal_5807, signal_4161}), .c ({signal_5906, signal_4193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3585 ( .a ({signal_7408, signal_7406}), .b ({signal_5714, signal_4129}), .c ({signal_5807, signal_4161}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3586 ( .a ({signal_7412, signal_7410}), .b ({signal_5907, signal_4194}), .c ({signal_5995, signal_4226}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3587 ( .a ({signal_7416, signal_7414}), .b ({signal_5808, signal_4162}), .c ({signal_5907, signal_4194}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3588 ( .a ({signal_7420, signal_7418}), .b ({signal_5715, signal_4130}), .c ({signal_5808, signal_4162}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3589 ( .a ({signal_7424, signal_7422}), .b ({signal_5809, signal_4195}), .c ({signal_5908, signal_4227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3590 ( .a ({signal_7428, signal_7426}), .b ({signal_5698, signal_4163}), .c ({signal_5809, signal_4195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3591 ( .a ({signal_7432, signal_7430}), .b ({signal_5368, signal_4131}), .c ({signal_5698, signal_4163}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3592 ( .a ({signal_7436, signal_7434}), .b ({signal_5810, signal_4196}), .c ({signal_5909, signal_4228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3593 ( .a ({signal_7440, signal_7438}), .b ({signal_5699, signal_4164}), .c ({signal_5810, signal_4196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3594 ( .a ({signal_7444, signal_7442}), .b ({signal_5369, signal_4132}), .c ({signal_5699, signal_4164}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3595 ( .a ({signal_7448, signal_7446}), .b ({signal_5811, signal_4197}), .c ({signal_5910, signal_4229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3596 ( .a ({signal_7452, signal_7450}), .b ({signal_5700, signal_4165}), .c ({signal_5811, signal_4197}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3597 ( .a ({signal_7456, signal_7454}), .b ({signal_5370, signal_4133}), .c ({signal_5700, signal_4165}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3598 ( .a ({signal_7460, signal_7458}), .b ({signal_5812, signal_4198}), .c ({signal_5911, signal_4230}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3599 ( .a ({signal_7464, signal_7462}), .b ({signal_5701, signal_4166}), .c ({signal_5812, signal_4198}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3600 ( .a ({signal_7468, signal_7466}), .b ({signal_5371, signal_4134}), .c ({signal_5701, signal_4166}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3601 ( .a ({signal_7472, signal_7470}), .b ({signal_5813, signal_4217}), .c ({signal_5912, signal_4249}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3602 ( .a ({signal_7476, signal_7474}), .b ({signal_5702, signal_4185}), .c ({signal_5813, signal_4217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3603 ( .a ({signal_7480, signal_7478}), .b ({signal_5367, signal_4153}), .c ({signal_5702, signal_4185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3604 ( .a ({signal_7484, signal_7482}), .b ({signal_5235, signal_4547}), .c ({signal_5367, signal_4153}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3605 ( .a ({signal_7488, signal_7486}), .b ({signal_5814, signal_4199}), .c ({signal_5913, signal_4231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3606 ( .a ({signal_7492, signal_7490}), .b ({signal_5703, signal_4167}), .c ({signal_5814, signal_4199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3607 ( .a ({signal_7496, signal_7494}), .b ({signal_5372, signal_4135}), .c ({signal_5703, signal_4167}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3608 ( .a ({signal_7500, signal_7498}), .b ({signal_5815, signal_4200}), .c ({signal_5914, signal_4232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3609 ( .a ({signal_7504, signal_7502}), .b ({signal_5704, signal_4168}), .c ({signal_5815, signal_4200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3610 ( .a ({signal_7508, signal_7506}), .b ({signal_5373, signal_4136}), .c ({signal_5704, signal_4168}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3611 ( .a ({signal_7512, signal_7510}), .b ({signal_5816, signal_4201}), .c ({signal_5915, signal_4233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3612 ( .a ({signal_7516, signal_7514}), .b ({signal_5705, signal_4169}), .c ({signal_5816, signal_4201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3613 ( .a ({signal_7520, signal_7518}), .b ({signal_5374, signal_4137}), .c ({signal_5705, signal_4169}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3614 ( .a ({signal_7524, signal_7522}), .b ({signal_5817, signal_4202}), .c ({signal_5916, signal_4234}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3615 ( .a ({signal_7528, signal_7526}), .b ({signal_5706, signal_4170}), .c ({signal_5817, signal_4202}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3616 ( .a ({signal_7532, signal_7530}), .b ({signal_5375, signal_4138}), .c ({signal_5706, signal_4170}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3617 ( .a ({signal_7536, signal_7534}), .b ({signal_5818, signal_4203}), .c ({signal_5917, signal_4235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3618 ( .a ({signal_7540, signal_7538}), .b ({signal_5707, signal_4171}), .c ({signal_5818, signal_4203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3619 ( .a ({signal_7544, signal_7542}), .b ({signal_5376, signal_4139}), .c ({signal_5707, signal_4171}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3620 ( .a ({signal_7548, signal_7546}), .b ({signal_5819, signal_4204}), .c ({signal_5918, signal_4236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3621 ( .a ({signal_7552, signal_7550}), .b ({signal_5708, signal_4172}), .c ({signal_5819, signal_4204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3622 ( .a ({signal_7556, signal_7554}), .b ({signal_5377, signal_4140}), .c ({signal_5708, signal_4172}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3623 ( .a ({signal_7560, signal_7558}), .b ({signal_5820, signal_4205}), .c ({signal_5919, signal_4237}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3624 ( .a ({signal_7564, signal_7562}), .b ({signal_5709, signal_4173}), .c ({signal_5820, signal_4205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3625 ( .a ({signal_7568, signal_7566}), .b ({signal_5378, signal_4141}), .c ({signal_5709, signal_4173}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3626 ( .a ({signal_7572, signal_7570}), .b ({signal_5821, signal_4206}), .c ({signal_5920, signal_4238}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3627 ( .a ({signal_7576, signal_7574}), .b ({signal_5710, signal_4174}), .c ({signal_5821, signal_4206}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3628 ( .a ({signal_7580, signal_7578}), .b ({signal_5379, signal_4142}), .c ({signal_5710, signal_4174}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3629 ( .a ({signal_7584, signal_7582}), .b ({signal_5389, signal_4517}), .c ({signal_5711, signal_4123}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3630 ( .a ({signal_7588, signal_7586}), .b ({signal_5390, signal_4518}), .c ({signal_5712, signal_4124}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3631 ( .a ({signal_7592, signal_7590}), .b ({signal_5719, signal_4519}), .c ({signal_5822, signal_4125}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3632 ( .a ({signal_7596, signal_7594}), .b ({signal_5391, signal_4520}), .c ({signal_5713, signal_4126}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3633 ( .a ({signal_7600, signal_7598}), .b ({signal_5720, signal_4521}), .c ({signal_5823, signal_4127}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3634 ( .a ({signal_7604, signal_7602}), .b ({signal_5721, signal_4522}), .c ({signal_5824, signal_4128}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3635 ( .a ({signal_7608, signal_7606}), .b ({signal_5392, signal_4523}), .c ({signal_5714, signal_4129}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3636 ( .a ({signal_7612, signal_7610}), .b ({signal_5393, signal_4524}), .c ({signal_5715, signal_4130}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3637 ( .a ({signal_7616, signal_7614}), .b ({signal_5825, signal_4207}), .c ({signal_5921, signal_4239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3638 ( .a ({signal_7620, signal_7618}), .b ({signal_5716, signal_4175}), .c ({signal_5825, signal_4207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3639 ( .a ({signal_7624, signal_7622}), .b ({signal_5380, signal_4143}), .c ({signal_5716, signal_4175}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3640 ( .a ({signal_7628, signal_7626}), .b ({signal_5213, signal_4525}), .c ({signal_5368, signal_4131}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3641 ( .a ({signal_7632, signal_7630}), .b ({signal_5214, signal_4526}), .c ({signal_5369, signal_4132}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3642 ( .a ({signal_7636, signal_7634}), .b ({signal_5215, signal_4527}), .c ({signal_5370, signal_4133}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3643 ( .a ({signal_7640, signal_7638}), .b ({signal_5216, signal_4528}), .c ({signal_5371, signal_4134}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3644 ( .a ({signal_7644, signal_7642}), .b ({signal_5217, signal_4529}), .c ({signal_5372, signal_4135}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3645 ( .a ({signal_7648, signal_7646}), .b ({signal_5218, signal_4530}), .c ({signal_5373, signal_4136}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3646 ( .a ({signal_7652, signal_7650}), .b ({signal_5219, signal_4531}), .c ({signal_5374, signal_4137}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3647 ( .a ({signal_7656, signal_7654}), .b ({signal_5220, signal_4532}), .c ({signal_5375, signal_4138}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3648 ( .a ({signal_7660, signal_7658}), .b ({signal_5221, signal_4533}), .c ({signal_5376, signal_4139}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3649 ( .a ({signal_7664, signal_7662}), .b ({signal_5222, signal_4534}), .c ({signal_5377, signal_4140}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3650 ( .a ({signal_7668, signal_7666}), .b ({signal_5826, signal_4208}), .c ({signal_5922, signal_4240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3651 ( .a ({signal_7672, signal_7670}), .b ({signal_5717, signal_4176}), .c ({signal_5826, signal_4208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3652 ( .a ({signal_7676, signal_7674}), .b ({signal_5381, signal_4144}), .c ({signal_5717, signal_4176}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3653 ( .a ({signal_7680, signal_7678}), .b ({signal_5223, signal_4535}), .c ({signal_5378, signal_4141}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3654 ( .a ({signal_7684, signal_7682}), .b ({signal_5224, signal_4536}), .c ({signal_5379, signal_4142}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3655 ( .a ({signal_7688, signal_7686}), .b ({signal_5225, signal_4537}), .c ({signal_5380, signal_4143}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3656 ( .a ({signal_7692, signal_7690}), .b ({signal_5226, signal_4538}), .c ({signal_5381, signal_4144}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3657 ( .a ({signal_7696, signal_7694}), .b ({signal_5227, signal_4539}), .c ({signal_5382, signal_4145}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3658 ( .a ({signal_7700, signal_7698}), .b ({signal_5228, signal_4540}), .c ({signal_5383, signal_4146}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3659 ( .a ({signal_7704, signal_7702}), .b ({signal_5229, signal_4541}), .c ({signal_5384, signal_4147}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3660 ( .a ({signal_7708, signal_7706}), .b ({signal_5230, signal_4542}), .c ({signal_5385, signal_4148}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3661 ( .a ({signal_7712, signal_7710}), .b ({signal_5231, signal_4543}), .c ({signal_5386, signal_4149}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3662 ( .a ({signal_7716, signal_7714}), .b ({signal_5232, signal_4544}), .c ({signal_5387, signal_4150}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3663 ( .a ({signal_7720, signal_7718}), .b ({signal_5827, signal_4218}), .c ({signal_5923, signal_4250}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3664 ( .a ({signal_7724, signal_7722}), .b ({signal_5718, signal_4186}), .c ({signal_5827, signal_4218}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3665 ( .a ({signal_7728, signal_7726}), .b ({signal_5388, signal_4154}), .c ({signal_5718, signal_4186}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3666 ( .a ({signal_7732, signal_7730}), .b ({signal_5236, signal_4548}), .c ({signal_5388, signal_4154}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3667 ( .a ({signal_4964, signal_3116}), .b ({1'b0, signal_7734}), .c ({signal_5389, signal_4517}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3668 ( .a ({signal_4963, signal_3115}), .b ({1'b0, signal_7736}), .c ({signal_5390, signal_4518}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3669 ( .a ({signal_4962, signal_3114}), .b ({1'b0, signal_7738}), .c ({signal_5719, signal_4519}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3670 ( .a ({signal_4961, signal_3113}), .b ({1'b0, signal_7740}), .c ({signal_5391, signal_4520}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3671 ( .a ({signal_4960, signal_3112}), .b ({1'b0, signal_7742}), .c ({signal_5720, signal_4521}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3672 ( .a ({signal_4959, signal_3111}), .b ({1'b0, signal_7744}), .c ({signal_5721, signal_4522}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3673 ( .a ({signal_4958, signal_3110}), .b ({1'b0, signal_7746}), .c ({signal_5392, signal_4523}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3674 ( .a ({signal_4957, signal_3109}), .b ({1'b0, signal_7748}), .c ({signal_5393, signal_4524}) ) ;
    AES_step2_ANF #(.low_latency(0), .pipeline(1)) cell_4209 ( .in0 ({signal_912, signal_792, signal_4378, signal_4377, signal_4376, signal_4375, signal_4374, signal_4373, signal_4372, signal_4371, signal_4370, signal_4369, signal_4368, signal_4367, signal_4366, signal_4365, signal_4364, signal_4363, signal_4362, signal_4361, signal_4360, signal_4359, signal_4358, signal_4357, signal_4356, signal_4355, signal_4354, signal_4353, signal_4352, signal_4351, signal_4350, signal_4349, signal_4348, signal_4347, ciphertext_s0[0], ciphertext_s0[1], ciphertext_s0[2], ciphertext_s0[4], ciphertext_s0[5], ciphertext_s0[6], ciphertext_s0[7], ciphertext_s0[8], ciphertext_s0[9], ciphertext_s0[10], ciphertext_s0[12], ciphertext_s0[13], ciphertext_s0[14], ciphertext_s0[15], ciphertext_s0[16], ciphertext_s0[17], ciphertext_s0[18], ciphertext_s0[20], ciphertext_s0[21], ciphertext_s0[22], ciphertext_s0[23], ciphertext_s0[24], ciphertext_s0[25], ciphertext_s0[26], ciphertext_s0[28], ciphertext_s0[29], ciphertext_s0[30], ciphertext_s0[31], ciphertext_s0[32], ciphertext_s0[33], ciphertext_s0[34], ciphertext_s0[36], ciphertext_s0[37], ciphertext_s0[38], ciphertext_s0[39], ciphertext_s0[40], ciphertext_s0[41], ciphertext_s0[42], ciphertext_s0[44], ciphertext_s0[45], ciphertext_s0[46], ciphertext_s0[47], ciphertext_s0[48], ciphertext_s0[49], ciphertext_s0[50], ciphertext_s0[52], ciphertext_s0[53], ciphertext_s0[54], ciphertext_s0[55], ciphertext_s0[56], ciphertext_s0[57], ciphertext_s0[58], ciphertext_s0[60], ciphertext_s0[61], ciphertext_s0[62], ciphertext_s0[63], ciphertext_s0[64], ciphertext_s0[65], ciphertext_s0[66], ciphertext_s0[68], ciphertext_s0[69], ciphertext_s0[70], ciphertext_s0[71], ciphertext_s0[72], ciphertext_s0[73], ciphertext_s0[74], ciphertext_s0[76], ciphertext_s0[77], ciphertext_s0[78], ciphertext_s0[79], ciphertext_s0[80], ciphertext_s0[81], ciphertext_s0[82], ciphertext_s0[84], ciphertext_s0[85], ciphertext_s0[86], ciphertext_s0[87], ciphertext_s0[88], ciphertext_s0[89], ciphertext_s0[90], ciphertext_s0[92], ciphertext_s0[93], ciphertext_s0[94], ciphertext_s0[95], ciphertext_s0[96], ciphertext_s0[97], ciphertext_s0[98], ciphertext_s0[100], ciphertext_s0[101], ciphertext_s0[102], ciphertext_s0[103], ciphertext_s0[104], ciphertext_s0[105], ciphertext_s0[106], ciphertext_s0[108], ciphertext_s0[109], ciphertext_s0[110], ciphertext_s0[111], ciphertext_s0[112], ciphertext_s0[113], ciphertext_s0[114], ciphertext_s0[116], ciphertext_s0[117], ciphertext_s0[118], ciphertext_s0[119], ciphertext_s0[120], ciphertext_s0[121], ciphertext_s0[122], ciphertext_s0[124], ciphertext_s0[125], ciphertext_s0[126], ciphertext_s0[127], signal_2592, signal_2472, signal_2352, signal_2232, signal_2112, signal_1992, signal_1872, signal_1752, signal_1632, signal_1512, signal_1392, signal_1272, signal_1152, signal_1032}), .in1 ({signal_4934, signal_4933, signal_4550, signal_4667, signal_4700, signal_4733, signal_4766, signal_4799, signal_4832, signal_4865, signal_4898, signal_4931, signal_4583, signal_4616, signal_4643, signal_4646, signal_4649, signal_4652, signal_4655, signal_4658, signal_4661, signal_4664, signal_4670, signal_4673, signal_4676, signal_4679, signal_4682, signal_4685, signal_4688, signal_4691, signal_4694, signal_4697, signal_4703, signal_4706, ciphertext_s1[0], ciphertext_s1[1], ciphertext_s1[2], ciphertext_s1[4], ciphertext_s1[5], ciphertext_s1[6], ciphertext_s1[7], ciphertext_s1[8], ciphertext_s1[9], ciphertext_s1[10], ciphertext_s1[12], ciphertext_s1[13], ciphertext_s1[14], ciphertext_s1[15], ciphertext_s1[16], ciphertext_s1[17], ciphertext_s1[18], ciphertext_s1[20], ciphertext_s1[21], ciphertext_s1[22], ciphertext_s1[23], ciphertext_s1[24], ciphertext_s1[25], ciphertext_s1[26], ciphertext_s1[28], ciphertext_s1[29], ciphertext_s1[30], ciphertext_s1[31], ciphertext_s1[32], ciphertext_s1[33], ciphertext_s1[34], ciphertext_s1[36], ciphertext_s1[37], ciphertext_s1[38], ciphertext_s1[39], ciphertext_s1[40], ciphertext_s1[41], ciphertext_s1[42], ciphertext_s1[44], ciphertext_s1[45], ciphertext_s1[46], ciphertext_s1[47], ciphertext_s1[48], ciphertext_s1[49], ciphertext_s1[50], ciphertext_s1[52], ciphertext_s1[53], ciphertext_s1[54], ciphertext_s1[55], ciphertext_s1[56], ciphertext_s1[57], ciphertext_s1[58], ciphertext_s1[60], ciphertext_s1[61], ciphertext_s1[62], ciphertext_s1[63], ciphertext_s1[64], ciphertext_s1[65], ciphertext_s1[66], ciphertext_s1[68], ciphertext_s1[69], ciphertext_s1[70], ciphertext_s1[71], ciphertext_s1[72], ciphertext_s1[73], ciphertext_s1[74], ciphertext_s1[76], ciphertext_s1[77], ciphertext_s1[78], ciphertext_s1[79], ciphertext_s1[80], ciphertext_s1[81], ciphertext_s1[82], ciphertext_s1[84], ciphertext_s1[85], ciphertext_s1[86], ciphertext_s1[87], ciphertext_s1[88], ciphertext_s1[89], ciphertext_s1[90], ciphertext_s1[92], ciphertext_s1[93], ciphertext_s1[94], ciphertext_s1[95], ciphertext_s1[96], ciphertext_s1[97], ciphertext_s1[98], ciphertext_s1[100], ciphertext_s1[101], ciphertext_s1[102], ciphertext_s1[103], ciphertext_s1[104], ciphertext_s1[105], ciphertext_s1[106], ciphertext_s1[108], ciphertext_s1[109], ciphertext_s1[110], ciphertext_s1[111], ciphertext_s1[112], ciphertext_s1[113], ciphertext_s1[114], ciphertext_s1[116], ciphertext_s1[117], ciphertext_s1[118], ciphertext_s1[119], ciphertext_s1[120], ciphertext_s1[121], ciphertext_s1[122], ciphertext_s1[124], ciphertext_s1[125], ciphertext_s1[126], ciphertext_s1[127], signal_4948, signal_4947, signal_4946, signal_4945, signal_4944, signal_4943, signal_4942, signal_4941, signal_4940, signal_4939, signal_4938, signal_4937, signal_4936, signal_4935}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_4548, signal_4547, signal_4546, signal_4545, signal_4544, signal_4543, signal_4542, signal_4541, signal_4540, signal_4539, signal_4538, signal_4537, signal_4536, signal_4535, signal_4534, signal_4533, signal_4532, signal_4531, signal_4530, signal_4529, signal_4528, signal_4527, signal_4526, signal_4525, signal_4516, signal_4514, signal_4511, signal_4510, signal_4509, signal_4508, signal_4506, signal_4503, signal_4502, signal_4501, signal_4500, signal_4498, signal_4495, signal_4494, signal_4493, signal_4492, signal_4490, signal_4487, signal_4486, signal_4485, signal_4484, signal_4482, signal_4479, signal_4478, signal_4477, signal_4476, signal_4474, signal_4471, signal_4470, signal_4469, signal_4468, signal_4466, signal_4463, signal_4462, signal_4461, signal_4460, signal_4458, signal_4455, signal_4454, signal_4453, signal_4452, signal_4450, signal_4447, signal_4446, signal_4445, signal_4444, signal_4442, signal_4439, signal_4438, signal_4437, signal_4436, signal_4434, signal_4431, signal_4430, signal_4429, signal_4428, signal_4426, signal_4423, signal_4422, signal_4421, signal_4420, signal_4418, signal_4415, signal_4414, signal_4413, signal_4412, signal_4410, signal_4407, signal_4406, signal_4405, signal_4404, signal_4402, signal_4399, signal_4398, signal_4397, signal_4396, signal_4394, signal_4391, signal_4390, signal_4389, signal_4121, signal_4120, signal_4119, signal_4118, signal_4117, signal_4116, signal_4115, signal_4114, signal_4112, signal_4111, signal_4110, signal_4109, signal_4108, signal_4107, signal_4106, signal_4105, signal_4104, signal_4103, signal_4102, signal_4101, signal_4100, signal_4099, signal_4098, signal_4097, signal_4096, signal_4095, signal_4094, signal_4093, signal_4092, signal_4091, signal_4089, signal_4088, signal_4087, signal_4086, signal_4085, signal_4084, signal_4083, signal_4082, signal_4080, signal_4079, signal_4078, signal_4077, signal_4076, signal_4075, signal_4074, signal_4073, signal_4072, signal_4071, signal_4070, signal_4069, signal_4068, signal_4067, signal_4066, signal_4065, signal_4064, signal_4063, signal_4062, signal_4061, signal_4060, signal_4059, signal_4057, signal_4056, signal_4055, signal_4054, signal_4053, signal_4052, signal_4051, signal_4050, signal_4048, signal_4047, signal_4046, signal_4045, signal_4044, signal_4043, signal_4042, signal_4041, signal_4040, signal_4039, signal_4038, signal_4037, signal_4036, signal_4035, signal_4034, signal_4033, signal_4032, signal_4031, signal_4030, signal_4029, signal_4028, signal_4027, signal_4025, signal_4024, signal_4023, signal_4022, signal_4021, signal_4020, signal_4019, signal_4018, signal_4016, signal_4015, signal_4014, signal_4013, signal_4012, signal_4011, signal_4010, signal_4009, signal_4008, signal_4007, signal_4006, signal_4005, signal_4004, signal_4003, signal_4002, signal_4001, signal_4000, signal_3999, signal_3998, signal_3997, signal_3996, signal_3995, signal_3994, signal_3992, signal_3991, signal_3986, signal_3984, signal_3983, signal_3978, signal_3976, signal_3975, signal_3970, signal_3968, signal_3967, signal_3962, signal_3960, signal_3959, signal_3954, signal_3952, signal_3951, signal_3946, signal_3944, signal_3943, signal_3938, signal_3936, signal_3935, signal_3930, signal_3928, signal_3927, signal_3922, signal_3920, signal_3919, signal_3914, signal_3912, signal_3911, signal_3906, signal_3904, signal_3903, signal_3898, signal_3896, signal_3895, signal_3890, signal_3888, signal_3887, signal_3882, signal_3880, signal_3879, signal_3874, signal_3872, signal_3871, signal_3116, signal_3115, signal_3114, signal_3113, signal_3112, signal_3111, signal_3110, signal_3109, signal_2852, signal_2789, signal_2788, signal_2725, signal_2724, signal_2661, signal_2660, signal_2597}), .out1 ({signal_5236, signal_5235, signal_5234, signal_5233, signal_5232, signal_5231, signal_5230, signal_5229, signal_5228, signal_5227, signal_5226, signal_5225, signal_5224, signal_5223, signal_5222, signal_5221, signal_5220, signal_5219, signal_5218, signal_5217, signal_5216, signal_5215, signal_5214, signal_5213, signal_5212, signal_5211, signal_5210, signal_5209, signal_5208, signal_5207, signal_5206, signal_5205, signal_5204, signal_5203, signal_5202, signal_5201, signal_5200, signal_5199, signal_5198, signal_5197, signal_5196, signal_5195, signal_5194, signal_5193, signal_5192, signal_5191, signal_5190, signal_5189, signal_5188, signal_5187, signal_5186, signal_5185, signal_5184, signal_5183, signal_5182, signal_5181, signal_5180, signal_5179, signal_5178, signal_5177, signal_5176, signal_5175, signal_5174, signal_5173, signal_5172, signal_5171, signal_5170, signal_5169, signal_5168, signal_5167, signal_5166, signal_5165, signal_5164, signal_5163, signal_5162, signal_5161, signal_5160, signal_5159, signal_5158, signal_5157, signal_5156, signal_5155, signal_5154, signal_5153, signal_5152, signal_5151, signal_5150, signal_5149, signal_5148, signal_5147, signal_5146, signal_5145, signal_5144, signal_5143, signal_5142, signal_5141, signal_5140, signal_5139, signal_5138, signal_5137, signal_5136, signal_5135, signal_5134, signal_5133, signal_5132, signal_5131, signal_5130, signal_5129, signal_5128, signal_5127, signal_5126, signal_5125, signal_5124, signal_5123, signal_5122, signal_5121, signal_5120, signal_5119, signal_5118, signal_5117, signal_5116, signal_5115, signal_5114, signal_5113, signal_5112, signal_5111, signal_5110, signal_5109, signal_5108, signal_5107, signal_5106, signal_5105, signal_5104, signal_5103, signal_5102, signal_5101, signal_5100, signal_5099, signal_5098, signal_5097, signal_5096, signal_5095, signal_5094, signal_5093, signal_5092, signal_5091, signal_5090, signal_5089, signal_5088, signal_5087, signal_5086, signal_5085, signal_5084, signal_5083, signal_5082, signal_5081, signal_5080, signal_5079, signal_5078, signal_5077, signal_5076, signal_5075, signal_5074, signal_5073, signal_5072, signal_5071, signal_5070, signal_5069, signal_5068, signal_5067, signal_5066, signal_5065, signal_5064, signal_5063, signal_5062, signal_5061, signal_5060, signal_5059, signal_5058, signal_5057, signal_5056, signal_5055, signal_5054, signal_5053, signal_5052, signal_5051, signal_5050, signal_5049, signal_5048, signal_5047, signal_5046, signal_5045, signal_5044, signal_5043, signal_5042, signal_5041, signal_5040, signal_5039, signal_5038, signal_5037, signal_5036, signal_5035, signal_5034, signal_5033, signal_5032, signal_5031, signal_5030, signal_5029, signal_5028, signal_5027, signal_5026, signal_5025, signal_5024, signal_5023, signal_5022, signal_5021, signal_5020, signal_5019, signal_5018, signal_5017, signal_5016, signal_5015, signal_5014, signal_5013, signal_5012, signal_5011, signal_5010, signal_5009, signal_5008, signal_5007, signal_5006, signal_5005, signal_5004, signal_5003, signal_5002, signal_5001, signal_5000, signal_4999, signal_4998, signal_4997, signal_4996, signal_4995, signal_4994, signal_4993, signal_4992, signal_4991, signal_4990, signal_4989, signal_4988, signal_4987, signal_4986, signal_4985, signal_4984, signal_4983, signal_4982, signal_4981, signal_4980, signal_4979, signal_4978, signal_4977, signal_4976, signal_4975, signal_4974, signal_4973, signal_4972, signal_4971, signal_4970, signal_4969, signal_4968, signal_4967, signal_4966, signal_4965, signal_4964, signal_4963, signal_4962, signal_4961, signal_4960, signal_4959, signal_4958, signal_4957, signal_4956, signal_4955, signal_4954, signal_4953, signal_4952, signal_4951, signal_4950, signal_4949}) ) ;
    buf_clk cell_4211 ( .C (clk), .D (signal_6181), .Q (signal_6182) ) ;
    buf_clk cell_4213 ( .C (clk), .D (signal_6183), .Q (signal_6184) ) ;
    buf_clk cell_4215 ( .C (clk), .D (signal_6185), .Q (signal_6186) ) ;
    buf_clk cell_4217 ( .C (clk), .D (signal_6187), .Q (signal_6188) ) ;
    buf_clk cell_4219 ( .C (clk), .D (signal_6189), .Q (signal_6190) ) ;
    buf_clk cell_4221 ( .C (clk), .D (signal_6191), .Q (signal_6192) ) ;
    buf_clk cell_4223 ( .C (clk), .D (signal_6193), .Q (signal_6194) ) ;
    buf_clk cell_4225 ( .C (clk), .D (signal_6195), .Q (signal_6196) ) ;
    buf_clk cell_4227 ( .C (clk), .D (signal_6197), .Q (signal_6198) ) ;
    buf_clk cell_4229 ( .C (clk), .D (signal_6199), .Q (signal_6200) ) ;
    buf_clk cell_4231 ( .C (clk), .D (signal_6201), .Q (signal_6202) ) ;
    buf_clk cell_4233 ( .C (clk), .D (signal_6203), .Q (signal_6204) ) ;
    buf_clk cell_4235 ( .C (clk), .D (signal_6205), .Q (signal_6206) ) ;
    buf_clk cell_4237 ( .C (clk), .D (signal_6207), .Q (signal_6208) ) ;
    buf_clk cell_4239 ( .C (clk), .D (signal_6209), .Q (signal_6210) ) ;
    buf_clk cell_4241 ( .C (clk), .D (signal_6211), .Q (signal_6212) ) ;
    buf_clk cell_4243 ( .C (clk), .D (signal_6213), .Q (signal_6214) ) ;
    buf_clk cell_4245 ( .C (clk), .D (signal_6215), .Q (signal_6216) ) ;
    buf_clk cell_4247 ( .C (clk), .D (signal_6217), .Q (signal_6218) ) ;
    buf_clk cell_4249 ( .C (clk), .D (signal_6219), .Q (signal_6220) ) ;
    buf_clk cell_4251 ( .C (clk), .D (signal_6221), .Q (signal_6222) ) ;
    buf_clk cell_4253 ( .C (clk), .D (signal_6223), .Q (signal_6224) ) ;
    buf_clk cell_4255 ( .C (clk), .D (signal_6225), .Q (signal_6226) ) ;
    buf_clk cell_4257 ( .C (clk), .D (signal_6227), .Q (signal_6228) ) ;
    buf_clk cell_4259 ( .C (clk), .D (signal_6229), .Q (signal_6230) ) ;
    buf_clk cell_4261 ( .C (clk), .D (signal_6231), .Q (signal_6232) ) ;
    buf_clk cell_4263 ( .C (clk), .D (signal_6233), .Q (signal_6234) ) ;
    buf_clk cell_4265 ( .C (clk), .D (signal_6235), .Q (signal_6236) ) ;
    buf_clk cell_4267 ( .C (clk), .D (signal_6237), .Q (signal_6238) ) ;
    buf_clk cell_4269 ( .C (clk), .D (signal_6239), .Q (signal_6240) ) ;
    buf_clk cell_4271 ( .C (clk), .D (signal_6241), .Q (signal_6242) ) ;
    buf_clk cell_4273 ( .C (clk), .D (signal_6243), .Q (signal_6244) ) ;
    buf_clk cell_4275 ( .C (clk), .D (signal_6245), .Q (signal_6246) ) ;
    buf_clk cell_4277 ( .C (clk), .D (signal_6247), .Q (signal_6248) ) ;
    buf_clk cell_4279 ( .C (clk), .D (signal_6249), .Q (signal_6250) ) ;
    buf_clk cell_4281 ( .C (clk), .D (signal_6251), .Q (signal_6252) ) ;
    buf_clk cell_4283 ( .C (clk), .D (signal_6253), .Q (signal_6254) ) ;
    buf_clk cell_4285 ( .C (clk), .D (signal_6255), .Q (signal_6256) ) ;
    buf_clk cell_4287 ( .C (clk), .D (signal_6257), .Q (signal_6258) ) ;
    buf_clk cell_4289 ( .C (clk), .D (signal_6259), .Q (signal_6260) ) ;
    buf_clk cell_4291 ( .C (clk), .D (signal_6261), .Q (signal_6262) ) ;
    buf_clk cell_4293 ( .C (clk), .D (signal_6263), .Q (signal_6264) ) ;
    buf_clk cell_4295 ( .C (clk), .D (signal_6265), .Q (signal_6266) ) ;
    buf_clk cell_4297 ( .C (clk), .D (signal_6267), .Q (signal_6268) ) ;
    buf_clk cell_4299 ( .C (clk), .D (signal_6269), .Q (signal_6270) ) ;
    buf_clk cell_4301 ( .C (clk), .D (signal_6271), .Q (signal_6272) ) ;
    buf_clk cell_4303 ( .C (clk), .D (signal_6273), .Q (signal_6274) ) ;
    buf_clk cell_4305 ( .C (clk), .D (signal_6275), .Q (signal_6276) ) ;
    buf_clk cell_4307 ( .C (clk), .D (signal_6277), .Q (signal_6278) ) ;
    buf_clk cell_4309 ( .C (clk), .D (signal_6279), .Q (signal_6280) ) ;
    buf_clk cell_4311 ( .C (clk), .D (signal_6281), .Q (signal_6282) ) ;
    buf_clk cell_4313 ( .C (clk), .D (signal_6283), .Q (signal_6284) ) ;
    buf_clk cell_4315 ( .C (clk), .D (signal_6285), .Q (signal_6286) ) ;
    buf_clk cell_4317 ( .C (clk), .D (signal_6287), .Q (signal_6288) ) ;
    buf_clk cell_4319 ( .C (clk), .D (signal_6289), .Q (signal_6290) ) ;
    buf_clk cell_4321 ( .C (clk), .D (signal_6291), .Q (signal_6292) ) ;
    buf_clk cell_4323 ( .C (clk), .D (signal_6293), .Q (signal_6294) ) ;
    buf_clk cell_4325 ( .C (clk), .D (signal_6295), .Q (signal_6296) ) ;
    buf_clk cell_4327 ( .C (clk), .D (signal_6297), .Q (signal_6298) ) ;
    buf_clk cell_4329 ( .C (clk), .D (signal_6299), .Q (signal_6300) ) ;
    buf_clk cell_4331 ( .C (clk), .D (signal_6301), .Q (signal_6302) ) ;
    buf_clk cell_4333 ( .C (clk), .D (signal_6303), .Q (signal_6304) ) ;
    buf_clk cell_4335 ( .C (clk), .D (signal_6305), .Q (signal_6306) ) ;
    buf_clk cell_4337 ( .C (clk), .D (signal_6307), .Q (signal_6308) ) ;
    buf_clk cell_4339 ( .C (clk), .D (signal_6309), .Q (signal_6310) ) ;
    buf_clk cell_4341 ( .C (clk), .D (signal_6311), .Q (signal_6312) ) ;
    buf_clk cell_4343 ( .C (clk), .D (signal_6313), .Q (signal_6314) ) ;
    buf_clk cell_4345 ( .C (clk), .D (signal_6315), .Q (signal_6316) ) ;
    buf_clk cell_4347 ( .C (clk), .D (signal_6317), .Q (signal_6318) ) ;
    buf_clk cell_4349 ( .C (clk), .D (signal_6319), .Q (signal_6320) ) ;
    buf_clk cell_4351 ( .C (clk), .D (signal_6321), .Q (signal_6322) ) ;
    buf_clk cell_4353 ( .C (clk), .D (signal_6323), .Q (signal_6324) ) ;
    buf_clk cell_4355 ( .C (clk), .D (signal_6325), .Q (signal_6326) ) ;
    buf_clk cell_4357 ( .C (clk), .D (signal_6327), .Q (signal_6328) ) ;
    buf_clk cell_4359 ( .C (clk), .D (signal_6329), .Q (signal_6330) ) ;
    buf_clk cell_4361 ( .C (clk), .D (signal_6331), .Q (signal_6332) ) ;
    buf_clk cell_4363 ( .C (clk), .D (signal_6333), .Q (signal_6334) ) ;
    buf_clk cell_4365 ( .C (clk), .D (signal_6335), .Q (signal_6336) ) ;
    buf_clk cell_4367 ( .C (clk), .D (signal_6337), .Q (signal_6338) ) ;
    buf_clk cell_4369 ( .C (clk), .D (signal_6339), .Q (signal_6340) ) ;
    buf_clk cell_4371 ( .C (clk), .D (signal_6341), .Q (signal_6342) ) ;
    buf_clk cell_4373 ( .C (clk), .D (signal_6343), .Q (signal_6344) ) ;
    buf_clk cell_4375 ( .C (clk), .D (signal_6345), .Q (signal_6346) ) ;
    buf_clk cell_4377 ( .C (clk), .D (signal_6347), .Q (signal_6348) ) ;
    buf_clk cell_4379 ( .C (clk), .D (signal_6349), .Q (signal_6350) ) ;
    buf_clk cell_4381 ( .C (clk), .D (signal_6351), .Q (signal_6352) ) ;
    buf_clk cell_4383 ( .C (clk), .D (signal_6353), .Q (signal_6354) ) ;
    buf_clk cell_4385 ( .C (clk), .D (signal_6355), .Q (signal_6356) ) ;
    buf_clk cell_4387 ( .C (clk), .D (signal_6357), .Q (signal_6358) ) ;
    buf_clk cell_4389 ( .C (clk), .D (signal_6359), .Q (signal_6360) ) ;
    buf_clk cell_4391 ( .C (clk), .D (signal_6361), .Q (signal_6362) ) ;
    buf_clk cell_4393 ( .C (clk), .D (signal_6363), .Q (signal_6364) ) ;
    buf_clk cell_4395 ( .C (clk), .D (signal_6365), .Q (signal_6366) ) ;
    buf_clk cell_4397 ( .C (clk), .D (signal_6367), .Q (signal_6368) ) ;
    buf_clk cell_4399 ( .C (clk), .D (signal_6369), .Q (signal_6370) ) ;
    buf_clk cell_4401 ( .C (clk), .D (signal_6371), .Q (signal_6372) ) ;
    buf_clk cell_4403 ( .C (clk), .D (signal_6373), .Q (signal_6374) ) ;
    buf_clk cell_4405 ( .C (clk), .D (signal_6375), .Q (signal_6376) ) ;
    buf_clk cell_4407 ( .C (clk), .D (signal_6377), .Q (signal_6378) ) ;
    buf_clk cell_4409 ( .C (clk), .D (signal_6379), .Q (signal_6380) ) ;
    buf_clk cell_4411 ( .C (clk), .D (signal_6381), .Q (signal_6382) ) ;
    buf_clk cell_4413 ( .C (clk), .D (signal_6383), .Q (signal_6384) ) ;
    buf_clk cell_4415 ( .C (clk), .D (signal_6385), .Q (signal_6386) ) ;
    buf_clk cell_4417 ( .C (clk), .D (signal_6387), .Q (signal_6388) ) ;
    buf_clk cell_4419 ( .C (clk), .D (signal_6389), .Q (signal_6390) ) ;
    buf_clk cell_4421 ( .C (clk), .D (signal_6391), .Q (signal_6392) ) ;
    buf_clk cell_4423 ( .C (clk), .D (signal_6393), .Q (signal_6394) ) ;
    buf_clk cell_4425 ( .C (clk), .D (signal_6395), .Q (signal_6396) ) ;
    buf_clk cell_4427 ( .C (clk), .D (signal_6397), .Q (signal_6398) ) ;
    buf_clk cell_4429 ( .C (clk), .D (signal_6399), .Q (signal_6400) ) ;
    buf_clk cell_4431 ( .C (clk), .D (signal_6401), .Q (signal_6402) ) ;
    buf_clk cell_4433 ( .C (clk), .D (signal_6403), .Q (signal_6404) ) ;
    buf_clk cell_4435 ( .C (clk), .D (signal_6405), .Q (signal_6406) ) ;
    buf_clk cell_4437 ( .C (clk), .D (signal_6407), .Q (signal_6408) ) ;
    buf_clk cell_4439 ( .C (clk), .D (signal_6409), .Q (signal_6410) ) ;
    buf_clk cell_4441 ( .C (clk), .D (signal_6411), .Q (signal_6412) ) ;
    buf_clk cell_4443 ( .C (clk), .D (signal_6413), .Q (signal_6414) ) ;
    buf_clk cell_4445 ( .C (clk), .D (signal_6415), .Q (signal_6416) ) ;
    buf_clk cell_4447 ( .C (clk), .D (signal_6417), .Q (signal_6418) ) ;
    buf_clk cell_4449 ( .C (clk), .D (signal_6419), .Q (signal_6420) ) ;
    buf_clk cell_4451 ( .C (clk), .D (signal_6421), .Q (signal_6422) ) ;
    buf_clk cell_4453 ( .C (clk), .D (signal_6423), .Q (signal_6424) ) ;
    buf_clk cell_4455 ( .C (clk), .D (signal_6425), .Q (signal_6426) ) ;
    buf_clk cell_4457 ( .C (clk), .D (signal_6427), .Q (signal_6428) ) ;
    buf_clk cell_4459 ( .C (clk), .D (signal_6429), .Q (signal_6430) ) ;
    buf_clk cell_4461 ( .C (clk), .D (signal_6431), .Q (signal_6432) ) ;
    buf_clk cell_4463 ( .C (clk), .D (signal_6433), .Q (signal_6434) ) ;
    buf_clk cell_4465 ( .C (clk), .D (signal_6435), .Q (signal_6436) ) ;
    buf_clk cell_4467 ( .C (clk), .D (signal_6437), .Q (signal_6438) ) ;
    buf_clk cell_4469 ( .C (clk), .D (signal_6439), .Q (signal_6440) ) ;
    buf_clk cell_4471 ( .C (clk), .D (signal_6441), .Q (signal_6442) ) ;
    buf_clk cell_4473 ( .C (clk), .D (signal_6443), .Q (signal_6444) ) ;
    buf_clk cell_4475 ( .C (clk), .D (signal_6445), .Q (signal_6446) ) ;
    buf_clk cell_4477 ( .C (clk), .D (signal_6447), .Q (signal_6448) ) ;
    buf_clk cell_4479 ( .C (clk), .D (signal_6449), .Q (signal_6450) ) ;
    buf_clk cell_4481 ( .C (clk), .D (signal_6451), .Q (signal_6452) ) ;
    buf_clk cell_4483 ( .C (clk), .D (signal_6453), .Q (signal_6454) ) ;
    buf_clk cell_4485 ( .C (clk), .D (signal_6455), .Q (signal_6456) ) ;
    buf_clk cell_4487 ( .C (clk), .D (signal_6457), .Q (signal_6458) ) ;
    buf_clk cell_4489 ( .C (clk), .D (signal_6459), .Q (signal_6460) ) ;
    buf_clk cell_4491 ( .C (clk), .D (signal_6461), .Q (signal_6462) ) ;
    buf_clk cell_4493 ( .C (clk), .D (signal_6463), .Q (signal_6464) ) ;
    buf_clk cell_4495 ( .C (clk), .D (signal_6465), .Q (signal_6466) ) ;
    buf_clk cell_4497 ( .C (clk), .D (signal_6467), .Q (signal_6468) ) ;
    buf_clk cell_4499 ( .C (clk), .D (signal_6469), .Q (signal_6470) ) ;
    buf_clk cell_4501 ( .C (clk), .D (signal_6471), .Q (signal_6472) ) ;
    buf_clk cell_4503 ( .C (clk), .D (signal_6473), .Q (signal_6474) ) ;
    buf_clk cell_4505 ( .C (clk), .D (signal_6475), .Q (signal_6476) ) ;
    buf_clk cell_4507 ( .C (clk), .D (signal_6477), .Q (signal_6478) ) ;
    buf_clk cell_4509 ( .C (clk), .D (signal_6479), .Q (signal_6480) ) ;
    buf_clk cell_4511 ( .C (clk), .D (signal_6481), .Q (signal_6482) ) ;
    buf_clk cell_4513 ( .C (clk), .D (signal_6483), .Q (signal_6484) ) ;
    buf_clk cell_4515 ( .C (clk), .D (signal_6485), .Q (signal_6486) ) ;
    buf_clk cell_4517 ( .C (clk), .D (signal_6487), .Q (signal_6488) ) ;
    buf_clk cell_4519 ( .C (clk), .D (signal_6489), .Q (signal_6490) ) ;
    buf_clk cell_4521 ( .C (clk), .D (signal_6491), .Q (signal_6492) ) ;
    buf_clk cell_4523 ( .C (clk), .D (signal_6493), .Q (signal_6494) ) ;
    buf_clk cell_4525 ( .C (clk), .D (signal_6495), .Q (signal_6496) ) ;
    buf_clk cell_4527 ( .C (clk), .D (signal_6497), .Q (signal_6498) ) ;
    buf_clk cell_4529 ( .C (clk), .D (signal_6499), .Q (signal_6500) ) ;
    buf_clk cell_4531 ( .C (clk), .D (signal_6501), .Q (signal_6502) ) ;
    buf_clk cell_4533 ( .C (clk), .D (signal_6503), .Q (signal_6504) ) ;
    buf_clk cell_4535 ( .C (clk), .D (signal_6505), .Q (signal_6506) ) ;
    buf_clk cell_4537 ( .C (clk), .D (signal_6507), .Q (signal_6508) ) ;
    buf_clk cell_4539 ( .C (clk), .D (signal_6509), .Q (signal_6510) ) ;
    buf_clk cell_4541 ( .C (clk), .D (signal_6511), .Q (signal_6512) ) ;
    buf_clk cell_4543 ( .C (clk), .D (signal_6513), .Q (signal_6514) ) ;
    buf_clk cell_4545 ( .C (clk), .D (signal_6515), .Q (signal_6516) ) ;
    buf_clk cell_4547 ( .C (clk), .D (signal_6517), .Q (signal_6518) ) ;
    buf_clk cell_4549 ( .C (clk), .D (signal_6519), .Q (signal_6520) ) ;
    buf_clk cell_4551 ( .C (clk), .D (signal_6521), .Q (signal_6522) ) ;
    buf_clk cell_4553 ( .C (clk), .D (signal_6523), .Q (signal_6524) ) ;
    buf_clk cell_4555 ( .C (clk), .D (signal_6525), .Q (signal_6526) ) ;
    buf_clk cell_4557 ( .C (clk), .D (signal_6527), .Q (signal_6528) ) ;
    buf_clk cell_4559 ( .C (clk), .D (signal_6529), .Q (signal_6530) ) ;
    buf_clk cell_4561 ( .C (clk), .D (signal_6531), .Q (signal_6532) ) ;
    buf_clk cell_4563 ( .C (clk), .D (signal_6533), .Q (signal_6534) ) ;
    buf_clk cell_4565 ( .C (clk), .D (signal_6535), .Q (signal_6536) ) ;
    buf_clk cell_4567 ( .C (clk), .D (signal_6537), .Q (signal_6538) ) ;
    buf_clk cell_4569 ( .C (clk), .D (signal_6539), .Q (signal_6540) ) ;
    buf_clk cell_4571 ( .C (clk), .D (signal_6541), .Q (signal_6542) ) ;
    buf_clk cell_4573 ( .C (clk), .D (signal_6543), .Q (signal_6544) ) ;
    buf_clk cell_4575 ( .C (clk), .D (signal_6545), .Q (signal_6546) ) ;
    buf_clk cell_4577 ( .C (clk), .D (signal_6547), .Q (signal_6548) ) ;
    buf_clk cell_4579 ( .C (clk), .D (signal_6549), .Q (signal_6550) ) ;
    buf_clk cell_4581 ( .C (clk), .D (signal_6551), .Q (signal_6552) ) ;
    buf_clk cell_4583 ( .C (clk), .D (signal_6553), .Q (signal_6554) ) ;
    buf_clk cell_4585 ( .C (clk), .D (signal_6555), .Q (signal_6556) ) ;
    buf_clk cell_4587 ( .C (clk), .D (signal_6557), .Q (signal_6558) ) ;
    buf_clk cell_4589 ( .C (clk), .D (signal_6559), .Q (signal_6560) ) ;
    buf_clk cell_4591 ( .C (clk), .D (signal_6561), .Q (signal_6562) ) ;
    buf_clk cell_4593 ( .C (clk), .D (signal_6563), .Q (signal_6564) ) ;
    buf_clk cell_4595 ( .C (clk), .D (signal_6565), .Q (signal_6566) ) ;
    buf_clk cell_4597 ( .C (clk), .D (signal_6567), .Q (signal_6568) ) ;
    buf_clk cell_4599 ( .C (clk), .D (signal_6569), .Q (signal_6570) ) ;
    buf_clk cell_4601 ( .C (clk), .D (signal_6571), .Q (signal_6572) ) ;
    buf_clk cell_4603 ( .C (clk), .D (signal_6573), .Q (signal_6574) ) ;
    buf_clk cell_4605 ( .C (clk), .D (signal_6575), .Q (signal_6576) ) ;
    buf_clk cell_4607 ( .C (clk), .D (signal_6577), .Q (signal_6578) ) ;
    buf_clk cell_4609 ( .C (clk), .D (signal_6579), .Q (signal_6580) ) ;
    buf_clk cell_4611 ( .C (clk), .D (signal_6581), .Q (signal_6582) ) ;
    buf_clk cell_4613 ( .C (clk), .D (signal_6583), .Q (signal_6584) ) ;
    buf_clk cell_4615 ( .C (clk), .D (signal_6585), .Q (signal_6586) ) ;
    buf_clk cell_4617 ( .C (clk), .D (signal_6587), .Q (signal_6588) ) ;
    buf_clk cell_4619 ( .C (clk), .D (signal_6589), .Q (signal_6590) ) ;
    buf_clk cell_4621 ( .C (clk), .D (signal_6591), .Q (signal_6592) ) ;
    buf_clk cell_4623 ( .C (clk), .D (signal_6593), .Q (signal_6594) ) ;
    buf_clk cell_4625 ( .C (clk), .D (signal_6595), .Q (signal_6596) ) ;
    buf_clk cell_4627 ( .C (clk), .D (signal_6597), .Q (signal_6598) ) ;
    buf_clk cell_4629 ( .C (clk), .D (signal_6599), .Q (signal_6600) ) ;
    buf_clk cell_4631 ( .C (clk), .D (signal_6601), .Q (signal_6602) ) ;
    buf_clk cell_4633 ( .C (clk), .D (signal_6603), .Q (signal_6604) ) ;
    buf_clk cell_4635 ( .C (clk), .D (signal_6605), .Q (signal_6606) ) ;
    buf_clk cell_4637 ( .C (clk), .D (signal_6607), .Q (signal_6608) ) ;
    buf_clk cell_4639 ( .C (clk), .D (signal_6609), .Q (signal_6610) ) ;
    buf_clk cell_4641 ( .C (clk), .D (signal_6611), .Q (signal_6612) ) ;
    buf_clk cell_4643 ( .C (clk), .D (signal_6613), .Q (signal_6614) ) ;
    buf_clk cell_4645 ( .C (clk), .D (signal_6615), .Q (signal_6616) ) ;
    buf_clk cell_4647 ( .C (clk), .D (signal_6617), .Q (signal_6618) ) ;
    buf_clk cell_4649 ( .C (clk), .D (signal_6619), .Q (signal_6620) ) ;
    buf_clk cell_4651 ( .C (clk), .D (signal_6621), .Q (signal_6622) ) ;
    buf_clk cell_4653 ( .C (clk), .D (signal_6623), .Q (signal_6624) ) ;
    buf_clk cell_4655 ( .C (clk), .D (signal_6625), .Q (signal_6626) ) ;
    buf_clk cell_4657 ( .C (clk), .D (signal_6627), .Q (signal_6628) ) ;
    buf_clk cell_4659 ( .C (clk), .D (signal_6629), .Q (signal_6630) ) ;
    buf_clk cell_4661 ( .C (clk), .D (signal_6631), .Q (signal_6632) ) ;
    buf_clk cell_4663 ( .C (clk), .D (signal_6633), .Q (signal_6634) ) ;
    buf_clk cell_4665 ( .C (clk), .D (signal_6635), .Q (signal_6636) ) ;
    buf_clk cell_4667 ( .C (clk), .D (signal_6637), .Q (signal_6638) ) ;
    buf_clk cell_4669 ( .C (clk), .D (signal_6639), .Q (signal_6640) ) ;
    buf_clk cell_4671 ( .C (clk), .D (signal_6641), .Q (signal_6642) ) ;
    buf_clk cell_4673 ( .C (clk), .D (signal_6643), .Q (signal_6644) ) ;
    buf_clk cell_4675 ( .C (clk), .D (signal_6645), .Q (signal_6646) ) ;
    buf_clk cell_4677 ( .C (clk), .D (signal_6647), .Q (signal_6648) ) ;
    buf_clk cell_4679 ( .C (clk), .D (signal_6649), .Q (signal_6650) ) ;
    buf_clk cell_4681 ( .C (clk), .D (signal_6651), .Q (signal_6652) ) ;
    buf_clk cell_4683 ( .C (clk), .D (signal_6653), .Q (signal_6654) ) ;
    buf_clk cell_4685 ( .C (clk), .D (signal_6655), .Q (signal_6656) ) ;
    buf_clk cell_4687 ( .C (clk), .D (signal_6657), .Q (signal_6658) ) ;
    buf_clk cell_4689 ( .C (clk), .D (signal_6659), .Q (signal_6660) ) ;
    buf_clk cell_4691 ( .C (clk), .D (signal_6661), .Q (signal_6662) ) ;
    buf_clk cell_4693 ( .C (clk), .D (signal_6663), .Q (signal_6664) ) ;
    buf_clk cell_4695 ( .C (clk), .D (signal_6665), .Q (signal_6666) ) ;
    buf_clk cell_4697 ( .C (clk), .D (signal_6667), .Q (signal_6668) ) ;
    buf_clk cell_4699 ( .C (clk), .D (signal_6669), .Q (signal_6670) ) ;
    buf_clk cell_4701 ( .C (clk), .D (signal_6671), .Q (signal_6672) ) ;
    buf_clk cell_4703 ( .C (clk), .D (signal_6673), .Q (signal_6674) ) ;
    buf_clk cell_4705 ( .C (clk), .D (signal_6675), .Q (signal_6676) ) ;
    buf_clk cell_4707 ( .C (clk), .D (signal_6677), .Q (signal_6678) ) ;
    buf_clk cell_4709 ( .C (clk), .D (signal_6679), .Q (signal_6680) ) ;
    buf_clk cell_4711 ( .C (clk), .D (signal_6681), .Q (signal_6682) ) ;
    buf_clk cell_4713 ( .C (clk), .D (signal_6683), .Q (signal_6684) ) ;
    buf_clk cell_4715 ( .C (clk), .D (signal_6685), .Q (signal_6686) ) ;
    buf_clk cell_4717 ( .C (clk), .D (signal_6687), .Q (signal_6688) ) ;
    buf_clk cell_4719 ( .C (clk), .D (signal_6689), .Q (signal_6690) ) ;
    buf_clk cell_4721 ( .C (clk), .D (signal_6691), .Q (signal_6692) ) ;
    buf_clk cell_4723 ( .C (clk), .D (signal_6693), .Q (signal_6694) ) ;
    buf_clk cell_4725 ( .C (clk), .D (signal_6695), .Q (signal_6696) ) ;
    buf_clk cell_4727 ( .C (clk), .D (signal_6697), .Q (signal_6698) ) ;
    buf_clk cell_4729 ( .C (clk), .D (signal_6699), .Q (signal_6700) ) ;
    buf_clk cell_4731 ( .C (clk), .D (signal_6701), .Q (signal_6702) ) ;
    buf_clk cell_4733 ( .C (clk), .D (signal_6703), .Q (signal_6704) ) ;
    buf_clk cell_4735 ( .C (clk), .D (signal_6705), .Q (signal_6706) ) ;
    buf_clk cell_4737 ( .C (clk), .D (signal_6707), .Q (signal_6708) ) ;
    buf_clk cell_4739 ( .C (clk), .D (signal_6709), .Q (signal_6710) ) ;
    buf_clk cell_4741 ( .C (clk), .D (signal_6711), .Q (signal_6712) ) ;
    buf_clk cell_4743 ( .C (clk), .D (signal_6713), .Q (signal_6714) ) ;
    buf_clk cell_4745 ( .C (clk), .D (signal_6715), .Q (signal_6716) ) ;
    buf_clk cell_4747 ( .C (clk), .D (signal_6717), .Q (signal_6718) ) ;
    buf_clk cell_4749 ( .C (clk), .D (signal_6719), .Q (signal_6720) ) ;
    buf_clk cell_4751 ( .C (clk), .D (signal_6721), .Q (signal_6722) ) ;
    buf_clk cell_4753 ( .C (clk), .D (signal_6723), .Q (signal_6724) ) ;
    buf_clk cell_4755 ( .C (clk), .D (signal_6725), .Q (signal_6726) ) ;
    buf_clk cell_4757 ( .C (clk), .D (signal_6727), .Q (signal_6728) ) ;
    buf_clk cell_4759 ( .C (clk), .D (signal_6729), .Q (signal_6730) ) ;
    buf_clk cell_4761 ( .C (clk), .D (signal_6731), .Q (signal_6732) ) ;
    buf_clk cell_4763 ( .C (clk), .D (signal_6733), .Q (signal_6734) ) ;
    buf_clk cell_4765 ( .C (clk), .D (signal_6735), .Q (signal_6736) ) ;
    buf_clk cell_4767 ( .C (clk), .D (signal_6737), .Q (signal_6738) ) ;
    buf_clk cell_4769 ( .C (clk), .D (signal_6739), .Q (signal_6740) ) ;
    buf_clk cell_4771 ( .C (clk), .D (signal_6741), .Q (signal_6742) ) ;
    buf_clk cell_4773 ( .C (clk), .D (signal_6743), .Q (signal_6744) ) ;
    buf_clk cell_4775 ( .C (clk), .D (signal_6745), .Q (signal_6746) ) ;
    buf_clk cell_4777 ( .C (clk), .D (signal_6747), .Q (signal_6748) ) ;
    buf_clk cell_4779 ( .C (clk), .D (signal_6749), .Q (signal_6750) ) ;
    buf_clk cell_4781 ( .C (clk), .D (signal_6751), .Q (signal_6752) ) ;
    buf_clk cell_4783 ( .C (clk), .D (signal_6753), .Q (signal_6754) ) ;
    buf_clk cell_4785 ( .C (clk), .D (signal_6755), .Q (signal_6756) ) ;
    buf_clk cell_4787 ( .C (clk), .D (signal_6757), .Q (signal_6758) ) ;
    buf_clk cell_4789 ( .C (clk), .D (signal_6759), .Q (signal_6760) ) ;
    buf_clk cell_4791 ( .C (clk), .D (signal_6761), .Q (signal_6762) ) ;
    buf_clk cell_4793 ( .C (clk), .D (signal_6763), .Q (signal_6764) ) ;
    buf_clk cell_4795 ( .C (clk), .D (signal_6765), .Q (signal_6766) ) ;
    buf_clk cell_4797 ( .C (clk), .D (signal_6767), .Q (signal_6768) ) ;
    buf_clk cell_4799 ( .C (clk), .D (signal_6769), .Q (signal_6770) ) ;
    buf_clk cell_4801 ( .C (clk), .D (signal_6771), .Q (signal_6772) ) ;
    buf_clk cell_4803 ( .C (clk), .D (signal_6773), .Q (signal_6774) ) ;
    buf_clk cell_4805 ( .C (clk), .D (signal_6775), .Q (signal_6776) ) ;
    buf_clk cell_4807 ( .C (clk), .D (signal_6777), .Q (signal_6778) ) ;
    buf_clk cell_4809 ( .C (clk), .D (signal_6779), .Q (signal_6780) ) ;
    buf_clk cell_4811 ( .C (clk), .D (signal_6781), .Q (signal_6782) ) ;
    buf_clk cell_4813 ( .C (clk), .D (signal_6783), .Q (signal_6784) ) ;
    buf_clk cell_4815 ( .C (clk), .D (signal_6785), .Q (signal_6786) ) ;
    buf_clk cell_4817 ( .C (clk), .D (signal_6787), .Q (signal_6788) ) ;
    buf_clk cell_4819 ( .C (clk), .D (signal_6789), .Q (signal_6790) ) ;
    buf_clk cell_4821 ( .C (clk), .D (signal_6791), .Q (signal_6792) ) ;
    buf_clk cell_4823 ( .C (clk), .D (signal_6793), .Q (signal_6794) ) ;
    buf_clk cell_4825 ( .C (clk), .D (signal_6795), .Q (signal_6796) ) ;
    buf_clk cell_4827 ( .C (clk), .D (signal_6797), .Q (signal_6798) ) ;
    buf_clk cell_4829 ( .C (clk), .D (signal_6799), .Q (signal_6800) ) ;
    buf_clk cell_4831 ( .C (clk), .D (signal_6801), .Q (signal_6802) ) ;
    buf_clk cell_4833 ( .C (clk), .D (signal_6803), .Q (signal_6804) ) ;
    buf_clk cell_4835 ( .C (clk), .D (signal_6805), .Q (signal_6806) ) ;
    buf_clk cell_4837 ( .C (clk), .D (signal_6807), .Q (signal_6808) ) ;
    buf_clk cell_4839 ( .C (clk), .D (signal_6809), .Q (signal_6810) ) ;
    buf_clk cell_4841 ( .C (clk), .D (signal_6811), .Q (signal_6812) ) ;
    buf_clk cell_4843 ( .C (clk), .D (signal_6813), .Q (signal_6814) ) ;
    buf_clk cell_4845 ( .C (clk), .D (signal_6815), .Q (signal_6816) ) ;
    buf_clk cell_4847 ( .C (clk), .D (signal_6817), .Q (signal_6818) ) ;
    buf_clk cell_4849 ( .C (clk), .D (signal_6819), .Q (signal_6820) ) ;
    buf_clk cell_4851 ( .C (clk), .D (signal_6821), .Q (signal_6822) ) ;
    buf_clk cell_4853 ( .C (clk), .D (signal_6823), .Q (signal_6824) ) ;
    buf_clk cell_4855 ( .C (clk), .D (signal_6825), .Q (signal_6826) ) ;
    buf_clk cell_4857 ( .C (clk), .D (signal_6827), .Q (signal_6828) ) ;
    buf_clk cell_4859 ( .C (clk), .D (signal_6829), .Q (signal_6830) ) ;
    buf_clk cell_4861 ( .C (clk), .D (signal_6831), .Q (signal_6832) ) ;
    buf_clk cell_4863 ( .C (clk), .D (signal_6833), .Q (signal_6834) ) ;
    buf_clk cell_4865 ( .C (clk), .D (signal_6835), .Q (signal_6836) ) ;
    buf_clk cell_4867 ( .C (clk), .D (signal_6837), .Q (signal_6838) ) ;
    buf_clk cell_4869 ( .C (clk), .D (signal_6839), .Q (signal_6840) ) ;
    buf_clk cell_4871 ( .C (clk), .D (signal_6841), .Q (signal_6842) ) ;
    buf_clk cell_4873 ( .C (clk), .D (signal_6843), .Q (signal_6844) ) ;
    buf_clk cell_4875 ( .C (clk), .D (signal_6845), .Q (signal_6846) ) ;
    buf_clk cell_4877 ( .C (clk), .D (signal_6847), .Q (signal_6848) ) ;
    buf_clk cell_4879 ( .C (clk), .D (signal_6849), .Q (signal_6850) ) ;
    buf_clk cell_4881 ( .C (clk), .D (signal_6851), .Q (signal_6852) ) ;
    buf_clk cell_4883 ( .C (clk), .D (signal_6853), .Q (signal_6854) ) ;
    buf_clk cell_4885 ( .C (clk), .D (signal_6855), .Q (signal_6856) ) ;
    buf_clk cell_4887 ( .C (clk), .D (signal_6857), .Q (signal_6858) ) ;
    buf_clk cell_4889 ( .C (clk), .D (signal_6859), .Q (signal_6860) ) ;
    buf_clk cell_4891 ( .C (clk), .D (signal_6861), .Q (signal_6862) ) ;
    buf_clk cell_4893 ( .C (clk), .D (signal_6863), .Q (signal_6864) ) ;
    buf_clk cell_4895 ( .C (clk), .D (signal_6865), .Q (signal_6866) ) ;
    buf_clk cell_4897 ( .C (clk), .D (signal_6867), .Q (signal_6868) ) ;
    buf_clk cell_4899 ( .C (clk), .D (signal_6869), .Q (signal_6870) ) ;
    buf_clk cell_4901 ( .C (clk), .D (signal_6871), .Q (signal_6872) ) ;
    buf_clk cell_4903 ( .C (clk), .D (signal_6873), .Q (signal_6874) ) ;
    buf_clk cell_4905 ( .C (clk), .D (signal_6875), .Q (signal_6876) ) ;
    buf_clk cell_4907 ( .C (clk), .D (signal_6877), .Q (signal_6878) ) ;
    buf_clk cell_4909 ( .C (clk), .D (signal_6879), .Q (signal_6880) ) ;
    buf_clk cell_4911 ( .C (clk), .D (signal_6881), .Q (signal_6882) ) ;
    buf_clk cell_4913 ( .C (clk), .D (signal_6883), .Q (signal_6884) ) ;
    buf_clk cell_4915 ( .C (clk), .D (signal_6885), .Q (signal_6886) ) ;
    buf_clk cell_4917 ( .C (clk), .D (signal_6887), .Q (signal_6888) ) ;
    buf_clk cell_4919 ( .C (clk), .D (signal_6889), .Q (signal_6890) ) ;
    buf_clk cell_4921 ( .C (clk), .D (signal_6891), .Q (signal_6892) ) ;
    buf_clk cell_4923 ( .C (clk), .D (signal_6893), .Q (signal_6894) ) ;
    buf_clk cell_4925 ( .C (clk), .D (signal_6895), .Q (signal_6896) ) ;
    buf_clk cell_4927 ( .C (clk), .D (signal_6897), .Q (signal_6898) ) ;
    buf_clk cell_4929 ( .C (clk), .D (signal_6899), .Q (signal_6900) ) ;
    buf_clk cell_4931 ( .C (clk), .D (signal_6901), .Q (signal_6902) ) ;
    buf_clk cell_4933 ( .C (clk), .D (signal_6903), .Q (signal_6904) ) ;
    buf_clk cell_4935 ( .C (clk), .D (signal_6905), .Q (signal_6906) ) ;
    buf_clk cell_4937 ( .C (clk), .D (signal_6907), .Q (signal_6908) ) ;
    buf_clk cell_4939 ( .C (clk), .D (signal_6909), .Q (signal_6910) ) ;
    buf_clk cell_4941 ( .C (clk), .D (signal_6911), .Q (signal_6912) ) ;
    buf_clk cell_4943 ( .C (clk), .D (signal_6913), .Q (signal_6914) ) ;
    buf_clk cell_4945 ( .C (clk), .D (signal_6915), .Q (signal_6916) ) ;
    buf_clk cell_4947 ( .C (clk), .D (signal_6917), .Q (signal_6918) ) ;
    buf_clk cell_4949 ( .C (clk), .D (signal_6919), .Q (signal_6920) ) ;
    buf_clk cell_4951 ( .C (clk), .D (signal_6921), .Q (signal_6922) ) ;
    buf_clk cell_4953 ( .C (clk), .D (signal_6923), .Q (signal_6924) ) ;
    buf_clk cell_4955 ( .C (clk), .D (signal_6925), .Q (signal_6926) ) ;
    buf_clk cell_4957 ( .C (clk), .D (signal_6927), .Q (signal_6928) ) ;
    buf_clk cell_4959 ( .C (clk), .D (signal_6929), .Q (signal_6930) ) ;
    buf_clk cell_4961 ( .C (clk), .D (signal_6931), .Q (signal_6932) ) ;
    buf_clk cell_4963 ( .C (clk), .D (signal_6933), .Q (signal_6934) ) ;
    buf_clk cell_4965 ( .C (clk), .D (signal_6935), .Q (signal_6936) ) ;
    buf_clk cell_4967 ( .C (clk), .D (signal_6937), .Q (signal_6938) ) ;
    buf_clk cell_4969 ( .C (clk), .D (signal_6939), .Q (signal_6940) ) ;
    buf_clk cell_4971 ( .C (clk), .D (signal_6941), .Q (signal_6942) ) ;
    buf_clk cell_4973 ( .C (clk), .D (signal_6943), .Q (signal_6944) ) ;
    buf_clk cell_4975 ( .C (clk), .D (signal_6945), .Q (signal_6946) ) ;
    buf_clk cell_4977 ( .C (clk), .D (signal_6947), .Q (signal_6948) ) ;
    buf_clk cell_4979 ( .C (clk), .D (signal_6949), .Q (signal_6950) ) ;
    buf_clk cell_4981 ( .C (clk), .D (signal_6951), .Q (signal_6952) ) ;
    buf_clk cell_4983 ( .C (clk), .D (signal_6953), .Q (signal_6954) ) ;
    buf_clk cell_4985 ( .C (clk), .D (signal_6955), .Q (signal_6956) ) ;
    buf_clk cell_4987 ( .C (clk), .D (signal_6957), .Q (signal_6958) ) ;
    buf_clk cell_4989 ( .C (clk), .D (signal_6959), .Q (signal_6960) ) ;
    buf_clk cell_4991 ( .C (clk), .D (signal_6961), .Q (signal_6962) ) ;
    buf_clk cell_4993 ( .C (clk), .D (signal_6963), .Q (signal_6964) ) ;
    buf_clk cell_4995 ( .C (clk), .D (signal_6965), .Q (signal_6966) ) ;
    buf_clk cell_4997 ( .C (clk), .D (signal_6967), .Q (signal_6968) ) ;
    buf_clk cell_4999 ( .C (clk), .D (signal_6969), .Q (signal_6970) ) ;
    buf_clk cell_5001 ( .C (clk), .D (signal_6971), .Q (signal_6972) ) ;
    buf_clk cell_5003 ( .C (clk), .D (signal_6973), .Q (signal_6974) ) ;
    buf_clk cell_5005 ( .C (clk), .D (signal_6975), .Q (signal_6976) ) ;
    buf_clk cell_5007 ( .C (clk), .D (signal_6977), .Q (signal_6978) ) ;
    buf_clk cell_5009 ( .C (clk), .D (signal_6979), .Q (signal_6980) ) ;
    buf_clk cell_5011 ( .C (clk), .D (signal_6981), .Q (signal_6982) ) ;
    buf_clk cell_5013 ( .C (clk), .D (signal_6983), .Q (signal_6984) ) ;
    buf_clk cell_5015 ( .C (clk), .D (signal_6985), .Q (signal_6986) ) ;
    buf_clk cell_5017 ( .C (clk), .D (signal_6987), .Q (signal_6988) ) ;
    buf_clk cell_5019 ( .C (clk), .D (signal_6989), .Q (signal_6990) ) ;
    buf_clk cell_5021 ( .C (clk), .D (signal_6991), .Q (signal_6992) ) ;
    buf_clk cell_5023 ( .C (clk), .D (signal_6993), .Q (signal_6994) ) ;
    buf_clk cell_5025 ( .C (clk), .D (signal_6995), .Q (signal_6996) ) ;
    buf_clk cell_5027 ( .C (clk), .D (signal_6997), .Q (signal_6998) ) ;
    buf_clk cell_5029 ( .C (clk), .D (signal_6999), .Q (signal_7000) ) ;
    buf_clk cell_5031 ( .C (clk), .D (signal_7001), .Q (signal_7002) ) ;
    buf_clk cell_5033 ( .C (clk), .D (signal_7003), .Q (signal_7004) ) ;
    buf_clk cell_5035 ( .C (clk), .D (signal_7005), .Q (signal_7006) ) ;
    buf_clk cell_5037 ( .C (clk), .D (signal_7007), .Q (signal_7008) ) ;
    buf_clk cell_5039 ( .C (clk), .D (signal_7009), .Q (signal_7010) ) ;
    buf_clk cell_5041 ( .C (clk), .D (signal_7011), .Q (signal_7012) ) ;
    buf_clk cell_5043 ( .C (clk), .D (signal_7013), .Q (signal_7014) ) ;
    buf_clk cell_5045 ( .C (clk), .D (signal_7015), .Q (signal_7016) ) ;
    buf_clk cell_5047 ( .C (clk), .D (signal_7017), .Q (signal_7018) ) ;
    buf_clk cell_5049 ( .C (clk), .D (signal_7019), .Q (signal_7020) ) ;
    buf_clk cell_5051 ( .C (clk), .D (signal_7021), .Q (signal_7022) ) ;
    buf_clk cell_5053 ( .C (clk), .D (signal_7023), .Q (signal_7024) ) ;
    buf_clk cell_5055 ( .C (clk), .D (signal_7025), .Q (signal_7026) ) ;
    buf_clk cell_5057 ( .C (clk), .D (signal_7027), .Q (signal_7028) ) ;
    buf_clk cell_5059 ( .C (clk), .D (signal_7029), .Q (signal_7030) ) ;
    buf_clk cell_5061 ( .C (clk), .D (signal_7031), .Q (signal_7032) ) ;
    buf_clk cell_5063 ( .C (clk), .D (signal_7033), .Q (signal_7034) ) ;
    buf_clk cell_5065 ( .C (clk), .D (signal_7035), .Q (signal_7036) ) ;
    buf_clk cell_5067 ( .C (clk), .D (signal_7037), .Q (signal_7038) ) ;
    buf_clk cell_5069 ( .C (clk), .D (signal_7039), .Q (signal_7040) ) ;
    buf_clk cell_5071 ( .C (clk), .D (signal_7041), .Q (signal_7042) ) ;
    buf_clk cell_5073 ( .C (clk), .D (signal_7043), .Q (signal_7044) ) ;
    buf_clk cell_5075 ( .C (clk), .D (signal_7045), .Q (signal_7046) ) ;
    buf_clk cell_5077 ( .C (clk), .D (signal_7047), .Q (signal_7048) ) ;
    buf_clk cell_5079 ( .C (clk), .D (signal_7049), .Q (signal_7050) ) ;
    buf_clk cell_5081 ( .C (clk), .D (signal_7051), .Q (signal_7052) ) ;
    buf_clk cell_5083 ( .C (clk), .D (signal_7053), .Q (signal_7054) ) ;
    buf_clk cell_5085 ( .C (clk), .D (signal_7055), .Q (signal_7056) ) ;
    buf_clk cell_5087 ( .C (clk), .D (signal_7057), .Q (signal_7058) ) ;
    buf_clk cell_5089 ( .C (clk), .D (signal_7059), .Q (signal_7060) ) ;
    buf_clk cell_5091 ( .C (clk), .D (signal_7061), .Q (signal_7062) ) ;
    buf_clk cell_5093 ( .C (clk), .D (signal_7063), .Q (signal_7064) ) ;
    buf_clk cell_5095 ( .C (clk), .D (signal_7065), .Q (signal_7066) ) ;
    buf_clk cell_5097 ( .C (clk), .D (signal_7067), .Q (signal_7068) ) ;
    buf_clk cell_5099 ( .C (clk), .D (signal_7069), .Q (signal_7070) ) ;
    buf_clk cell_5101 ( .C (clk), .D (signal_7071), .Q (signal_7072) ) ;
    buf_clk cell_5103 ( .C (clk), .D (signal_7073), .Q (signal_7074) ) ;
    buf_clk cell_5105 ( .C (clk), .D (signal_7075), .Q (signal_7076) ) ;
    buf_clk cell_5107 ( .C (clk), .D (signal_7077), .Q (signal_7078) ) ;
    buf_clk cell_5109 ( .C (clk), .D (signal_7079), .Q (signal_7080) ) ;
    buf_clk cell_5111 ( .C (clk), .D (signal_7081), .Q (signal_7082) ) ;
    buf_clk cell_5113 ( .C (clk), .D (signal_7083), .Q (signal_7084) ) ;
    buf_clk cell_5115 ( .C (clk), .D (signal_7085), .Q (signal_7086) ) ;
    buf_clk cell_5117 ( .C (clk), .D (signal_7087), .Q (signal_7088) ) ;
    buf_clk cell_5119 ( .C (clk), .D (signal_7089), .Q (signal_7090) ) ;
    buf_clk cell_5121 ( .C (clk), .D (signal_7091), .Q (signal_7092) ) ;
    buf_clk cell_5123 ( .C (clk), .D (signal_7093), .Q (signal_7094) ) ;
    buf_clk cell_5125 ( .C (clk), .D (signal_7095), .Q (signal_7096) ) ;
    buf_clk cell_5127 ( .C (clk), .D (signal_7097), .Q (signal_7098) ) ;
    buf_clk cell_5129 ( .C (clk), .D (signal_7099), .Q (signal_7100) ) ;
    buf_clk cell_5131 ( .C (clk), .D (signal_7101), .Q (signal_7102) ) ;
    buf_clk cell_5133 ( .C (clk), .D (signal_7103), .Q (signal_7104) ) ;
    buf_clk cell_5135 ( .C (clk), .D (signal_7105), .Q (signal_7106) ) ;
    buf_clk cell_5137 ( .C (clk), .D (signal_7107), .Q (signal_7108) ) ;
    buf_clk cell_5139 ( .C (clk), .D (signal_7109), .Q (signal_7110) ) ;
    buf_clk cell_5141 ( .C (clk), .D (signal_7111), .Q (signal_7112) ) ;
    buf_clk cell_5143 ( .C (clk), .D (signal_7113), .Q (signal_7114) ) ;
    buf_clk cell_5145 ( .C (clk), .D (signal_7115), .Q (signal_7116) ) ;
    buf_clk cell_5147 ( .C (clk), .D (signal_7117), .Q (signal_7118) ) ;
    buf_clk cell_5149 ( .C (clk), .D (signal_7119), .Q (signal_7120) ) ;
    buf_clk cell_5151 ( .C (clk), .D (signal_7121), .Q (signal_7122) ) ;
    buf_clk cell_5153 ( .C (clk), .D (signal_7123), .Q (signal_7124) ) ;
    buf_clk cell_5155 ( .C (clk), .D (signal_7125), .Q (signal_7126) ) ;
    buf_clk cell_5157 ( .C (clk), .D (signal_7127), .Q (signal_7128) ) ;
    buf_clk cell_5159 ( .C (clk), .D (signal_7129), .Q (signal_7130) ) ;
    buf_clk cell_5161 ( .C (clk), .D (signal_7131), .Q (signal_7132) ) ;
    buf_clk cell_5163 ( .C (clk), .D (signal_7133), .Q (signal_7134) ) ;
    buf_clk cell_5165 ( .C (clk), .D (signal_7135), .Q (signal_7136) ) ;
    buf_clk cell_5167 ( .C (clk), .D (signal_7137), .Q (signal_7138) ) ;
    buf_clk cell_5169 ( .C (clk), .D (signal_7139), .Q (signal_7140) ) ;
    buf_clk cell_5171 ( .C (clk), .D (signal_7141), .Q (signal_7142) ) ;
    buf_clk cell_5173 ( .C (clk), .D (signal_7143), .Q (signal_7144) ) ;
    buf_clk cell_5175 ( .C (clk), .D (signal_7145), .Q (signal_7146) ) ;
    buf_clk cell_5177 ( .C (clk), .D (signal_7147), .Q (signal_7148) ) ;
    buf_clk cell_5179 ( .C (clk), .D (signal_7149), .Q (signal_7150) ) ;
    buf_clk cell_5181 ( .C (clk), .D (signal_7151), .Q (signal_7152) ) ;
    buf_clk cell_5183 ( .C (clk), .D (signal_7153), .Q (signal_7154) ) ;
    buf_clk cell_5185 ( .C (clk), .D (signal_7155), .Q (signal_7156) ) ;
    buf_clk cell_5187 ( .C (clk), .D (signal_7157), .Q (signal_7158) ) ;
    buf_clk cell_5189 ( .C (clk), .D (signal_7159), .Q (signal_7160) ) ;
    buf_clk cell_5191 ( .C (clk), .D (signal_7161), .Q (signal_7162) ) ;
    buf_clk cell_5193 ( .C (clk), .D (signal_7163), .Q (signal_7164) ) ;
    buf_clk cell_5195 ( .C (clk), .D (signal_7165), .Q (signal_7166) ) ;
    buf_clk cell_5197 ( .C (clk), .D (signal_7167), .Q (signal_7168) ) ;
    buf_clk cell_5199 ( .C (clk), .D (signal_7169), .Q (signal_7170) ) ;
    buf_clk cell_5201 ( .C (clk), .D (signal_7171), .Q (signal_7172) ) ;
    buf_clk cell_5203 ( .C (clk), .D (signal_7173), .Q (signal_7174) ) ;
    buf_clk cell_5205 ( .C (clk), .D (signal_7175), .Q (signal_7176) ) ;
    buf_clk cell_5207 ( .C (clk), .D (signal_7177), .Q (signal_7178) ) ;
    buf_clk cell_5209 ( .C (clk), .D (signal_7179), .Q (signal_7180) ) ;
    buf_clk cell_5211 ( .C (clk), .D (signal_7181), .Q (signal_7182) ) ;
    buf_clk cell_5213 ( .C (clk), .D (signal_7183), .Q (signal_7184) ) ;
    buf_clk cell_5215 ( .C (clk), .D (signal_7185), .Q (signal_7186) ) ;
    buf_clk cell_5217 ( .C (clk), .D (signal_7187), .Q (signal_7188) ) ;
    buf_clk cell_5219 ( .C (clk), .D (signal_7189), .Q (signal_7190) ) ;
    buf_clk cell_5221 ( .C (clk), .D (signal_7191), .Q (signal_7192) ) ;
    buf_clk cell_5223 ( .C (clk), .D (signal_7193), .Q (signal_7194) ) ;
    buf_clk cell_5225 ( .C (clk), .D (signal_7195), .Q (signal_7196) ) ;
    buf_clk cell_5227 ( .C (clk), .D (signal_7197), .Q (signal_7198) ) ;
    buf_clk cell_5229 ( .C (clk), .D (signal_7199), .Q (signal_7200) ) ;
    buf_clk cell_5231 ( .C (clk), .D (signal_7201), .Q (signal_7202) ) ;
    buf_clk cell_5233 ( .C (clk), .D (signal_7203), .Q (signal_7204) ) ;
    buf_clk cell_5235 ( .C (clk), .D (signal_7205), .Q (signal_7206) ) ;
    buf_clk cell_5237 ( .C (clk), .D (signal_7207), .Q (signal_7208) ) ;
    buf_clk cell_5239 ( .C (clk), .D (signal_7209), .Q (signal_7210) ) ;
    buf_clk cell_5241 ( .C (clk), .D (signal_7211), .Q (signal_7212) ) ;
    buf_clk cell_5243 ( .C (clk), .D (signal_7213), .Q (signal_7214) ) ;
    buf_clk cell_5245 ( .C (clk), .D (signal_7215), .Q (signal_7216) ) ;
    buf_clk cell_5247 ( .C (clk), .D (signal_7217), .Q (signal_7218) ) ;
    buf_clk cell_5249 ( .C (clk), .D (signal_7219), .Q (signal_7220) ) ;
    buf_clk cell_5251 ( .C (clk), .D (signal_7221), .Q (signal_7222) ) ;
    buf_clk cell_5253 ( .C (clk), .D (signal_7223), .Q (signal_7224) ) ;
    buf_clk cell_5255 ( .C (clk), .D (signal_7225), .Q (signal_7226) ) ;
    buf_clk cell_5257 ( .C (clk), .D (signal_7227), .Q (signal_7228) ) ;
    buf_clk cell_5259 ( .C (clk), .D (signal_7229), .Q (signal_7230) ) ;
    buf_clk cell_5261 ( .C (clk), .D (signal_7231), .Q (signal_7232) ) ;
    buf_clk cell_5263 ( .C (clk), .D (signal_7233), .Q (signal_7234) ) ;
    buf_clk cell_5265 ( .C (clk), .D (signal_7235), .Q (signal_7236) ) ;
    buf_clk cell_5267 ( .C (clk), .D (signal_7237), .Q (signal_7238) ) ;
    buf_clk cell_5269 ( .C (clk), .D (signal_7239), .Q (signal_7240) ) ;
    buf_clk cell_5271 ( .C (clk), .D (signal_7241), .Q (signal_7242) ) ;
    buf_clk cell_5273 ( .C (clk), .D (signal_7243), .Q (signal_7244) ) ;
    buf_clk cell_5275 ( .C (clk), .D (signal_7245), .Q (signal_7246) ) ;
    buf_clk cell_5277 ( .C (clk), .D (signal_7247), .Q (signal_7248) ) ;
    buf_clk cell_5279 ( .C (clk), .D (signal_7249), .Q (signal_7250) ) ;
    buf_clk cell_5281 ( .C (clk), .D (signal_7251), .Q (signal_7252) ) ;
    buf_clk cell_5283 ( .C (clk), .D (signal_7253), .Q (signal_7254) ) ;
    buf_clk cell_5285 ( .C (clk), .D (signal_7255), .Q (signal_7256) ) ;
    buf_clk cell_5287 ( .C (clk), .D (signal_7257), .Q (signal_7258) ) ;
    buf_clk cell_5289 ( .C (clk), .D (signal_7259), .Q (signal_7260) ) ;
    buf_clk cell_5291 ( .C (clk), .D (signal_7261), .Q (signal_7262) ) ;
    buf_clk cell_5293 ( .C (clk), .D (signal_7263), .Q (signal_7264) ) ;
    buf_clk cell_5295 ( .C (clk), .D (signal_7265), .Q (signal_7266) ) ;
    buf_clk cell_5297 ( .C (clk), .D (signal_7267), .Q (signal_7268) ) ;
    buf_clk cell_5299 ( .C (clk), .D (signal_7269), .Q (signal_7270) ) ;
    buf_clk cell_5301 ( .C (clk), .D (signal_7271), .Q (signal_7272) ) ;
    buf_clk cell_5303 ( .C (clk), .D (signal_7273), .Q (signal_7274) ) ;
    buf_clk cell_5305 ( .C (clk), .D (signal_7275), .Q (signal_7276) ) ;
    buf_clk cell_5307 ( .C (clk), .D (signal_7277), .Q (signal_7278) ) ;
    buf_clk cell_5309 ( .C (clk), .D (signal_7279), .Q (signal_7280) ) ;
    buf_clk cell_5311 ( .C (clk), .D (signal_7281), .Q (signal_7282) ) ;
    buf_clk cell_5313 ( .C (clk), .D (signal_7283), .Q (signal_7284) ) ;
    buf_clk cell_5315 ( .C (clk), .D (signal_7285), .Q (signal_7286) ) ;
    buf_clk cell_5317 ( .C (clk), .D (signal_7287), .Q (signal_7288) ) ;
    buf_clk cell_5319 ( .C (clk), .D (signal_7289), .Q (signal_7290) ) ;
    buf_clk cell_5321 ( .C (clk), .D (signal_7291), .Q (signal_7292) ) ;
    buf_clk cell_5323 ( .C (clk), .D (signal_7293), .Q (signal_7294) ) ;
    buf_clk cell_5325 ( .C (clk), .D (signal_7295), .Q (signal_7296) ) ;
    buf_clk cell_5327 ( .C (clk), .D (signal_7297), .Q (signal_7298) ) ;
    buf_clk cell_5329 ( .C (clk), .D (signal_7299), .Q (signal_7300) ) ;
    buf_clk cell_5331 ( .C (clk), .D (signal_7301), .Q (signal_7302) ) ;
    buf_clk cell_5333 ( .C (clk), .D (signal_7303), .Q (signal_7304) ) ;
    buf_clk cell_5335 ( .C (clk), .D (signal_7305), .Q (signal_7306) ) ;
    buf_clk cell_5337 ( .C (clk), .D (signal_7307), .Q (signal_7308) ) ;
    buf_clk cell_5339 ( .C (clk), .D (signal_7309), .Q (signal_7310) ) ;
    buf_clk cell_5341 ( .C (clk), .D (signal_7311), .Q (signal_7312) ) ;
    buf_clk cell_5343 ( .C (clk), .D (signal_7313), .Q (signal_7314) ) ;
    buf_clk cell_5345 ( .C (clk), .D (signal_7315), .Q (signal_7316) ) ;
    buf_clk cell_5347 ( .C (clk), .D (signal_7317), .Q (signal_7318) ) ;
    buf_clk cell_5349 ( .C (clk), .D (signal_7319), .Q (signal_7320) ) ;
    buf_clk cell_5351 ( .C (clk), .D (signal_7321), .Q (signal_7322) ) ;
    buf_clk cell_5353 ( .C (clk), .D (signal_7323), .Q (signal_7324) ) ;
    buf_clk cell_5355 ( .C (clk), .D (signal_7325), .Q (signal_7326) ) ;
    buf_clk cell_5357 ( .C (clk), .D (signal_7327), .Q (signal_7328) ) ;
    buf_clk cell_5359 ( .C (clk), .D (signal_7329), .Q (signal_7330) ) ;
    buf_clk cell_5361 ( .C (clk), .D (signal_7331), .Q (signal_7332) ) ;
    buf_clk cell_5363 ( .C (clk), .D (signal_7333), .Q (signal_7334) ) ;
    buf_clk cell_5365 ( .C (clk), .D (signal_7335), .Q (signal_7336) ) ;
    buf_clk cell_5367 ( .C (clk), .D (signal_7337), .Q (signal_7338) ) ;
    buf_clk cell_5369 ( .C (clk), .D (signal_7339), .Q (signal_7340) ) ;
    buf_clk cell_5371 ( .C (clk), .D (signal_7341), .Q (signal_7342) ) ;
    buf_clk cell_5373 ( .C (clk), .D (signal_7343), .Q (signal_7344) ) ;
    buf_clk cell_5375 ( .C (clk), .D (signal_7345), .Q (signal_7346) ) ;
    buf_clk cell_5377 ( .C (clk), .D (signal_7347), .Q (signal_7348) ) ;
    buf_clk cell_5379 ( .C (clk), .D (signal_7349), .Q (signal_7350) ) ;
    buf_clk cell_5381 ( .C (clk), .D (signal_7351), .Q (signal_7352) ) ;
    buf_clk cell_5383 ( .C (clk), .D (signal_7353), .Q (signal_7354) ) ;
    buf_clk cell_5385 ( .C (clk), .D (signal_7355), .Q (signal_7356) ) ;
    buf_clk cell_5387 ( .C (clk), .D (signal_7357), .Q (signal_7358) ) ;
    buf_clk cell_5389 ( .C (clk), .D (signal_7359), .Q (signal_7360) ) ;
    buf_clk cell_5391 ( .C (clk), .D (signal_7361), .Q (signal_7362) ) ;
    buf_clk cell_5393 ( .C (clk), .D (signal_7363), .Q (signal_7364) ) ;
    buf_clk cell_5395 ( .C (clk), .D (signal_7365), .Q (signal_7366) ) ;
    buf_clk cell_5397 ( .C (clk), .D (signal_7367), .Q (signal_7368) ) ;
    buf_clk cell_5399 ( .C (clk), .D (signal_7369), .Q (signal_7370) ) ;
    buf_clk cell_5401 ( .C (clk), .D (signal_7371), .Q (signal_7372) ) ;
    buf_clk cell_5403 ( .C (clk), .D (signal_7373), .Q (signal_7374) ) ;
    buf_clk cell_5405 ( .C (clk), .D (signal_7375), .Q (signal_7376) ) ;
    buf_clk cell_5407 ( .C (clk), .D (signal_7377), .Q (signal_7378) ) ;
    buf_clk cell_5409 ( .C (clk), .D (signal_7379), .Q (signal_7380) ) ;
    buf_clk cell_5411 ( .C (clk), .D (signal_7381), .Q (signal_7382) ) ;
    buf_clk cell_5413 ( .C (clk), .D (signal_7383), .Q (signal_7384) ) ;
    buf_clk cell_5415 ( .C (clk), .D (signal_7385), .Q (signal_7386) ) ;
    buf_clk cell_5417 ( .C (clk), .D (signal_7387), .Q (signal_7388) ) ;
    buf_clk cell_5419 ( .C (clk), .D (signal_7389), .Q (signal_7390) ) ;
    buf_clk cell_5421 ( .C (clk), .D (signal_7391), .Q (signal_7392) ) ;
    buf_clk cell_5423 ( .C (clk), .D (signal_7393), .Q (signal_7394) ) ;
    buf_clk cell_5425 ( .C (clk), .D (signal_7395), .Q (signal_7396) ) ;
    buf_clk cell_5427 ( .C (clk), .D (signal_7397), .Q (signal_7398) ) ;
    buf_clk cell_5429 ( .C (clk), .D (signal_7399), .Q (signal_7400) ) ;
    buf_clk cell_5431 ( .C (clk), .D (signal_7401), .Q (signal_7402) ) ;
    buf_clk cell_5433 ( .C (clk), .D (signal_7403), .Q (signal_7404) ) ;
    buf_clk cell_5435 ( .C (clk), .D (signal_7405), .Q (signal_7406) ) ;
    buf_clk cell_5437 ( .C (clk), .D (signal_7407), .Q (signal_7408) ) ;
    buf_clk cell_5439 ( .C (clk), .D (signal_7409), .Q (signal_7410) ) ;
    buf_clk cell_5441 ( .C (clk), .D (signal_7411), .Q (signal_7412) ) ;
    buf_clk cell_5443 ( .C (clk), .D (signal_7413), .Q (signal_7414) ) ;
    buf_clk cell_5445 ( .C (clk), .D (signal_7415), .Q (signal_7416) ) ;
    buf_clk cell_5447 ( .C (clk), .D (signal_7417), .Q (signal_7418) ) ;
    buf_clk cell_5449 ( .C (clk), .D (signal_7419), .Q (signal_7420) ) ;
    buf_clk cell_5451 ( .C (clk), .D (signal_7421), .Q (signal_7422) ) ;
    buf_clk cell_5453 ( .C (clk), .D (signal_7423), .Q (signal_7424) ) ;
    buf_clk cell_5455 ( .C (clk), .D (signal_7425), .Q (signal_7426) ) ;
    buf_clk cell_5457 ( .C (clk), .D (signal_7427), .Q (signal_7428) ) ;
    buf_clk cell_5459 ( .C (clk), .D (signal_7429), .Q (signal_7430) ) ;
    buf_clk cell_5461 ( .C (clk), .D (signal_7431), .Q (signal_7432) ) ;
    buf_clk cell_5463 ( .C (clk), .D (signal_7433), .Q (signal_7434) ) ;
    buf_clk cell_5465 ( .C (clk), .D (signal_7435), .Q (signal_7436) ) ;
    buf_clk cell_5467 ( .C (clk), .D (signal_7437), .Q (signal_7438) ) ;
    buf_clk cell_5469 ( .C (clk), .D (signal_7439), .Q (signal_7440) ) ;
    buf_clk cell_5471 ( .C (clk), .D (signal_7441), .Q (signal_7442) ) ;
    buf_clk cell_5473 ( .C (clk), .D (signal_7443), .Q (signal_7444) ) ;
    buf_clk cell_5475 ( .C (clk), .D (signal_7445), .Q (signal_7446) ) ;
    buf_clk cell_5477 ( .C (clk), .D (signal_7447), .Q (signal_7448) ) ;
    buf_clk cell_5479 ( .C (clk), .D (signal_7449), .Q (signal_7450) ) ;
    buf_clk cell_5481 ( .C (clk), .D (signal_7451), .Q (signal_7452) ) ;
    buf_clk cell_5483 ( .C (clk), .D (signal_7453), .Q (signal_7454) ) ;
    buf_clk cell_5485 ( .C (clk), .D (signal_7455), .Q (signal_7456) ) ;
    buf_clk cell_5487 ( .C (clk), .D (signal_7457), .Q (signal_7458) ) ;
    buf_clk cell_5489 ( .C (clk), .D (signal_7459), .Q (signal_7460) ) ;
    buf_clk cell_5491 ( .C (clk), .D (signal_7461), .Q (signal_7462) ) ;
    buf_clk cell_5493 ( .C (clk), .D (signal_7463), .Q (signal_7464) ) ;
    buf_clk cell_5495 ( .C (clk), .D (signal_7465), .Q (signal_7466) ) ;
    buf_clk cell_5497 ( .C (clk), .D (signal_7467), .Q (signal_7468) ) ;
    buf_clk cell_5499 ( .C (clk), .D (signal_7469), .Q (signal_7470) ) ;
    buf_clk cell_5501 ( .C (clk), .D (signal_7471), .Q (signal_7472) ) ;
    buf_clk cell_5503 ( .C (clk), .D (signal_7473), .Q (signal_7474) ) ;
    buf_clk cell_5505 ( .C (clk), .D (signal_7475), .Q (signal_7476) ) ;
    buf_clk cell_5507 ( .C (clk), .D (signal_7477), .Q (signal_7478) ) ;
    buf_clk cell_5509 ( .C (clk), .D (signal_7479), .Q (signal_7480) ) ;
    buf_clk cell_5511 ( .C (clk), .D (signal_7481), .Q (signal_7482) ) ;
    buf_clk cell_5513 ( .C (clk), .D (signal_7483), .Q (signal_7484) ) ;
    buf_clk cell_5515 ( .C (clk), .D (signal_7485), .Q (signal_7486) ) ;
    buf_clk cell_5517 ( .C (clk), .D (signal_7487), .Q (signal_7488) ) ;
    buf_clk cell_5519 ( .C (clk), .D (signal_7489), .Q (signal_7490) ) ;
    buf_clk cell_5521 ( .C (clk), .D (signal_7491), .Q (signal_7492) ) ;
    buf_clk cell_5523 ( .C (clk), .D (signal_7493), .Q (signal_7494) ) ;
    buf_clk cell_5525 ( .C (clk), .D (signal_7495), .Q (signal_7496) ) ;
    buf_clk cell_5527 ( .C (clk), .D (signal_7497), .Q (signal_7498) ) ;
    buf_clk cell_5529 ( .C (clk), .D (signal_7499), .Q (signal_7500) ) ;
    buf_clk cell_5531 ( .C (clk), .D (signal_7501), .Q (signal_7502) ) ;
    buf_clk cell_5533 ( .C (clk), .D (signal_7503), .Q (signal_7504) ) ;
    buf_clk cell_5535 ( .C (clk), .D (signal_7505), .Q (signal_7506) ) ;
    buf_clk cell_5537 ( .C (clk), .D (signal_7507), .Q (signal_7508) ) ;
    buf_clk cell_5539 ( .C (clk), .D (signal_7509), .Q (signal_7510) ) ;
    buf_clk cell_5541 ( .C (clk), .D (signal_7511), .Q (signal_7512) ) ;
    buf_clk cell_5543 ( .C (clk), .D (signal_7513), .Q (signal_7514) ) ;
    buf_clk cell_5545 ( .C (clk), .D (signal_7515), .Q (signal_7516) ) ;
    buf_clk cell_5547 ( .C (clk), .D (signal_7517), .Q (signal_7518) ) ;
    buf_clk cell_5549 ( .C (clk), .D (signal_7519), .Q (signal_7520) ) ;
    buf_clk cell_5551 ( .C (clk), .D (signal_7521), .Q (signal_7522) ) ;
    buf_clk cell_5553 ( .C (clk), .D (signal_7523), .Q (signal_7524) ) ;
    buf_clk cell_5555 ( .C (clk), .D (signal_7525), .Q (signal_7526) ) ;
    buf_clk cell_5557 ( .C (clk), .D (signal_7527), .Q (signal_7528) ) ;
    buf_clk cell_5559 ( .C (clk), .D (signal_7529), .Q (signal_7530) ) ;
    buf_clk cell_5561 ( .C (clk), .D (signal_7531), .Q (signal_7532) ) ;
    buf_clk cell_5563 ( .C (clk), .D (signal_7533), .Q (signal_7534) ) ;
    buf_clk cell_5565 ( .C (clk), .D (signal_7535), .Q (signal_7536) ) ;
    buf_clk cell_5567 ( .C (clk), .D (signal_7537), .Q (signal_7538) ) ;
    buf_clk cell_5569 ( .C (clk), .D (signal_7539), .Q (signal_7540) ) ;
    buf_clk cell_5571 ( .C (clk), .D (signal_7541), .Q (signal_7542) ) ;
    buf_clk cell_5573 ( .C (clk), .D (signal_7543), .Q (signal_7544) ) ;
    buf_clk cell_5575 ( .C (clk), .D (signal_7545), .Q (signal_7546) ) ;
    buf_clk cell_5577 ( .C (clk), .D (signal_7547), .Q (signal_7548) ) ;
    buf_clk cell_5579 ( .C (clk), .D (signal_7549), .Q (signal_7550) ) ;
    buf_clk cell_5581 ( .C (clk), .D (signal_7551), .Q (signal_7552) ) ;
    buf_clk cell_5583 ( .C (clk), .D (signal_7553), .Q (signal_7554) ) ;
    buf_clk cell_5585 ( .C (clk), .D (signal_7555), .Q (signal_7556) ) ;
    buf_clk cell_5587 ( .C (clk), .D (signal_7557), .Q (signal_7558) ) ;
    buf_clk cell_5589 ( .C (clk), .D (signal_7559), .Q (signal_7560) ) ;
    buf_clk cell_5591 ( .C (clk), .D (signal_7561), .Q (signal_7562) ) ;
    buf_clk cell_5593 ( .C (clk), .D (signal_7563), .Q (signal_7564) ) ;
    buf_clk cell_5595 ( .C (clk), .D (signal_7565), .Q (signal_7566) ) ;
    buf_clk cell_5597 ( .C (clk), .D (signal_7567), .Q (signal_7568) ) ;
    buf_clk cell_5599 ( .C (clk), .D (signal_7569), .Q (signal_7570) ) ;
    buf_clk cell_5601 ( .C (clk), .D (signal_7571), .Q (signal_7572) ) ;
    buf_clk cell_5603 ( .C (clk), .D (signal_7573), .Q (signal_7574) ) ;
    buf_clk cell_5605 ( .C (clk), .D (signal_7575), .Q (signal_7576) ) ;
    buf_clk cell_5607 ( .C (clk), .D (signal_7577), .Q (signal_7578) ) ;
    buf_clk cell_5609 ( .C (clk), .D (signal_7579), .Q (signal_7580) ) ;
    buf_clk cell_5611 ( .C (clk), .D (signal_7581), .Q (signal_7582) ) ;
    buf_clk cell_5613 ( .C (clk), .D (signal_7583), .Q (signal_7584) ) ;
    buf_clk cell_5615 ( .C (clk), .D (signal_7585), .Q (signal_7586) ) ;
    buf_clk cell_5617 ( .C (clk), .D (signal_7587), .Q (signal_7588) ) ;
    buf_clk cell_5619 ( .C (clk), .D (signal_7589), .Q (signal_7590) ) ;
    buf_clk cell_5621 ( .C (clk), .D (signal_7591), .Q (signal_7592) ) ;
    buf_clk cell_5623 ( .C (clk), .D (signal_7593), .Q (signal_7594) ) ;
    buf_clk cell_5625 ( .C (clk), .D (signal_7595), .Q (signal_7596) ) ;
    buf_clk cell_5627 ( .C (clk), .D (signal_7597), .Q (signal_7598) ) ;
    buf_clk cell_5629 ( .C (clk), .D (signal_7599), .Q (signal_7600) ) ;
    buf_clk cell_5631 ( .C (clk), .D (signal_7601), .Q (signal_7602) ) ;
    buf_clk cell_5633 ( .C (clk), .D (signal_7603), .Q (signal_7604) ) ;
    buf_clk cell_5635 ( .C (clk), .D (signal_7605), .Q (signal_7606) ) ;
    buf_clk cell_5637 ( .C (clk), .D (signal_7607), .Q (signal_7608) ) ;
    buf_clk cell_5639 ( .C (clk), .D (signal_7609), .Q (signal_7610) ) ;
    buf_clk cell_5641 ( .C (clk), .D (signal_7611), .Q (signal_7612) ) ;
    buf_clk cell_5643 ( .C (clk), .D (signal_7613), .Q (signal_7614) ) ;
    buf_clk cell_5645 ( .C (clk), .D (signal_7615), .Q (signal_7616) ) ;
    buf_clk cell_5647 ( .C (clk), .D (signal_7617), .Q (signal_7618) ) ;
    buf_clk cell_5649 ( .C (clk), .D (signal_7619), .Q (signal_7620) ) ;
    buf_clk cell_5651 ( .C (clk), .D (signal_7621), .Q (signal_7622) ) ;
    buf_clk cell_5653 ( .C (clk), .D (signal_7623), .Q (signal_7624) ) ;
    buf_clk cell_5655 ( .C (clk), .D (signal_7625), .Q (signal_7626) ) ;
    buf_clk cell_5657 ( .C (clk), .D (signal_7627), .Q (signal_7628) ) ;
    buf_clk cell_5659 ( .C (clk), .D (signal_7629), .Q (signal_7630) ) ;
    buf_clk cell_5661 ( .C (clk), .D (signal_7631), .Q (signal_7632) ) ;
    buf_clk cell_5663 ( .C (clk), .D (signal_7633), .Q (signal_7634) ) ;
    buf_clk cell_5665 ( .C (clk), .D (signal_7635), .Q (signal_7636) ) ;
    buf_clk cell_5667 ( .C (clk), .D (signal_7637), .Q (signal_7638) ) ;
    buf_clk cell_5669 ( .C (clk), .D (signal_7639), .Q (signal_7640) ) ;
    buf_clk cell_5671 ( .C (clk), .D (signal_7641), .Q (signal_7642) ) ;
    buf_clk cell_5673 ( .C (clk), .D (signal_7643), .Q (signal_7644) ) ;
    buf_clk cell_5675 ( .C (clk), .D (signal_7645), .Q (signal_7646) ) ;
    buf_clk cell_5677 ( .C (clk), .D (signal_7647), .Q (signal_7648) ) ;
    buf_clk cell_5679 ( .C (clk), .D (signal_7649), .Q (signal_7650) ) ;
    buf_clk cell_5681 ( .C (clk), .D (signal_7651), .Q (signal_7652) ) ;
    buf_clk cell_5683 ( .C (clk), .D (signal_7653), .Q (signal_7654) ) ;
    buf_clk cell_5685 ( .C (clk), .D (signal_7655), .Q (signal_7656) ) ;
    buf_clk cell_5687 ( .C (clk), .D (signal_7657), .Q (signal_7658) ) ;
    buf_clk cell_5689 ( .C (clk), .D (signal_7659), .Q (signal_7660) ) ;
    buf_clk cell_5691 ( .C (clk), .D (signal_7661), .Q (signal_7662) ) ;
    buf_clk cell_5693 ( .C (clk), .D (signal_7663), .Q (signal_7664) ) ;
    buf_clk cell_5695 ( .C (clk), .D (signal_7665), .Q (signal_7666) ) ;
    buf_clk cell_5697 ( .C (clk), .D (signal_7667), .Q (signal_7668) ) ;
    buf_clk cell_5699 ( .C (clk), .D (signal_7669), .Q (signal_7670) ) ;
    buf_clk cell_5701 ( .C (clk), .D (signal_7671), .Q (signal_7672) ) ;
    buf_clk cell_5703 ( .C (clk), .D (signal_7673), .Q (signal_7674) ) ;
    buf_clk cell_5705 ( .C (clk), .D (signal_7675), .Q (signal_7676) ) ;
    buf_clk cell_5707 ( .C (clk), .D (signal_7677), .Q (signal_7678) ) ;
    buf_clk cell_5709 ( .C (clk), .D (signal_7679), .Q (signal_7680) ) ;
    buf_clk cell_5711 ( .C (clk), .D (signal_7681), .Q (signal_7682) ) ;
    buf_clk cell_5713 ( .C (clk), .D (signal_7683), .Q (signal_7684) ) ;
    buf_clk cell_5715 ( .C (clk), .D (signal_7685), .Q (signal_7686) ) ;
    buf_clk cell_5717 ( .C (clk), .D (signal_7687), .Q (signal_7688) ) ;
    buf_clk cell_5719 ( .C (clk), .D (signal_7689), .Q (signal_7690) ) ;
    buf_clk cell_5721 ( .C (clk), .D (signal_7691), .Q (signal_7692) ) ;
    buf_clk cell_5723 ( .C (clk), .D (signal_7693), .Q (signal_7694) ) ;
    buf_clk cell_5725 ( .C (clk), .D (signal_7695), .Q (signal_7696) ) ;
    buf_clk cell_5727 ( .C (clk), .D (signal_7697), .Q (signal_7698) ) ;
    buf_clk cell_5729 ( .C (clk), .D (signal_7699), .Q (signal_7700) ) ;
    buf_clk cell_5731 ( .C (clk), .D (signal_7701), .Q (signal_7702) ) ;
    buf_clk cell_5733 ( .C (clk), .D (signal_7703), .Q (signal_7704) ) ;
    buf_clk cell_5735 ( .C (clk), .D (signal_7705), .Q (signal_7706) ) ;
    buf_clk cell_5737 ( .C (clk), .D (signal_7707), .Q (signal_7708) ) ;
    buf_clk cell_5739 ( .C (clk), .D (signal_7709), .Q (signal_7710) ) ;
    buf_clk cell_5741 ( .C (clk), .D (signal_7711), .Q (signal_7712) ) ;
    buf_clk cell_5743 ( .C (clk), .D (signal_7713), .Q (signal_7714) ) ;
    buf_clk cell_5745 ( .C (clk), .D (signal_7715), .Q (signal_7716) ) ;
    buf_clk cell_5747 ( .C (clk), .D (signal_7717), .Q (signal_7718) ) ;
    buf_clk cell_5749 ( .C (clk), .D (signal_7719), .Q (signal_7720) ) ;
    buf_clk cell_5751 ( .C (clk), .D (signal_7721), .Q (signal_7722) ) ;
    buf_clk cell_5753 ( .C (clk), .D (signal_7723), .Q (signal_7724) ) ;
    buf_clk cell_5755 ( .C (clk), .D (signal_7725), .Q (signal_7726) ) ;
    buf_clk cell_5757 ( .C (clk), .D (signal_7727), .Q (signal_7728) ) ;
    buf_clk cell_5759 ( .C (clk), .D (signal_7729), .Q (signal_7730) ) ;
    buf_clk cell_5761 ( .C (clk), .D (signal_7731), .Q (signal_7732) ) ;
    buf_clk cell_5763 ( .C (clk), .D (signal_7733), .Q (signal_7734) ) ;
    buf_clk cell_5765 ( .C (clk), .D (signal_7735), .Q (signal_7736) ) ;
    buf_clk cell_5767 ( .C (clk), .D (signal_7737), .Q (signal_7738) ) ;
    buf_clk cell_5769 ( .C (clk), .D (signal_7739), .Q (signal_7740) ) ;
    buf_clk cell_5771 ( .C (clk), .D (signal_7741), .Q (signal_7742) ) ;
    buf_clk cell_5773 ( .C (clk), .D (signal_7743), .Q (signal_7744) ) ;
    buf_clk cell_5775 ( .C (clk), .D (signal_7745), .Q (signal_7746) ) ;
    buf_clk cell_5777 ( .C (clk), .D (signal_7747), .Q (signal_7748) ) ;
    buf_clk cell_5779 ( .C (clk), .D (signal_7749), .Q (signal_7750) ) ;
    buf_clk cell_5781 ( .C (clk), .D (signal_7751), .Q (signal_7752) ) ;
    buf_clk cell_5783 ( .C (clk), .D (signal_7753), .Q (signal_7754) ) ;
    buf_clk cell_5785 ( .C (clk), .D (signal_7755), .Q (signal_7756) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(1)) cell_293 ( .clk (clk), .D ({signal_5723, signal_421}), .Q ({signal_4549, signal_3870}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_296 ( .clk (clk), .D ({signal_5403, signal_423}), .Q ({signal_4666, signal_3869}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_299 ( .clk (clk), .D ({signal_5405, signal_425}), .Q ({signal_4699, signal_3868}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_302 ( .clk (clk), .D ({signal_5407, signal_427}), .Q ({signal_4732, signal_3867}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_305 ( .clk (clk), .D ({signal_5409, signal_429}), .Q ({signal_4765, signal_3866}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_308 ( .clk (clk), .D ({signal_5411, signal_431}), .Q ({signal_4798, signal_3865}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_311 ( .clk (clk), .D ({signal_5413, signal_433}), .Q ({signal_4831, signal_3864}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_314 ( .clk (clk), .D ({signal_5415, signal_435}), .Q ({signal_4864, signal_3863}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_317 ( .clk (clk), .D ({signal_5417, signal_437}), .Q ({signal_4897, signal_3862}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_320 ( .clk (clk), .D ({signal_5725, signal_439}), .Q ({signal_4930, signal_3861}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_323 ( .clk (clk), .D ({signal_5419, signal_441}), .Q ({signal_4582, signal_3860}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_326 ( .clk (clk), .D ({signal_5421, signal_443}), .Q ({signal_4615, signal_3859}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_329 ( .clk (clk), .D ({signal_5423, signal_445}), .Q ({signal_4642, signal_3858}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_332 ( .clk (clk), .D ({signal_5425, signal_447}), .Q ({signal_4645, signal_3857}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_335 ( .clk (clk), .D ({signal_5427, signal_449}), .Q ({signal_4648, signal_3856}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_338 ( .clk (clk), .D ({signal_5429, signal_451}), .Q ({signal_4651, signal_3855}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_341 ( .clk (clk), .D ({signal_5431, signal_453}), .Q ({signal_4654, signal_3854}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_344 ( .clk (clk), .D ({signal_5433, signal_455}), .Q ({signal_4657, signal_3853}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_347 ( .clk (clk), .D ({signal_5435, signal_457}), .Q ({signal_4660, signal_3852}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_350 ( .clk (clk), .D ({signal_5437, signal_459}), .Q ({signal_4663, signal_3851}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_353 ( .clk (clk), .D ({signal_5439, signal_461}), .Q ({signal_4669, signal_3850}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_356 ( .clk (clk), .D ({signal_5441, signal_463}), .Q ({signal_4672, signal_3849}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_359 ( .clk (clk), .D ({signal_5443, signal_465}), .Q ({signal_4675, signal_3848}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_362 ( .clk (clk), .D ({signal_5445, signal_467}), .Q ({signal_4678, signal_3847}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_365 ( .clk (clk), .D ({signal_5447, signal_469}), .Q ({signal_4681, signal_3846}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_368 ( .clk (clk), .D ({signal_5449, signal_471}), .Q ({signal_4684, signal_3845}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_371 ( .clk (clk), .D ({signal_5451, signal_473}), .Q ({signal_4687, signal_3844}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_374 ( .clk (clk), .D ({signal_5453, signal_475}), .Q ({signal_4690, signal_3843}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_377 ( .clk (clk), .D ({signal_5455, signal_477}), .Q ({signal_4693, signal_3842}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_380 ( .clk (clk), .D ({signal_5457, signal_479}), .Q ({signal_4696, signal_3841}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_383 ( .clk (clk), .D ({signal_5459, signal_481}), .Q ({signal_4702, signal_3840}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_386 ( .clk (clk), .D ({signal_5461, signal_483}), .Q ({signal_4705, signal_3839}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_389 ( .clk (clk), .D ({signal_5727, signal_485}), .Q ({signal_4708, signal_3838}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_392 ( .clk (clk), .D ({signal_5463, signal_487}), .Q ({signal_4711, signal_3837}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_395 ( .clk (clk), .D ({signal_5465, signal_489}), .Q ({signal_4714, signal_3836}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_398 ( .clk (clk), .D ({signal_5467, signal_491}), .Q ({signal_4717, signal_3835}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_401 ( .clk (clk), .D ({signal_5469, signal_493}), .Q ({signal_4720, signal_3834}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_404 ( .clk (clk), .D ({signal_5471, signal_495}), .Q ({signal_4723, signal_3833}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_407 ( .clk (clk), .D ({signal_5473, signal_497}), .Q ({signal_4726, signal_3832}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_410 ( .clk (clk), .D ({signal_5475, signal_499}), .Q ({signal_4729, signal_3831}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_413 ( .clk (clk), .D ({signal_5477, signal_501}), .Q ({signal_4735, signal_3830}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_416 ( .clk (clk), .D ({signal_5729, signal_503}), .Q ({signal_4738, signal_3829}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_419 ( .clk (clk), .D ({signal_5479, signal_505}), .Q ({signal_4741, signal_3828}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_422 ( .clk (clk), .D ({signal_5481, signal_507}), .Q ({signal_4744, signal_3827}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_425 ( .clk (clk), .D ({signal_5483, signal_509}), .Q ({signal_4747, signal_3826}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_428 ( .clk (clk), .D ({signal_5485, signal_511}), .Q ({signal_4750, signal_3825}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_431 ( .clk (clk), .D ({signal_5487, signal_513}), .Q ({signal_4753, signal_3824}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_434 ( .clk (clk), .D ({signal_5489, signal_515}), .Q ({signal_4756, signal_3823}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_437 ( .clk (clk), .D ({signal_5491, signal_517}), .Q ({signal_4759, signal_3822}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_440 ( .clk (clk), .D ({signal_5493, signal_519}), .Q ({signal_4762, signal_3821}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_443 ( .clk (clk), .D ({signal_5495, signal_521}), .Q ({signal_4768, signal_3820}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_446 ( .clk (clk), .D ({signal_5497, signal_523}), .Q ({signal_4771, signal_3819}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_449 ( .clk (clk), .D ({signal_5499, signal_525}), .Q ({signal_4774, signal_3818}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_452 ( .clk (clk), .D ({signal_5501, signal_527}), .Q ({signal_4777, signal_3817}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_455 ( .clk (clk), .D ({signal_5503, signal_529}), .Q ({signal_4780, signal_3816}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_458 ( .clk (clk), .D ({signal_5505, signal_531}), .Q ({signal_4783, signal_3815}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_461 ( .clk (clk), .D ({signal_5507, signal_533}), .Q ({signal_4786, signal_3814}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_464 ( .clk (clk), .D ({signal_5509, signal_535}), .Q ({signal_4789, signal_3813}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_467 ( .clk (clk), .D ({signal_5511, signal_537}), .Q ({signal_4792, signal_3812}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_470 ( .clk (clk), .D ({signal_5513, signal_539}), .Q ({signal_4795, signal_3811}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_473 ( .clk (clk), .D ({signal_5515, signal_541}), .Q ({signal_4801, signal_3810}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_476 ( .clk (clk), .D ({signal_5517, signal_543}), .Q ({signal_4804, signal_3809}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_479 ( .clk (clk), .D ({signal_5519, signal_545}), .Q ({signal_4807, signal_3808}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_482 ( .clk (clk), .D ({signal_5521, signal_547}), .Q ({signal_4810, signal_3807}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_485 ( .clk (clk), .D ({signal_5731, signal_549}), .Q ({signal_4813, signal_3806}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_488 ( .clk (clk), .D ({signal_5523, signal_551}), .Q ({signal_4816, signal_3805}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_491 ( .clk (clk), .D ({signal_5525, signal_553}), .Q ({signal_4819, signal_3804}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_494 ( .clk (clk), .D ({signal_5527, signal_555}), .Q ({signal_4822, signal_3803}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_497 ( .clk (clk), .D ({signal_5529, signal_557}), .Q ({signal_4825, signal_3802}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_500 ( .clk (clk), .D ({signal_5531, signal_559}), .Q ({signal_4828, signal_3801}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_503 ( .clk (clk), .D ({signal_5533, signal_561}), .Q ({signal_4834, signal_3800}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_506 ( .clk (clk), .D ({signal_5535, signal_563}), .Q ({signal_4837, signal_3799}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_509 ( .clk (clk), .D ({signal_5537, signal_565}), .Q ({signal_4840, signal_3798}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_512 ( .clk (clk), .D ({signal_5733, signal_567}), .Q ({signal_4843, signal_3797}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_515 ( .clk (clk), .D ({signal_5539, signal_569}), .Q ({signal_4846, signal_3796}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_518 ( .clk (clk), .D ({signal_5541, signal_571}), .Q ({signal_4849, signal_3795}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_521 ( .clk (clk), .D ({signal_5543, signal_573}), .Q ({signal_4852, signal_3794}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_524 ( .clk (clk), .D ({signal_5545, signal_575}), .Q ({signal_4855, signal_3793}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_527 ( .clk (clk), .D ({signal_5547, signal_577}), .Q ({signal_4858, signal_3792}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_530 ( .clk (clk), .D ({signal_5549, signal_579}), .Q ({signal_4861, signal_3791}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_533 ( .clk (clk), .D ({signal_5551, signal_581}), .Q ({signal_4867, signal_3790}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_536 ( .clk (clk), .D ({signal_5553, signal_583}), .Q ({signal_4870, signal_3789}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_539 ( .clk (clk), .D ({signal_5555, signal_585}), .Q ({signal_4873, signal_3788}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_542 ( .clk (clk), .D ({signal_5557, signal_587}), .Q ({signal_4876, signal_3787}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_545 ( .clk (clk), .D ({signal_5559, signal_589}), .Q ({signal_4879, signal_3786}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_548 ( .clk (clk), .D ({signal_5561, signal_591}), .Q ({signal_4882, signal_3785}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_551 ( .clk (clk), .D ({signal_5563, signal_593}), .Q ({signal_4885, signal_3784}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_554 ( .clk (clk), .D ({signal_5565, signal_595}), .Q ({signal_4888, signal_3783}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_557 ( .clk (clk), .D ({signal_5567, signal_597}), .Q ({signal_4891, signal_3782}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_560 ( .clk (clk), .D ({signal_5569, signal_599}), .Q ({signal_4894, signal_3781}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_563 ( .clk (clk), .D ({signal_5571, signal_601}), .Q ({signal_4900, signal_3780}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_566 ( .clk (clk), .D ({signal_5573, signal_603}), .Q ({signal_4903, signal_3779}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_569 ( .clk (clk), .D ({signal_5575, signal_605}), .Q ({signal_4906, signal_3778}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_572 ( .clk (clk), .D ({signal_5577, signal_607}), .Q ({signal_4909, signal_3777}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_575 ( .clk (clk), .D ({signal_5579, signal_609}), .Q ({signal_4912, signal_3776}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_578 ( .clk (clk), .D ({signal_5581, signal_611}), .Q ({signal_4915, signal_3775}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_581 ( .clk (clk), .D ({signal_5735, signal_613}), .Q ({signal_4918, signal_3774}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_584 ( .clk (clk), .D ({signal_5583, signal_615}), .Q ({signal_4921, signal_3773}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_587 ( .clk (clk), .D ({signal_5585, signal_617}), .Q ({signal_4924, signal_3772}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_590 ( .clk (clk), .D ({signal_5587, signal_619}), .Q ({signal_4927, signal_3771}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_593 ( .clk (clk), .D ({signal_5589, signal_621}), .Q ({signal_4552, signal_3770}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_596 ( .clk (clk), .D ({signal_5591, signal_623}), .Q ({signal_4555, signal_3769}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_599 ( .clk (clk), .D ({signal_5593, signal_625}), .Q ({signal_4558, signal_3768}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_602 ( .clk (clk), .D ({signal_5595, signal_627}), .Q ({signal_4561, signal_3767}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_605 ( .clk (clk), .D ({signal_5597, signal_629}), .Q ({signal_4564, signal_3766}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_608 ( .clk (clk), .D ({signal_5737, signal_631}), .Q ({signal_4567, signal_3765}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_611 ( .clk (clk), .D ({signal_5599, signal_633}), .Q ({signal_4570, signal_3764}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_614 ( .clk (clk), .D ({signal_5601, signal_635}), .Q ({signal_4573, signal_3763}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_617 ( .clk (clk), .D ({signal_5603, signal_637}), .Q ({signal_4576, signal_3762}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_620 ( .clk (clk), .D ({signal_5605, signal_639}), .Q ({signal_4579, signal_3761}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_623 ( .clk (clk), .D ({signal_5607, signal_641}), .Q ({signal_4585, signal_3760}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_626 ( .clk (clk), .D ({signal_5609, signal_643}), .Q ({signal_4588, signal_3759}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_629 ( .clk (clk), .D ({signal_5611, signal_645}), .Q ({signal_4591, signal_3758}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_632 ( .clk (clk), .D ({signal_5613, signal_647}), .Q ({signal_4594, signal_3757}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_635 ( .clk (clk), .D ({signal_5615, signal_649}), .Q ({signal_4597, signal_3756}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_638 ( .clk (clk), .D ({signal_5617, signal_651}), .Q ({signal_4600, signal_3755}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_641 ( .clk (clk), .D ({signal_5619, signal_653}), .Q ({signal_4603, signal_3754}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_644 ( .clk (clk), .D ({signal_5621, signal_655}), .Q ({signal_4606, signal_3753}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_647 ( .clk (clk), .D ({signal_5623, signal_657}), .Q ({signal_4609, signal_3752}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_650 ( .clk (clk), .D ({signal_5625, signal_659}), .Q ({signal_4612, signal_3751}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_653 ( .clk (clk), .D ({signal_5627, signal_661}), .Q ({signal_4618, signal_3750}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_656 ( .clk (clk), .D ({signal_5629, signal_663}), .Q ({signal_4621, signal_3749}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_659 ( .clk (clk), .D ({signal_5631, signal_665}), .Q ({signal_4624, signal_3748}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_662 ( .clk (clk), .D ({signal_5633, signal_667}), .Q ({signal_4627, signal_3747}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_665 ( .clk (clk), .D ({signal_5635, signal_669}), .Q ({signal_4630, signal_3746}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_668 ( .clk (clk), .D ({signal_5637, signal_671}), .Q ({signal_4633, signal_3745}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_671 ( .clk (clk), .D ({signal_5639, signal_673}), .Q ({signal_4636, signal_3744}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_674 ( .clk (clk), .D ({signal_5641, signal_675}), .Q ({signal_4639, signal_3743}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3157 ( .clk (clk), .D ({signal_5925, signal_2853}), .Q ({signal_4550, signal_4378}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3160 ( .clk (clk), .D ({signal_5927, signal_2855}), .Q ({signal_4667, signal_4377}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3163 ( .clk (clk), .D ({signal_5929, signal_2857}), .Q ({signal_4700, signal_4376}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3166 ( .clk (clk), .D ({signal_5931, signal_2859}), .Q ({signal_4733, signal_4375}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3169 ( .clk (clk), .D ({signal_5933, signal_2861}), .Q ({signal_4766, signal_4374}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3172 ( .clk (clk), .D ({signal_5935, signal_2863}), .Q ({signal_4799, signal_4373}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3175 ( .clk (clk), .D ({signal_5937, signal_2865}), .Q ({signal_4832, signal_4372}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3178 ( .clk (clk), .D ({signal_5939, signal_2867}), .Q ({signal_4865, signal_4371}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3181 ( .clk (clk), .D ({signal_5941, signal_2869}), .Q ({signal_4898, signal_4370}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3184 ( .clk (clk), .D ({signal_5943, signal_2871}), .Q ({signal_4931, signal_4369}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3187 ( .clk (clk), .D ({signal_5945, signal_2873}), .Q ({signal_4583, signal_4368}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3190 ( .clk (clk), .D ({signal_5947, signal_2875}), .Q ({signal_4616, signal_4367}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3193 ( .clk (clk), .D ({signal_5949, signal_2877}), .Q ({signal_4643, signal_4366}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3196 ( .clk (clk), .D ({signal_5951, signal_2879}), .Q ({signal_4646, signal_4365}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3199 ( .clk (clk), .D ({signal_5953, signal_2881}), .Q ({signal_4649, signal_4364}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3202 ( .clk (clk), .D ({signal_5955, signal_2883}), .Q ({signal_4652, signal_4363}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3205 ( .clk (clk), .D ({signal_5957, signal_2885}), .Q ({signal_4655, signal_4362}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3208 ( .clk (clk), .D ({signal_5959, signal_2887}), .Q ({signal_4658, signal_4361}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3211 ( .clk (clk), .D ({signal_5961, signal_2889}), .Q ({signal_4661, signal_4360}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3214 ( .clk (clk), .D ({signal_5963, signal_2891}), .Q ({signal_4664, signal_4359}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3217 ( .clk (clk), .D ({signal_5965, signal_2893}), .Q ({signal_4670, signal_4358}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3220 ( .clk (clk), .D ({signal_5967, signal_2895}), .Q ({signal_4673, signal_4357}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3223 ( .clk (clk), .D ({signal_5969, signal_2897}), .Q ({signal_4676, signal_4356}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3226 ( .clk (clk), .D ({signal_5971, signal_2899}), .Q ({signal_4679, signal_4355}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3229 ( .clk (clk), .D ({signal_5997, signal_2901}), .Q ({signal_4682, signal_4354}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3232 ( .clk (clk), .D ({signal_5999, signal_2903}), .Q ({signal_4685, signal_4353}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3235 ( .clk (clk), .D ({signal_6016, signal_2905}), .Q ({signal_4688, signal_4352}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3238 ( .clk (clk), .D ({signal_6018, signal_2907}), .Q ({signal_4691, signal_4351}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3241 ( .clk (clk), .D ({signal_6001, signal_2909}), .Q ({signal_4694, signal_4350}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3244 ( .clk (clk), .D ({signal_6020, signal_2911}), .Q ({signal_4697, signal_4349}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3247 ( .clk (clk), .D ({signal_6003, signal_2913}), .Q ({signal_4703, signal_4348}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3250 ( .clk (clk), .D ({signal_6005, signal_2915}), .Q ({signal_4706, signal_4347}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3253 ( .clk (clk), .D ({signal_5829, signal_2917}), .Q ({signal_4709, signal_4346}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3256 ( .clk (clk), .D ({signal_5831, signal_2919}), .Q ({signal_4712, signal_4345}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3259 ( .clk (clk), .D ({signal_5833, signal_2921}), .Q ({signal_4715, signal_4344}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3262 ( .clk (clk), .D ({signal_5835, signal_2923}), .Q ({signal_4718, signal_4343}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3265 ( .clk (clk), .D ({signal_5837, signal_2925}), .Q ({signal_4721, signal_4342}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3268 ( .clk (clk), .D ({signal_5839, signal_2927}), .Q ({signal_4724, signal_4341}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3271 ( .clk (clk), .D ({signal_5841, signal_2929}), .Q ({signal_4727, signal_4340}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3274 ( .clk (clk), .D ({signal_5843, signal_2931}), .Q ({signal_4730, signal_4339}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3277 ( .clk (clk), .D ({signal_5845, signal_2933}), .Q ({signal_4736, signal_4338}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3280 ( .clk (clk), .D ({signal_5847, signal_2935}), .Q ({signal_4739, signal_4337}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3283 ( .clk (clk), .D ({signal_5849, signal_2937}), .Q ({signal_4742, signal_4336}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3286 ( .clk (clk), .D ({signal_5851, signal_2939}), .Q ({signal_4745, signal_4335}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3289 ( .clk (clk), .D ({signal_5853, signal_2941}), .Q ({signal_4748, signal_4334}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3292 ( .clk (clk), .D ({signal_5855, signal_2943}), .Q ({signal_4751, signal_4333}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3295 ( .clk (clk), .D ({signal_5857, signal_2945}), .Q ({signal_4754, signal_4332}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3298 ( .clk (clk), .D ({signal_5859, signal_2947}), .Q ({signal_4757, signal_4331}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3301 ( .clk (clk), .D ({signal_5861, signal_2949}), .Q ({signal_4760, signal_4330}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3304 ( .clk (clk), .D ({signal_5863, signal_2951}), .Q ({signal_4763, signal_4329}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3307 ( .clk (clk), .D ({signal_5865, signal_2953}), .Q ({signal_4769, signal_4328}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3310 ( .clk (clk), .D ({signal_5867, signal_2955}), .Q ({signal_4772, signal_4327}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3313 ( .clk (clk), .D ({signal_5869, signal_2957}), .Q ({signal_4775, signal_4326}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3316 ( .clk (clk), .D ({signal_5871, signal_2959}), .Q ({signal_4778, signal_4325}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3319 ( .clk (clk), .D ({signal_5873, signal_2961}), .Q ({signal_4781, signal_4324}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3322 ( .clk (clk), .D ({signal_5875, signal_2963}), .Q ({signal_4784, signal_4323}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3325 ( .clk (clk), .D ({signal_5973, signal_2965}), .Q ({signal_4787, signal_4322}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3328 ( .clk (clk), .D ({signal_5975, signal_2967}), .Q ({signal_4790, signal_4321}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3331 ( .clk (clk), .D ({signal_6007, signal_2969}), .Q ({signal_4793, signal_4320}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3334 ( .clk (clk), .D ({signal_6009, signal_2971}), .Q ({signal_4796, signal_4319}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3337 ( .clk (clk), .D ({signal_5977, signal_2973}), .Q ({signal_4802, signal_4318}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3340 ( .clk (clk), .D ({signal_6011, signal_2975}), .Q ({signal_4805, signal_4317}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3343 ( .clk (clk), .D ({signal_5979, signal_2977}), .Q ({signal_4808, signal_4316}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3346 ( .clk (clk), .D ({signal_5981, signal_2979}), .Q ({signal_4811, signal_4315}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3349 ( .clk (clk), .D ({signal_5739, signal_2981}), .Q ({signal_4814, signal_4314}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3352 ( .clk (clk), .D ({signal_5741, signal_2983}), .Q ({signal_4817, signal_4313}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3355 ( .clk (clk), .D ({signal_5743, signal_2985}), .Q ({signal_4820, signal_4312}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3358 ( .clk (clk), .D ({signal_5745, signal_2987}), .Q ({signal_4823, signal_4311}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3361 ( .clk (clk), .D ({signal_5747, signal_2989}), .Q ({signal_4826, signal_4310}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3364 ( .clk (clk), .D ({signal_5749, signal_2991}), .Q ({signal_4829, signal_4309}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3367 ( .clk (clk), .D ({signal_5751, signal_2993}), .Q ({signal_4835, signal_4308}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3370 ( .clk (clk), .D ({signal_5753, signal_2995}), .Q ({signal_4838, signal_4307}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3373 ( .clk (clk), .D ({signal_5755, signal_2997}), .Q ({signal_4841, signal_4306}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3376 ( .clk (clk), .D ({signal_5757, signal_2999}), .Q ({signal_4844, signal_4305}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3379 ( .clk (clk), .D ({signal_5759, signal_3001}), .Q ({signal_4847, signal_4304}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3382 ( .clk (clk), .D ({signal_5761, signal_3003}), .Q ({signal_4850, signal_4303}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3385 ( .clk (clk), .D ({signal_5763, signal_3005}), .Q ({signal_4853, signal_4302}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3388 ( .clk (clk), .D ({signal_5765, signal_3007}), .Q ({signal_4856, signal_4301}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3391 ( .clk (clk), .D ({signal_5767, signal_3009}), .Q ({signal_4859, signal_4300}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3394 ( .clk (clk), .D ({signal_5769, signal_3011}), .Q ({signal_4862, signal_4299}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3397 ( .clk (clk), .D ({signal_5771, signal_3013}), .Q ({signal_4868, signal_4298}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3400 ( .clk (clk), .D ({signal_5773, signal_3015}), .Q ({signal_4871, signal_4297}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3403 ( .clk (clk), .D ({signal_5775, signal_3017}), .Q ({signal_4874, signal_4296}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3406 ( .clk (clk), .D ({signal_5777, signal_3019}), .Q ({signal_4877, signal_4295}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3409 ( .clk (clk), .D ({signal_5779, signal_3021}), .Q ({signal_4880, signal_4294}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3412 ( .clk (clk), .D ({signal_5781, signal_3023}), .Q ({signal_4883, signal_4293}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3415 ( .clk (clk), .D ({signal_5783, signal_3025}), .Q ({signal_4886, signal_4292}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3418 ( .clk (clk), .D ({signal_5785, signal_3027}), .Q ({signal_4889, signal_4291}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3421 ( .clk (clk), .D ({signal_5877, signal_3029}), .Q ({signal_4892, signal_4290}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3424 ( .clk (clk), .D ({signal_5879, signal_3031}), .Q ({signal_4895, signal_4289}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3427 ( .clk (clk), .D ({signal_5983, signal_3033}), .Q ({signal_4901, signal_4288}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3430 ( .clk (clk), .D ({signal_5985, signal_3035}), .Q ({signal_4904, signal_4287}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3433 ( .clk (clk), .D ({signal_5881, signal_3037}), .Q ({signal_4907, signal_4286}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3436 ( .clk (clk), .D ({signal_5987, signal_3039}), .Q ({signal_4910, signal_4285}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3439 ( .clk (clk), .D ({signal_5883, signal_3041}), .Q ({signal_4913, signal_4284}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3442 ( .clk (clk), .D ({signal_5885, signal_3043}), .Q ({signal_4916, signal_4283}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3445 ( .clk (clk), .D ({signal_5643, signal_3045}), .Q ({signal_4919, signal_4282}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3448 ( .clk (clk), .D ({signal_5645, signal_3047}), .Q ({signal_4922, signal_4281}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3451 ( .clk (clk), .D ({signal_5647, signal_3049}), .Q ({signal_4925, signal_4280}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3454 ( .clk (clk), .D ({signal_5649, signal_3051}), .Q ({signal_4928, signal_4279}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3457 ( .clk (clk), .D ({signal_5651, signal_3053}), .Q ({signal_4553, signal_4278}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3460 ( .clk (clk), .D ({signal_5653, signal_3055}), .Q ({signal_4556, signal_4277}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3463 ( .clk (clk), .D ({signal_5655, signal_3057}), .Q ({signal_4559, signal_4276}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3466 ( .clk (clk), .D ({signal_5657, signal_3059}), .Q ({signal_4562, signal_4275}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3469 ( .clk (clk), .D ({signal_5659, signal_3061}), .Q ({signal_4565, signal_4274}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3472 ( .clk (clk), .D ({signal_5661, signal_3063}), .Q ({signal_4568, signal_4273}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3475 ( .clk (clk), .D ({signal_5663, signal_3065}), .Q ({signal_4571, signal_4272}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3478 ( .clk (clk), .D ({signal_5665, signal_3067}), .Q ({signal_4574, signal_4271}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3481 ( .clk (clk), .D ({signal_5667, signal_3069}), .Q ({signal_4577, signal_4270}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3484 ( .clk (clk), .D ({signal_5669, signal_3071}), .Q ({signal_4580, signal_4269}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3487 ( .clk (clk), .D ({signal_5671, signal_3073}), .Q ({signal_4586, signal_4268}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3490 ( .clk (clk), .D ({signal_5673, signal_3075}), .Q ({signal_4589, signal_4267}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3493 ( .clk (clk), .D ({signal_5675, signal_3077}), .Q ({signal_4592, signal_4266}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3496 ( .clk (clk), .D ({signal_5677, signal_3079}), .Q ({signal_4595, signal_4265}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3499 ( .clk (clk), .D ({signal_5679, signal_3081}), .Q ({signal_4598, signal_4264}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3502 ( .clk (clk), .D ({signal_5681, signal_3083}), .Q ({signal_4601, signal_4263}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3505 ( .clk (clk), .D ({signal_5683, signal_3085}), .Q ({signal_4604, signal_4262}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3508 ( .clk (clk), .D ({signal_5685, signal_3087}), .Q ({signal_4607, signal_4261}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3511 ( .clk (clk), .D ({signal_5687, signal_3089}), .Q ({signal_4610, signal_4260}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3514 ( .clk (clk), .D ({signal_5689, signal_3091}), .Q ({signal_4613, signal_4259}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3517 ( .clk (clk), .D ({signal_5787, signal_3093}), .Q ({signal_4619, signal_4258}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3520 ( .clk (clk), .D ({signal_5789, signal_3095}), .Q ({signal_4622, signal_4257}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3523 ( .clk (clk), .D ({signal_5887, signal_3097}), .Q ({signal_4625, signal_4256}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3526 ( .clk (clk), .D ({signal_5889, signal_3099}), .Q ({signal_4628, signal_4255}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3529 ( .clk (clk), .D ({signal_5791, signal_3101}), .Q ({signal_4631, signal_4254}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3532 ( .clk (clk), .D ({signal_5891, signal_3103}), .Q ({signal_4634, signal_4253}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3535 ( .clk (clk), .D ({signal_5793, signal_3105}), .Q ({signal_4637, signal_4252}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_3538 ( .clk (clk), .D ({signal_5795, signal_3107}), .Q ({signal_4640, signal_4251}) ) ;
    DFF_X1 cell_4202 ( .CK (clk), .D (signal_7750), .Q (signal_4388), .QN () ) ;
    DFF_X1 cell_4204 ( .CK (clk), .D (signal_7752), .Q (signal_4387), .QN () ) ;
    DFF_X1 cell_4206 ( .CK (clk), .D (signal_7754), .Q (signal_4386), .QN () ) ;
    DFF_X1 cell_4208 ( .CK (clk), .D (signal_7756), .Q (signal_4385), .QN () ) ;
endmodule
