/* modified netlist. Source: module SkinnyTop in file Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* 1 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 2 register stage(s) in total */

module SkinnyTop_GHPCLL_ANF_Pipeline_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [1023:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_943 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1485 ;
    wire signal_1487 ;
    wire signal_1489 ;
    wire signal_1491 ;
    wire signal_1493 ;
    wire signal_1495 ;
    wire signal_1497 ;
    wire signal_1499 ;
    wire signal_1501 ;
    wire signal_1503 ;
    wire signal_1505 ;
    wire signal_1507 ;
    wire signal_1509 ;
    wire signal_1511 ;
    wire signal_1513 ;
    wire signal_1515 ;
    wire signal_1517 ;
    wire signal_1519 ;
    wire signal_1521 ;
    wire signal_1523 ;
    wire signal_1525 ;
    wire signal_1527 ;
    wire signal_1529 ;
    wire signal_1531 ;
    wire signal_1533 ;
    wire signal_1535 ;
    wire signal_1537 ;
    wire signal_1539 ;
    wire signal_1541 ;
    wire signal_1543 ;
    wire signal_1545 ;
    wire signal_1547 ;
    wire signal_1549 ;
    wire signal_1551 ;
    wire signal_1553 ;
    wire signal_1555 ;
    wire signal_1557 ;
    wire signal_1559 ;
    wire signal_1561 ;
    wire signal_1563 ;
    wire signal_1565 ;
    wire signal_1567 ;
    wire signal_1569 ;
    wire signal_1571 ;
    wire signal_1573 ;
    wire signal_1575 ;
    wire signal_1577 ;
    wire signal_1579 ;
    wire signal_1581 ;
    wire signal_1583 ;
    wire signal_1585 ;
    wire signal_1587 ;
    wire signal_1589 ;
    wire signal_1591 ;
    wire signal_1593 ;
    wire signal_1595 ;
    wire signal_1597 ;
    wire signal_1599 ;
    wire signal_1601 ;
    wire signal_1603 ;
    wire signal_1605 ;
    wire signal_1607 ;
    wire signal_1609 ;
    wire signal_1611 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;

    /* cells in depth 0 */
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_769 ( .s (rst), .b ({signal_1164, signal_1163}), .a ({Key_s1[0], Key_s0[0]}), .c ({signal_1166, signal_1099}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_770 ( .s (rst), .b ({signal_1167, signal_1162}), .a ({Key_s1[1], Key_s0[1]}), .c ({signal_1169, signal_1098}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_771 ( .s (rst), .b ({signal_1170, signal_1161}), .a ({Key_s1[2], Key_s0[2]}), .c ({signal_1172, signal_1097}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_772 ( .s (rst), .b ({signal_1173, signal_1160}), .a ({Key_s1[3], Key_s0[3]}), .c ({signal_1175, signal_1096}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_773 ( .s (rst), .b ({signal_1176, signal_1159}), .a ({Key_s1[4], Key_s0[4]}), .c ({signal_1178, signal_1095}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_774 ( .s (rst), .b ({signal_1179, signal_1158}), .a ({Key_s1[5], Key_s0[5]}), .c ({signal_1181, signal_1094}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_775 ( .s (rst), .b ({signal_1182, signal_1157}), .a ({Key_s1[6], Key_s0[6]}), .c ({signal_1184, signal_1093}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_776 ( .s (rst), .b ({signal_1185, signal_1156}), .a ({Key_s1[7], Key_s0[7]}), .c ({signal_1187, signal_1092}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_777 ( .s (rst), .b ({signal_1188, signal_1155}), .a ({Key_s1[8], Key_s0[8]}), .c ({signal_1190, signal_1091}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_778 ( .s (rst), .b ({signal_1191, signal_1154}), .a ({Key_s1[9], Key_s0[9]}), .c ({signal_1193, signal_1090}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_779 ( .s (rst), .b ({signal_1194, signal_1153}), .a ({Key_s1[10], Key_s0[10]}), .c ({signal_1196, signal_1089}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_780 ( .s (rst), .b ({signal_1197, signal_1152}), .a ({Key_s1[11], Key_s0[11]}), .c ({signal_1199, signal_1088}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_781 ( .s (rst), .b ({signal_1200, signal_1151}), .a ({Key_s1[12], Key_s0[12]}), .c ({signal_1202, signal_1087}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_782 ( .s (rst), .b ({signal_1203, signal_1150}), .a ({Key_s1[13], Key_s0[13]}), .c ({signal_1205, signal_1086}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_783 ( .s (rst), .b ({signal_1206, signal_1149}), .a ({Key_s1[14], Key_s0[14]}), .c ({signal_1208, signal_1085}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_784 ( .s (rst), .b ({signal_1209, signal_1148}), .a ({Key_s1[15], Key_s0[15]}), .c ({signal_1211, signal_1084}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_785 ( .s (rst), .b ({signal_1212, signal_1147}), .a ({Key_s1[16], Key_s0[16]}), .c ({signal_1214, signal_1083}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_786 ( .s (rst), .b ({signal_1215, signal_1146}), .a ({Key_s1[17], Key_s0[17]}), .c ({signal_1217, signal_1082}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_787 ( .s (rst), .b ({signal_1218, signal_1145}), .a ({Key_s1[18], Key_s0[18]}), .c ({signal_1220, signal_1081}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_788 ( .s (rst), .b ({signal_1221, signal_1144}), .a ({Key_s1[19], Key_s0[19]}), .c ({signal_1223, signal_1080}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_789 ( .s (rst), .b ({signal_1224, signal_1143}), .a ({Key_s1[20], Key_s0[20]}), .c ({signal_1226, signal_1079}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_790 ( .s (rst), .b ({signal_1227, signal_1142}), .a ({Key_s1[21], Key_s0[21]}), .c ({signal_1229, signal_1078}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_791 ( .s (rst), .b ({signal_1230, signal_1141}), .a ({Key_s1[22], Key_s0[22]}), .c ({signal_1232, signal_1077}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_792 ( .s (rst), .b ({signal_1233, signal_1140}), .a ({Key_s1[23], Key_s0[23]}), .c ({signal_1235, signal_1076}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_793 ( .s (rst), .b ({signal_1236, signal_1139}), .a ({Key_s1[24], Key_s0[24]}), .c ({signal_1238, signal_1075}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_794 ( .s (rst), .b ({signal_1239, signal_1138}), .a ({Key_s1[25], Key_s0[25]}), .c ({signal_1241, signal_1074}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_795 ( .s (rst), .b ({signal_1242, signal_1137}), .a ({Key_s1[26], Key_s0[26]}), .c ({signal_1244, signal_1073}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_796 ( .s (rst), .b ({signal_1245, signal_1136}), .a ({Key_s1[27], Key_s0[27]}), .c ({signal_1247, signal_1072}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_797 ( .s (rst), .b ({signal_1248, signal_1135}), .a ({Key_s1[28], Key_s0[28]}), .c ({signal_1250, signal_1071}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_798 ( .s (rst), .b ({signal_1251, signal_1134}), .a ({Key_s1[29], Key_s0[29]}), .c ({signal_1253, signal_1070}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_799 ( .s (rst), .b ({signal_1254, signal_1133}), .a ({Key_s1[30], Key_s0[30]}), .c ({signal_1256, signal_1069}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_800 ( .s (rst), .b ({signal_1257, signal_1132}), .a ({Key_s1[31], Key_s0[31]}), .c ({signal_1259, signal_1068}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_801 ( .s (rst), .b ({signal_1260, signal_1131}), .a ({Key_s1[32], Key_s0[32]}), .c ({signal_1262, signal_1067}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_802 ( .s (rst), .b ({signal_1263, signal_1130}), .a ({Key_s1[33], Key_s0[33]}), .c ({signal_1265, signal_1066}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_803 ( .s (rst), .b ({signal_1266, signal_1129}), .a ({Key_s1[34], Key_s0[34]}), .c ({signal_1268, signal_1065}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_804 ( .s (rst), .b ({signal_1269, signal_1128}), .a ({Key_s1[35], Key_s0[35]}), .c ({signal_1271, signal_1064}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_805 ( .s (rst), .b ({signal_1272, signal_1127}), .a ({Key_s1[36], Key_s0[36]}), .c ({signal_1274, signal_1063}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_806 ( .s (rst), .b ({signal_1275, signal_1126}), .a ({Key_s1[37], Key_s0[37]}), .c ({signal_1277, signal_1062}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_807 ( .s (rst), .b ({signal_1278, signal_1125}), .a ({Key_s1[38], Key_s0[38]}), .c ({signal_1280, signal_1061}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_808 ( .s (rst), .b ({signal_1281, signal_1124}), .a ({Key_s1[39], Key_s0[39]}), .c ({signal_1283, signal_1060}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_809 ( .s (rst), .b ({signal_1284, signal_1123}), .a ({Key_s1[40], Key_s0[40]}), .c ({signal_1286, signal_1059}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_810 ( .s (rst), .b ({signal_1287, signal_1122}), .a ({Key_s1[41], Key_s0[41]}), .c ({signal_1289, signal_1058}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_811 ( .s (rst), .b ({signal_1290, signal_1121}), .a ({Key_s1[42], Key_s0[42]}), .c ({signal_1292, signal_1057}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_812 ( .s (rst), .b ({signal_1293, signal_1120}), .a ({Key_s1[43], Key_s0[43]}), .c ({signal_1295, signal_1056}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_813 ( .s (rst), .b ({signal_1296, signal_1119}), .a ({Key_s1[44], Key_s0[44]}), .c ({signal_1298, signal_1055}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_814 ( .s (rst), .b ({signal_1299, signal_1118}), .a ({Key_s1[45], Key_s0[45]}), .c ({signal_1301, signal_1054}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_815 ( .s (rst), .b ({signal_1302, signal_1117}), .a ({Key_s1[46], Key_s0[46]}), .c ({signal_1304, signal_1053}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_816 ( .s (rst), .b ({signal_1305, signal_1116}), .a ({Key_s1[47], Key_s0[47]}), .c ({signal_1307, signal_1052}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_817 ( .s (rst), .b ({signal_1308, signal_1115}), .a ({Key_s1[48], Key_s0[48]}), .c ({signal_1310, signal_1051}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_818 ( .s (rst), .b ({signal_1311, signal_1114}), .a ({Key_s1[49], Key_s0[49]}), .c ({signal_1313, signal_1050}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_819 ( .s (rst), .b ({signal_1314, signal_1113}), .a ({Key_s1[50], Key_s0[50]}), .c ({signal_1316, signal_1049}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_820 ( .s (rst), .b ({signal_1317, signal_1112}), .a ({Key_s1[51], Key_s0[51]}), .c ({signal_1319, signal_1048}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_821 ( .s (rst), .b ({signal_1320, signal_1111}), .a ({Key_s1[52], Key_s0[52]}), .c ({signal_1322, signal_1047}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_822 ( .s (rst), .b ({signal_1323, signal_1110}), .a ({Key_s1[53], Key_s0[53]}), .c ({signal_1325, signal_1046}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_823 ( .s (rst), .b ({signal_1326, signal_1109}), .a ({Key_s1[54], Key_s0[54]}), .c ({signal_1328, signal_1045}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_824 ( .s (rst), .b ({signal_1329, signal_1108}), .a ({Key_s1[55], Key_s0[55]}), .c ({signal_1331, signal_1044}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_825 ( .s (rst), .b ({signal_1332, signal_1107}), .a ({Key_s1[56], Key_s0[56]}), .c ({signal_1334, signal_1043}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_826 ( .s (rst), .b ({signal_1335, signal_1106}), .a ({Key_s1[57], Key_s0[57]}), .c ({signal_1337, signal_1042}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_827 ( .s (rst), .b ({signal_1338, signal_1105}), .a ({Key_s1[58], Key_s0[58]}), .c ({signal_1340, signal_1041}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_828 ( .s (rst), .b ({signal_1341, signal_1104}), .a ({Key_s1[59], Key_s0[59]}), .c ({signal_1343, signal_1040}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_829 ( .s (rst), .b ({signal_1344, signal_1103}), .a ({Key_s1[60], Key_s0[60]}), .c ({signal_1346, signal_1039}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_830 ( .s (rst), .b ({signal_1347, signal_1102}), .a ({Key_s1[61], Key_s0[61]}), .c ({signal_1349, signal_1038}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_831 ( .s (rst), .b ({signal_1350, signal_1101}), .a ({Key_s1[62], Key_s0[62]}), .c ({signal_1352, signal_1037}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_832 ( .s (rst), .b ({signal_1353, signal_1100}), .a ({Key_s1[63], Key_s0[63]}), .c ({signal_1355, signal_1036}) ) ;
    MUX2_X1 cell_961 ( .S (rst), .A (signal_1029), .B (1'b1), .Z (signal_1035) ) ;
    MUX2_X1 cell_962 ( .S (rst), .A (signal_1028), .B (1'b0), .Z (signal_1034) ) ;
    MUX2_X1 cell_963 ( .S (rst), .A (signal_1027), .B (1'b0), .Z (signal_1033) ) ;
    MUX2_X1 cell_964 ( .S (rst), .A (signal_1026), .B (1'b0), .Z (signal_1032) ) ;
    MUX2_X1 cell_965 ( .S (rst), .A (signal_1025), .B (1'b0), .Z (signal_1031) ) ;
    MUX2_X1 cell_966 ( .S (rst), .A (signal_1024), .B (1'b0), .Z (signal_1030) ) ;
    MUX2_X1 cell_979 ( .S (signal_940), .A (signal_759), .B (signal_939), .Z (signal_1029) ) ;
    NAND2_X1 cell_980 ( .A1 (signal_939), .A2 (signal_760), .ZN (signal_759) ) ;
    NAND2_X1 cell_981 ( .A1 (signal_761), .A2 (signal_762), .ZN (signal_760) ) ;
    NOR2_X1 cell_982 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_762) ) ;
    AND2_X1 cell_983 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_761) ) ;
    AND2_X1 cell_984 ( .A1 (signal_763), .A2 (signal_943), .ZN (signal_1027) ) ;
    NAND2_X1 cell_985 ( .A1 (signal_764), .A2 (signal_939), .ZN (signal_763) ) ;
    NOR2_X1 cell_986 ( .A1 (signal_940), .A2 (signal_765), .ZN (signal_764) ) ;
    NAND2_X1 cell_987 ( .A1 (signal_1028), .A2 (signal_766), .ZN (signal_765) ) ;
    NOR2_X1 cell_988 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_766) ) ;
    OR2_X1 cell_989 ( .A1 (signal_940), .A2 (signal_767), .ZN (signal_1024) ) ;
    NOR2_X1 cell_990 ( .A1 (signal_1025), .A2 (signal_768), .ZN (signal_767) ) ;
    NAND2_X1 cell_991 ( .A1 (signal_939), .A2 (signal_769), .ZN (signal_768) ) ;
    NOR2_X1 cell_992 ( .A1 (signal_1026), .A2 (signal_770), .ZN (signal_769) ) ;
    NAND2_X1 cell_993 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_770) ) ;
    NOR2_X1 cell_994 ( .A1 (signal_771), .A2 (signal_772), .ZN (done) ) ;
    NAND2_X1 cell_995 ( .A1 (signal_940), .A2 (signal_939), .ZN (signal_772) ) ;
    NAND2_X1 cell_996 ( .A1 (signal_773), .A2 (signal_774), .ZN (signal_771) ) ;
    NOR2_X1 cell_997 ( .A1 (signal_1025), .A2 (signal_775), .ZN (signal_774) ) ;
    INV_X1 cell_998 ( .A (signal_1028), .ZN (signal_775) ) ;
    NOR2_X1 cell_999 ( .A1 (signal_943), .A2 (signal_1026), .ZN (signal_773) ) ;

    /* cells in depth 1 */
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_0 ( .s (signal_2636), .b ({signal_1483, signal_839}), .a ({signal_2638, signal_2637}), .c ({signal_1485, signal_903}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1 ( .s (signal_2636), .b ({signal_1482, signal_838}), .a ({signal_2640, signal_2639}), .c ({signal_1487, signal_902}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2 ( .s (signal_2636), .b ({signal_1481, signal_837}), .a ({signal_2642, signal_2641}), .c ({signal_1489, signal_901}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_3 ( .s (signal_2636), .b ({signal_1480, signal_836}), .a ({signal_2644, signal_2643}), .c ({signal_1491, signal_900}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_4 ( .s (signal_2636), .b ({signal_1479, signal_835}), .a ({signal_2646, signal_2645}), .c ({signal_1493, signal_899}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_5 ( .s (signal_2636), .b ({signal_1478, signal_834}), .a ({signal_2648, signal_2647}), .c ({signal_1495, signal_898}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_6 ( .s (signal_2636), .b ({signal_1477, signal_833}), .a ({signal_2650, signal_2649}), .c ({signal_1497, signal_897}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_7 ( .s (signal_2636), .b ({signal_1476, signal_832}), .a ({signal_2652, signal_2651}), .c ({signal_1499, signal_896}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_8 ( .s (signal_2636), .b ({signal_1475, signal_831}), .a ({signal_2654, signal_2653}), .c ({signal_1501, signal_895}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_9 ( .s (signal_2636), .b ({signal_1474, signal_830}), .a ({signal_2656, signal_2655}), .c ({signal_1503, signal_894}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_10 ( .s (signal_2636), .b ({signal_1473, signal_829}), .a ({signal_2658, signal_2657}), .c ({signal_1505, signal_893}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_11 ( .s (signal_2636), .b ({signal_1472, signal_828}), .a ({signal_2660, signal_2659}), .c ({signal_1507, signal_892}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_12 ( .s (signal_2636), .b ({signal_1471, signal_827}), .a ({signal_2662, signal_2661}), .c ({signal_1509, signal_891}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_13 ( .s (signal_2636), .b ({signal_1470, signal_826}), .a ({signal_2664, signal_2663}), .c ({signal_1511, signal_890}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_14 ( .s (signal_2636), .b ({signal_1469, signal_825}), .a ({signal_2666, signal_2665}), .c ({signal_1513, signal_889}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_15 ( .s (signal_2636), .b ({signal_1468, signal_824}), .a ({signal_2668, signal_2667}), .c ({signal_1515, signal_888}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_16 ( .s (signal_2636), .b ({signal_1467, signal_823}), .a ({signal_2670, signal_2669}), .c ({signal_1517, signal_887}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_17 ( .s (signal_2636), .b ({signal_1466, signal_822}), .a ({signal_2672, signal_2671}), .c ({signal_1519, signal_886}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_18 ( .s (signal_2636), .b ({signal_1465, signal_821}), .a ({signal_2674, signal_2673}), .c ({signal_1521, signal_885}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_19 ( .s (signal_2636), .b ({signal_1464, signal_820}), .a ({signal_2676, signal_2675}), .c ({signal_1523, signal_884}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_20 ( .s (signal_2636), .b ({signal_1463, signal_819}), .a ({signal_2678, signal_2677}), .c ({signal_1525, signal_883}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_21 ( .s (signal_2636), .b ({signal_1462, signal_818}), .a ({signal_2680, signal_2679}), .c ({signal_1527, signal_882}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_22 ( .s (signal_2636), .b ({signal_1461, signal_817}), .a ({signal_2682, signal_2681}), .c ({signal_1529, signal_881}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_23 ( .s (signal_2636), .b ({signal_1460, signal_816}), .a ({signal_2684, signal_2683}), .c ({signal_1531, signal_880}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_24 ( .s (signal_2636), .b ({signal_1459, signal_815}), .a ({signal_2686, signal_2685}), .c ({signal_1533, signal_879}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_25 ( .s (signal_2636), .b ({signal_1458, signal_814}), .a ({signal_2688, signal_2687}), .c ({signal_1535, signal_878}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_26 ( .s (signal_2636), .b ({signal_1457, signal_813}), .a ({signal_2690, signal_2689}), .c ({signal_1537, signal_877}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_27 ( .s (signal_2636), .b ({signal_1456, signal_812}), .a ({signal_2692, signal_2691}), .c ({signal_1539, signal_876}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_28 ( .s (signal_2636), .b ({signal_1455, signal_811}), .a ({signal_2694, signal_2693}), .c ({signal_1541, signal_875}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_29 ( .s (signal_2636), .b ({signal_1454, signal_810}), .a ({signal_2696, signal_2695}), .c ({signal_1543, signal_874}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_30 ( .s (signal_2636), .b ({signal_1453, signal_809}), .a ({signal_2698, signal_2697}), .c ({signal_1545, signal_873}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_31 ( .s (signal_2636), .b ({signal_1452, signal_808}), .a ({signal_2700, signal_2699}), .c ({signal_1547, signal_872}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_32 ( .s (signal_2636), .b ({signal_1451, signal_807}), .a ({signal_2702, signal_2701}), .c ({signal_1549, signal_871}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_33 ( .s (signal_2636), .b ({signal_1450, signal_806}), .a ({signal_2704, signal_2703}), .c ({signal_1551, signal_870}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_34 ( .s (signal_2636), .b ({signal_1449, signal_805}), .a ({signal_2706, signal_2705}), .c ({signal_1553, signal_869}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_35 ( .s (signal_2636), .b ({signal_1448, signal_804}), .a ({signal_2708, signal_2707}), .c ({signal_1555, signal_868}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_36 ( .s (signal_2636), .b ({signal_1447, signal_803}), .a ({signal_2710, signal_2709}), .c ({signal_1557, signal_867}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_37 ( .s (signal_2636), .b ({signal_1446, signal_802}), .a ({signal_2712, signal_2711}), .c ({signal_1559, signal_866}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_38 ( .s (signal_2636), .b ({signal_1445, signal_801}), .a ({signal_2714, signal_2713}), .c ({signal_1561, signal_865}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_39 ( .s (signal_2636), .b ({signal_1444, signal_800}), .a ({signal_2716, signal_2715}), .c ({signal_1563, signal_864}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_40 ( .s (signal_2636), .b ({signal_1443, signal_799}), .a ({signal_2718, signal_2717}), .c ({signal_1565, signal_863}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_41 ( .s (signal_2636), .b ({signal_1442, signal_798}), .a ({signal_2720, signal_2719}), .c ({signal_1567, signal_862}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_42 ( .s (signal_2636), .b ({signal_1441, signal_797}), .a ({signal_2722, signal_2721}), .c ({signal_1569, signal_861}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_43 ( .s (signal_2636), .b ({signal_1440, signal_796}), .a ({signal_2724, signal_2723}), .c ({signal_1571, signal_860}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_44 ( .s (signal_2636), .b ({signal_1439, signal_795}), .a ({signal_2726, signal_2725}), .c ({signal_1573, signal_859}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_45 ( .s (signal_2636), .b ({signal_1438, signal_794}), .a ({signal_2728, signal_2727}), .c ({signal_1575, signal_858}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_46 ( .s (signal_2636), .b ({signal_1437, signal_793}), .a ({signal_2730, signal_2729}), .c ({signal_1577, signal_857}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_47 ( .s (signal_2636), .b ({signal_1436, signal_792}), .a ({signal_2732, signal_2731}), .c ({signal_1579, signal_856}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_48 ( .s (signal_2636), .b ({signal_1435, signal_791}), .a ({signal_2734, signal_2733}), .c ({signal_1581, signal_855}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_49 ( .s (signal_2636), .b ({signal_1434, signal_790}), .a ({signal_2736, signal_2735}), .c ({signal_1583, signal_854}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_50 ( .s (signal_2636), .b ({signal_1433, signal_789}), .a ({signal_2738, signal_2737}), .c ({signal_1585, signal_853}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_51 ( .s (signal_2636), .b ({signal_1432, signal_788}), .a ({signal_2740, signal_2739}), .c ({signal_1587, signal_852}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_52 ( .s (signal_2636), .b ({signal_1431, signal_787}), .a ({signal_2742, signal_2741}), .c ({signal_1589, signal_851}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_53 ( .s (signal_2636), .b ({signal_1430, signal_786}), .a ({signal_2744, signal_2743}), .c ({signal_1591, signal_850}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_54 ( .s (signal_2636), .b ({signal_1429, signal_785}), .a ({signal_2746, signal_2745}), .c ({signal_1593, signal_849}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_55 ( .s (signal_2636), .b ({signal_1428, signal_784}), .a ({signal_2748, signal_2747}), .c ({signal_1595, signal_848}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_56 ( .s (signal_2636), .b ({signal_1427, signal_783}), .a ({signal_2750, signal_2749}), .c ({signal_1597, signal_847}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_57 ( .s (signal_2636), .b ({signal_1426, signal_782}), .a ({signal_2752, signal_2751}), .c ({signal_1599, signal_846}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_58 ( .s (signal_2636), .b ({signal_1425, signal_781}), .a ({signal_2754, signal_2753}), .c ({signal_1601, signal_845}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_59 ( .s (signal_2636), .b ({signal_1424, signal_780}), .a ({signal_2756, signal_2755}), .c ({signal_1603, signal_844}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_60 ( .s (signal_2636), .b ({signal_1423, signal_779}), .a ({signal_2758, signal_2757}), .c ({signal_1605, signal_843}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_61 ( .s (signal_2636), .b ({signal_1422, signal_778}), .a ({signal_2760, signal_2759}), .c ({signal_1607, signal_842}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_62 ( .s (signal_2636), .b ({signal_1421, signal_777}), .a ({signal_2762, signal_2761}), .c ({signal_1609, signal_841}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_63 ( .s (signal_2636), .b ({signal_1420, signal_776}), .a ({signal_2764, signal_2763}), .c ({signal_1611, signal_840}) ) ;
    SkinnyTop_step2_ANF #(.low_latency(1), .pipeline(1)) cell_1000 ( .in0 ({signal_943, signal_940, signal_939, Ciphertext_s0[0], Ciphertext_s0[1], Ciphertext_s0[2], Ciphertext_s0[3], Ciphertext_s0[4], Ciphertext_s0[5], Ciphertext_s0[6], Ciphertext_s0[7], Ciphertext_s0[8], Ciphertext_s0[9], Ciphertext_s0[10], Ciphertext_s0[11], Ciphertext_s0[12], Ciphertext_s0[13], Ciphertext_s0[14], Ciphertext_s0[15], Ciphertext_s0[16], Ciphertext_s0[17], Ciphertext_s0[18], Ciphertext_s0[19], Ciphertext_s0[20], Ciphertext_s0[21], Ciphertext_s0[22], Ciphertext_s0[23], Ciphertext_s0[24], Ciphertext_s0[25], Ciphertext_s0[26], Ciphertext_s0[27], Ciphertext_s0[28], Ciphertext_s0[29], Ciphertext_s0[30], Ciphertext_s0[31], Ciphertext_s0[32], Ciphertext_s0[33], Ciphertext_s0[34], Ciphertext_s0[35], Ciphertext_s0[36], Ciphertext_s0[37], Ciphertext_s0[38], Ciphertext_s0[39], Ciphertext_s0[40], Ciphertext_s0[41], Ciphertext_s0[42], Ciphertext_s0[43], Ciphertext_s0[44], Ciphertext_s0[45], Ciphertext_s0[46], Ciphertext_s0[47], Ciphertext_s0[48], Ciphertext_s0[49], Ciphertext_s0[50], Ciphertext_s0[51], Ciphertext_s0[52], Ciphertext_s0[53], Ciphertext_s0[54], Ciphertext_s0[55], Ciphertext_s0[56], Ciphertext_s0[57], Ciphertext_s0[58], Ciphertext_s0[59], Ciphertext_s0[60], Ciphertext_s0[61], Ciphertext_s0[62], Ciphertext_s0[63], signal_1163, signal_1162, signal_1161, signal_1160, signal_1159, signal_1158, signal_1157, signal_1156, signal_1155, signal_1154, signal_1153, signal_1152, signal_1151, signal_1150, signal_1149, signal_1148, signal_1147, signal_1146, signal_1145, signal_1144, signal_1143, signal_1142, signal_1141, signal_1140, signal_1139, signal_1138, signal_1137, signal_1136, signal_1135, signal_1134, signal_1133, signal_1132, signal_1028, signal_1026, signal_1025, 1'b0}), .in1 ({1'b0, 1'b0, 1'b0, Ciphertext_s1[0], Ciphertext_s1[1], Ciphertext_s1[2], Ciphertext_s1[3], Ciphertext_s1[4], Ciphertext_s1[5], Ciphertext_s1[6], Ciphertext_s1[7], Ciphertext_s1[8], Ciphertext_s1[9], Ciphertext_s1[10], Ciphertext_s1[11], Ciphertext_s1[12], Ciphertext_s1[13], Ciphertext_s1[14], Ciphertext_s1[15], Ciphertext_s1[16], Ciphertext_s1[17], Ciphertext_s1[18], Ciphertext_s1[19], Ciphertext_s1[20], Ciphertext_s1[21], Ciphertext_s1[22], Ciphertext_s1[23], Ciphertext_s1[24], Ciphertext_s1[25], Ciphertext_s1[26], Ciphertext_s1[27], Ciphertext_s1[28], Ciphertext_s1[29], Ciphertext_s1[30], Ciphertext_s1[31], Ciphertext_s1[32], Ciphertext_s1[33], Ciphertext_s1[34], Ciphertext_s1[35], Ciphertext_s1[36], Ciphertext_s1[37], Ciphertext_s1[38], Ciphertext_s1[39], Ciphertext_s1[40], Ciphertext_s1[41], Ciphertext_s1[42], Ciphertext_s1[43], Ciphertext_s1[44], Ciphertext_s1[45], Ciphertext_s1[46], Ciphertext_s1[47], Ciphertext_s1[48], Ciphertext_s1[49], Ciphertext_s1[50], Ciphertext_s1[51], Ciphertext_s1[52], Ciphertext_s1[53], Ciphertext_s1[54], Ciphertext_s1[55], Ciphertext_s1[56], Ciphertext_s1[57], Ciphertext_s1[58], Ciphertext_s1[59], Ciphertext_s1[60], Ciphertext_s1[61], Ciphertext_s1[62], Ciphertext_s1[63], signal_1164, signal_1167, signal_1170, signal_1173, signal_1176, signal_1179, signal_1182, signal_1185, signal_1188, signal_1191, signal_1194, signal_1197, signal_1200, signal_1203, signal_1206, signal_1209, signal_1212, signal_1215, signal_1218, signal_1221, signal_1224, signal_1227, signal_1230, signal_1233, signal_1236, signal_1239, signal_1242, signal_1245, signal_1248, signal_1251, signal_1254, signal_1257, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960], Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720], Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480], Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240], Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_839, signal_838, signal_837, signal_836, signal_835, signal_834, signal_833, signal_832, signal_831, signal_830, signal_829, signal_828, signal_827, signal_826, signal_825, signal_824, signal_823, signal_822, signal_821, signal_820, signal_819, signal_818, signal_817, signal_816, signal_815, signal_814, signal_813, signal_812, signal_811, signal_810, signal_809, signal_808, signal_807, signal_806, signal_805, signal_804, signal_803, signal_802, signal_801, signal_800, signal_799, signal_798, signal_797, signal_796, signal_795, signal_794, signal_793, signal_792, signal_791, signal_790, signal_789, signal_788, signal_787, signal_786, signal_785, signal_784, signal_783, signal_782, signal_781, signal_780, signal_779, signal_778, signal_777, signal_776}), .out1 ({signal_1483, signal_1482, signal_1481, signal_1480, signal_1479, signal_1478, signal_1477, signal_1476, signal_1475, signal_1474, signal_1473, signal_1472, signal_1471, signal_1470, signal_1469, signal_1468, signal_1467, signal_1466, signal_1465, signal_1464, signal_1463, signal_1462, signal_1461, signal_1460, signal_1459, signal_1458, signal_1457, signal_1456, signal_1455, signal_1454, signal_1453, signal_1452, signal_1451, signal_1450, signal_1449, signal_1448, signal_1447, signal_1446, signal_1445, signal_1444, signal_1443, signal_1442, signal_1441, signal_1440, signal_1439, signal_1438, signal_1437, signal_1436, signal_1435, signal_1434, signal_1433, signal_1432, signal_1431, signal_1430, signal_1429, signal_1428, signal_1427, signal_1426, signal_1425, signal_1424, signal_1423, signal_1422, signal_1421, signal_1420}) ) ;
    buf_clk cell_1001 ( .C (clk), .D (rst), .Q (signal_2636) ) ;
    buf_clk cell_1002 ( .C (clk), .D (Plaintext_s0[0]), .Q (signal_2637) ) ;
    buf_clk cell_1003 ( .C (clk), .D (Plaintext_s1[0]), .Q (signal_2638) ) ;
    buf_clk cell_1004 ( .C (clk), .D (Plaintext_s0[1]), .Q (signal_2639) ) ;
    buf_clk cell_1005 ( .C (clk), .D (Plaintext_s1[1]), .Q (signal_2640) ) ;
    buf_clk cell_1006 ( .C (clk), .D (Plaintext_s0[2]), .Q (signal_2641) ) ;
    buf_clk cell_1007 ( .C (clk), .D (Plaintext_s1[2]), .Q (signal_2642) ) ;
    buf_clk cell_1008 ( .C (clk), .D (Plaintext_s0[3]), .Q (signal_2643) ) ;
    buf_clk cell_1009 ( .C (clk), .D (Plaintext_s1[3]), .Q (signal_2644) ) ;
    buf_clk cell_1010 ( .C (clk), .D (Plaintext_s0[4]), .Q (signal_2645) ) ;
    buf_clk cell_1011 ( .C (clk), .D (Plaintext_s1[4]), .Q (signal_2646) ) ;
    buf_clk cell_1012 ( .C (clk), .D (Plaintext_s0[5]), .Q (signal_2647) ) ;
    buf_clk cell_1013 ( .C (clk), .D (Plaintext_s1[5]), .Q (signal_2648) ) ;
    buf_clk cell_1014 ( .C (clk), .D (Plaintext_s0[6]), .Q (signal_2649) ) ;
    buf_clk cell_1015 ( .C (clk), .D (Plaintext_s1[6]), .Q (signal_2650) ) ;
    buf_clk cell_1016 ( .C (clk), .D (Plaintext_s0[7]), .Q (signal_2651) ) ;
    buf_clk cell_1017 ( .C (clk), .D (Plaintext_s1[7]), .Q (signal_2652) ) ;
    buf_clk cell_1018 ( .C (clk), .D (Plaintext_s0[8]), .Q (signal_2653) ) ;
    buf_clk cell_1019 ( .C (clk), .D (Plaintext_s1[8]), .Q (signal_2654) ) ;
    buf_clk cell_1020 ( .C (clk), .D (Plaintext_s0[9]), .Q (signal_2655) ) ;
    buf_clk cell_1021 ( .C (clk), .D (Plaintext_s1[9]), .Q (signal_2656) ) ;
    buf_clk cell_1022 ( .C (clk), .D (Plaintext_s0[10]), .Q (signal_2657) ) ;
    buf_clk cell_1023 ( .C (clk), .D (Plaintext_s1[10]), .Q (signal_2658) ) ;
    buf_clk cell_1024 ( .C (clk), .D (Plaintext_s0[11]), .Q (signal_2659) ) ;
    buf_clk cell_1025 ( .C (clk), .D (Plaintext_s1[11]), .Q (signal_2660) ) ;
    buf_clk cell_1026 ( .C (clk), .D (Plaintext_s0[12]), .Q (signal_2661) ) ;
    buf_clk cell_1027 ( .C (clk), .D (Plaintext_s1[12]), .Q (signal_2662) ) ;
    buf_clk cell_1028 ( .C (clk), .D (Plaintext_s0[13]), .Q (signal_2663) ) ;
    buf_clk cell_1029 ( .C (clk), .D (Plaintext_s1[13]), .Q (signal_2664) ) ;
    buf_clk cell_1030 ( .C (clk), .D (Plaintext_s0[14]), .Q (signal_2665) ) ;
    buf_clk cell_1031 ( .C (clk), .D (Plaintext_s1[14]), .Q (signal_2666) ) ;
    buf_clk cell_1032 ( .C (clk), .D (Plaintext_s0[15]), .Q (signal_2667) ) ;
    buf_clk cell_1033 ( .C (clk), .D (Plaintext_s1[15]), .Q (signal_2668) ) ;
    buf_clk cell_1034 ( .C (clk), .D (Plaintext_s0[16]), .Q (signal_2669) ) ;
    buf_clk cell_1035 ( .C (clk), .D (Plaintext_s1[16]), .Q (signal_2670) ) ;
    buf_clk cell_1036 ( .C (clk), .D (Plaintext_s0[17]), .Q (signal_2671) ) ;
    buf_clk cell_1037 ( .C (clk), .D (Plaintext_s1[17]), .Q (signal_2672) ) ;
    buf_clk cell_1038 ( .C (clk), .D (Plaintext_s0[18]), .Q (signal_2673) ) ;
    buf_clk cell_1039 ( .C (clk), .D (Plaintext_s1[18]), .Q (signal_2674) ) ;
    buf_clk cell_1040 ( .C (clk), .D (Plaintext_s0[19]), .Q (signal_2675) ) ;
    buf_clk cell_1041 ( .C (clk), .D (Plaintext_s1[19]), .Q (signal_2676) ) ;
    buf_clk cell_1042 ( .C (clk), .D (Plaintext_s0[20]), .Q (signal_2677) ) ;
    buf_clk cell_1043 ( .C (clk), .D (Plaintext_s1[20]), .Q (signal_2678) ) ;
    buf_clk cell_1044 ( .C (clk), .D (Plaintext_s0[21]), .Q (signal_2679) ) ;
    buf_clk cell_1045 ( .C (clk), .D (Plaintext_s1[21]), .Q (signal_2680) ) ;
    buf_clk cell_1046 ( .C (clk), .D (Plaintext_s0[22]), .Q (signal_2681) ) ;
    buf_clk cell_1047 ( .C (clk), .D (Plaintext_s1[22]), .Q (signal_2682) ) ;
    buf_clk cell_1048 ( .C (clk), .D (Plaintext_s0[23]), .Q (signal_2683) ) ;
    buf_clk cell_1049 ( .C (clk), .D (Plaintext_s1[23]), .Q (signal_2684) ) ;
    buf_clk cell_1050 ( .C (clk), .D (Plaintext_s0[24]), .Q (signal_2685) ) ;
    buf_clk cell_1051 ( .C (clk), .D (Plaintext_s1[24]), .Q (signal_2686) ) ;
    buf_clk cell_1052 ( .C (clk), .D (Plaintext_s0[25]), .Q (signal_2687) ) ;
    buf_clk cell_1053 ( .C (clk), .D (Plaintext_s1[25]), .Q (signal_2688) ) ;
    buf_clk cell_1054 ( .C (clk), .D (Plaintext_s0[26]), .Q (signal_2689) ) ;
    buf_clk cell_1055 ( .C (clk), .D (Plaintext_s1[26]), .Q (signal_2690) ) ;
    buf_clk cell_1056 ( .C (clk), .D (Plaintext_s0[27]), .Q (signal_2691) ) ;
    buf_clk cell_1057 ( .C (clk), .D (Plaintext_s1[27]), .Q (signal_2692) ) ;
    buf_clk cell_1058 ( .C (clk), .D (Plaintext_s0[28]), .Q (signal_2693) ) ;
    buf_clk cell_1059 ( .C (clk), .D (Plaintext_s1[28]), .Q (signal_2694) ) ;
    buf_clk cell_1060 ( .C (clk), .D (Plaintext_s0[29]), .Q (signal_2695) ) ;
    buf_clk cell_1061 ( .C (clk), .D (Plaintext_s1[29]), .Q (signal_2696) ) ;
    buf_clk cell_1062 ( .C (clk), .D (Plaintext_s0[30]), .Q (signal_2697) ) ;
    buf_clk cell_1063 ( .C (clk), .D (Plaintext_s1[30]), .Q (signal_2698) ) ;
    buf_clk cell_1064 ( .C (clk), .D (Plaintext_s0[31]), .Q (signal_2699) ) ;
    buf_clk cell_1065 ( .C (clk), .D (Plaintext_s1[31]), .Q (signal_2700) ) ;
    buf_clk cell_1066 ( .C (clk), .D (Plaintext_s0[32]), .Q (signal_2701) ) ;
    buf_clk cell_1067 ( .C (clk), .D (Plaintext_s1[32]), .Q (signal_2702) ) ;
    buf_clk cell_1068 ( .C (clk), .D (Plaintext_s0[33]), .Q (signal_2703) ) ;
    buf_clk cell_1069 ( .C (clk), .D (Plaintext_s1[33]), .Q (signal_2704) ) ;
    buf_clk cell_1070 ( .C (clk), .D (Plaintext_s0[34]), .Q (signal_2705) ) ;
    buf_clk cell_1071 ( .C (clk), .D (Plaintext_s1[34]), .Q (signal_2706) ) ;
    buf_clk cell_1072 ( .C (clk), .D (Plaintext_s0[35]), .Q (signal_2707) ) ;
    buf_clk cell_1073 ( .C (clk), .D (Plaintext_s1[35]), .Q (signal_2708) ) ;
    buf_clk cell_1074 ( .C (clk), .D (Plaintext_s0[36]), .Q (signal_2709) ) ;
    buf_clk cell_1075 ( .C (clk), .D (Plaintext_s1[36]), .Q (signal_2710) ) ;
    buf_clk cell_1076 ( .C (clk), .D (Plaintext_s0[37]), .Q (signal_2711) ) ;
    buf_clk cell_1077 ( .C (clk), .D (Plaintext_s1[37]), .Q (signal_2712) ) ;
    buf_clk cell_1078 ( .C (clk), .D (Plaintext_s0[38]), .Q (signal_2713) ) ;
    buf_clk cell_1079 ( .C (clk), .D (Plaintext_s1[38]), .Q (signal_2714) ) ;
    buf_clk cell_1080 ( .C (clk), .D (Plaintext_s0[39]), .Q (signal_2715) ) ;
    buf_clk cell_1081 ( .C (clk), .D (Plaintext_s1[39]), .Q (signal_2716) ) ;
    buf_clk cell_1082 ( .C (clk), .D (Plaintext_s0[40]), .Q (signal_2717) ) ;
    buf_clk cell_1083 ( .C (clk), .D (Plaintext_s1[40]), .Q (signal_2718) ) ;
    buf_clk cell_1084 ( .C (clk), .D (Plaintext_s0[41]), .Q (signal_2719) ) ;
    buf_clk cell_1085 ( .C (clk), .D (Plaintext_s1[41]), .Q (signal_2720) ) ;
    buf_clk cell_1086 ( .C (clk), .D (Plaintext_s0[42]), .Q (signal_2721) ) ;
    buf_clk cell_1087 ( .C (clk), .D (Plaintext_s1[42]), .Q (signal_2722) ) ;
    buf_clk cell_1088 ( .C (clk), .D (Plaintext_s0[43]), .Q (signal_2723) ) ;
    buf_clk cell_1089 ( .C (clk), .D (Plaintext_s1[43]), .Q (signal_2724) ) ;
    buf_clk cell_1090 ( .C (clk), .D (Plaintext_s0[44]), .Q (signal_2725) ) ;
    buf_clk cell_1091 ( .C (clk), .D (Plaintext_s1[44]), .Q (signal_2726) ) ;
    buf_clk cell_1092 ( .C (clk), .D (Plaintext_s0[45]), .Q (signal_2727) ) ;
    buf_clk cell_1093 ( .C (clk), .D (Plaintext_s1[45]), .Q (signal_2728) ) ;
    buf_clk cell_1094 ( .C (clk), .D (Plaintext_s0[46]), .Q (signal_2729) ) ;
    buf_clk cell_1095 ( .C (clk), .D (Plaintext_s1[46]), .Q (signal_2730) ) ;
    buf_clk cell_1096 ( .C (clk), .D (Plaintext_s0[47]), .Q (signal_2731) ) ;
    buf_clk cell_1097 ( .C (clk), .D (Plaintext_s1[47]), .Q (signal_2732) ) ;
    buf_clk cell_1098 ( .C (clk), .D (Plaintext_s0[48]), .Q (signal_2733) ) ;
    buf_clk cell_1099 ( .C (clk), .D (Plaintext_s1[48]), .Q (signal_2734) ) ;
    buf_clk cell_1100 ( .C (clk), .D (Plaintext_s0[49]), .Q (signal_2735) ) ;
    buf_clk cell_1101 ( .C (clk), .D (Plaintext_s1[49]), .Q (signal_2736) ) ;
    buf_clk cell_1102 ( .C (clk), .D (Plaintext_s0[50]), .Q (signal_2737) ) ;
    buf_clk cell_1103 ( .C (clk), .D (Plaintext_s1[50]), .Q (signal_2738) ) ;
    buf_clk cell_1104 ( .C (clk), .D (Plaintext_s0[51]), .Q (signal_2739) ) ;
    buf_clk cell_1105 ( .C (clk), .D (Plaintext_s1[51]), .Q (signal_2740) ) ;
    buf_clk cell_1106 ( .C (clk), .D (Plaintext_s0[52]), .Q (signal_2741) ) ;
    buf_clk cell_1107 ( .C (clk), .D (Plaintext_s1[52]), .Q (signal_2742) ) ;
    buf_clk cell_1108 ( .C (clk), .D (Plaintext_s0[53]), .Q (signal_2743) ) ;
    buf_clk cell_1109 ( .C (clk), .D (Plaintext_s1[53]), .Q (signal_2744) ) ;
    buf_clk cell_1110 ( .C (clk), .D (Plaintext_s0[54]), .Q (signal_2745) ) ;
    buf_clk cell_1111 ( .C (clk), .D (Plaintext_s1[54]), .Q (signal_2746) ) ;
    buf_clk cell_1112 ( .C (clk), .D (Plaintext_s0[55]), .Q (signal_2747) ) ;
    buf_clk cell_1113 ( .C (clk), .D (Plaintext_s1[55]), .Q (signal_2748) ) ;
    buf_clk cell_1114 ( .C (clk), .D (Plaintext_s0[56]), .Q (signal_2749) ) ;
    buf_clk cell_1115 ( .C (clk), .D (Plaintext_s1[56]), .Q (signal_2750) ) ;
    buf_clk cell_1116 ( .C (clk), .D (Plaintext_s0[57]), .Q (signal_2751) ) ;
    buf_clk cell_1117 ( .C (clk), .D (Plaintext_s1[57]), .Q (signal_2752) ) ;
    buf_clk cell_1118 ( .C (clk), .D (Plaintext_s0[58]), .Q (signal_2753) ) ;
    buf_clk cell_1119 ( .C (clk), .D (Plaintext_s1[58]), .Q (signal_2754) ) ;
    buf_clk cell_1120 ( .C (clk), .D (Plaintext_s0[59]), .Q (signal_2755) ) ;
    buf_clk cell_1121 ( .C (clk), .D (Plaintext_s1[59]), .Q (signal_2756) ) ;
    buf_clk cell_1122 ( .C (clk), .D (Plaintext_s0[60]), .Q (signal_2757) ) ;
    buf_clk cell_1123 ( .C (clk), .D (Plaintext_s1[60]), .Q (signal_2758) ) ;
    buf_clk cell_1124 ( .C (clk), .D (Plaintext_s0[61]), .Q (signal_2759) ) ;
    buf_clk cell_1125 ( .C (clk), .D (Plaintext_s1[61]), .Q (signal_2760) ) ;
    buf_clk cell_1126 ( .C (clk), .D (Plaintext_s0[62]), .Q (signal_2761) ) ;
    buf_clk cell_1127 ( .C (clk), .D (Plaintext_s1[62]), .Q (signal_2762) ) ;
    buf_clk cell_1128 ( .C (clk), .D (Plaintext_s0[63]), .Q (signal_2763) ) ;
    buf_clk cell_1129 ( .C (clk), .D (Plaintext_s1[63]), .Q (signal_2764) ) ;
    buf_clk cell_1130 ( .C (clk), .D (signal_1036), .Q (signal_2765) ) ;
    buf_clk cell_1131 ( .C (clk), .D (signal_1355), .Q (signal_2766) ) ;
    buf_clk cell_1132 ( .C (clk), .D (signal_1037), .Q (signal_2767) ) ;
    buf_clk cell_1133 ( .C (clk), .D (signal_1352), .Q (signal_2768) ) ;
    buf_clk cell_1134 ( .C (clk), .D (signal_1038), .Q (signal_2769) ) ;
    buf_clk cell_1135 ( .C (clk), .D (signal_1349), .Q (signal_2770) ) ;
    buf_clk cell_1136 ( .C (clk), .D (signal_1039), .Q (signal_2771) ) ;
    buf_clk cell_1137 ( .C (clk), .D (signal_1346), .Q (signal_2772) ) ;
    buf_clk cell_1138 ( .C (clk), .D (signal_1040), .Q (signal_2773) ) ;
    buf_clk cell_1139 ( .C (clk), .D (signal_1343), .Q (signal_2774) ) ;
    buf_clk cell_1140 ( .C (clk), .D (signal_1041), .Q (signal_2775) ) ;
    buf_clk cell_1141 ( .C (clk), .D (signal_1340), .Q (signal_2776) ) ;
    buf_clk cell_1142 ( .C (clk), .D (signal_1042), .Q (signal_2777) ) ;
    buf_clk cell_1143 ( .C (clk), .D (signal_1337), .Q (signal_2778) ) ;
    buf_clk cell_1144 ( .C (clk), .D (signal_1043), .Q (signal_2779) ) ;
    buf_clk cell_1145 ( .C (clk), .D (signal_1334), .Q (signal_2780) ) ;
    buf_clk cell_1146 ( .C (clk), .D (signal_1044), .Q (signal_2781) ) ;
    buf_clk cell_1147 ( .C (clk), .D (signal_1331), .Q (signal_2782) ) ;
    buf_clk cell_1148 ( .C (clk), .D (signal_1045), .Q (signal_2783) ) ;
    buf_clk cell_1149 ( .C (clk), .D (signal_1328), .Q (signal_2784) ) ;
    buf_clk cell_1150 ( .C (clk), .D (signal_1046), .Q (signal_2785) ) ;
    buf_clk cell_1151 ( .C (clk), .D (signal_1325), .Q (signal_2786) ) ;
    buf_clk cell_1152 ( .C (clk), .D (signal_1047), .Q (signal_2787) ) ;
    buf_clk cell_1153 ( .C (clk), .D (signal_1322), .Q (signal_2788) ) ;
    buf_clk cell_1154 ( .C (clk), .D (signal_1048), .Q (signal_2789) ) ;
    buf_clk cell_1155 ( .C (clk), .D (signal_1319), .Q (signal_2790) ) ;
    buf_clk cell_1156 ( .C (clk), .D (signal_1049), .Q (signal_2791) ) ;
    buf_clk cell_1157 ( .C (clk), .D (signal_1316), .Q (signal_2792) ) ;
    buf_clk cell_1158 ( .C (clk), .D (signal_1050), .Q (signal_2793) ) ;
    buf_clk cell_1159 ( .C (clk), .D (signal_1313), .Q (signal_2794) ) ;
    buf_clk cell_1160 ( .C (clk), .D (signal_1051), .Q (signal_2795) ) ;
    buf_clk cell_1161 ( .C (clk), .D (signal_1310), .Q (signal_2796) ) ;
    buf_clk cell_1162 ( .C (clk), .D (signal_1052), .Q (signal_2797) ) ;
    buf_clk cell_1163 ( .C (clk), .D (signal_1307), .Q (signal_2798) ) ;
    buf_clk cell_1164 ( .C (clk), .D (signal_1053), .Q (signal_2799) ) ;
    buf_clk cell_1165 ( .C (clk), .D (signal_1304), .Q (signal_2800) ) ;
    buf_clk cell_1166 ( .C (clk), .D (signal_1054), .Q (signal_2801) ) ;
    buf_clk cell_1167 ( .C (clk), .D (signal_1301), .Q (signal_2802) ) ;
    buf_clk cell_1168 ( .C (clk), .D (signal_1055), .Q (signal_2803) ) ;
    buf_clk cell_1169 ( .C (clk), .D (signal_1298), .Q (signal_2804) ) ;
    buf_clk cell_1170 ( .C (clk), .D (signal_1056), .Q (signal_2805) ) ;
    buf_clk cell_1171 ( .C (clk), .D (signal_1295), .Q (signal_2806) ) ;
    buf_clk cell_1172 ( .C (clk), .D (signal_1057), .Q (signal_2807) ) ;
    buf_clk cell_1173 ( .C (clk), .D (signal_1292), .Q (signal_2808) ) ;
    buf_clk cell_1174 ( .C (clk), .D (signal_1058), .Q (signal_2809) ) ;
    buf_clk cell_1175 ( .C (clk), .D (signal_1289), .Q (signal_2810) ) ;
    buf_clk cell_1176 ( .C (clk), .D (signal_1059), .Q (signal_2811) ) ;
    buf_clk cell_1177 ( .C (clk), .D (signal_1286), .Q (signal_2812) ) ;
    buf_clk cell_1178 ( .C (clk), .D (signal_1060), .Q (signal_2813) ) ;
    buf_clk cell_1179 ( .C (clk), .D (signal_1283), .Q (signal_2814) ) ;
    buf_clk cell_1180 ( .C (clk), .D (signal_1061), .Q (signal_2815) ) ;
    buf_clk cell_1181 ( .C (clk), .D (signal_1280), .Q (signal_2816) ) ;
    buf_clk cell_1182 ( .C (clk), .D (signal_1062), .Q (signal_2817) ) ;
    buf_clk cell_1183 ( .C (clk), .D (signal_1277), .Q (signal_2818) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_1063), .Q (signal_2819) ) ;
    buf_clk cell_1185 ( .C (clk), .D (signal_1274), .Q (signal_2820) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_1064), .Q (signal_2821) ) ;
    buf_clk cell_1187 ( .C (clk), .D (signal_1271), .Q (signal_2822) ) ;
    buf_clk cell_1188 ( .C (clk), .D (signal_1065), .Q (signal_2823) ) ;
    buf_clk cell_1189 ( .C (clk), .D (signal_1268), .Q (signal_2824) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_1066), .Q (signal_2825) ) ;
    buf_clk cell_1191 ( .C (clk), .D (signal_1265), .Q (signal_2826) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_1067), .Q (signal_2827) ) ;
    buf_clk cell_1193 ( .C (clk), .D (signal_1262), .Q (signal_2828) ) ;
    buf_clk cell_1194 ( .C (clk), .D (signal_1068), .Q (signal_2829) ) ;
    buf_clk cell_1195 ( .C (clk), .D (signal_1259), .Q (signal_2830) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_1069), .Q (signal_2831) ) ;
    buf_clk cell_1197 ( .C (clk), .D (signal_1256), .Q (signal_2832) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_1070), .Q (signal_2833) ) ;
    buf_clk cell_1199 ( .C (clk), .D (signal_1253), .Q (signal_2834) ) ;
    buf_clk cell_1200 ( .C (clk), .D (signal_1071), .Q (signal_2835) ) ;
    buf_clk cell_1201 ( .C (clk), .D (signal_1250), .Q (signal_2836) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_1072), .Q (signal_2837) ) ;
    buf_clk cell_1203 ( .C (clk), .D (signal_1247), .Q (signal_2838) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_1073), .Q (signal_2839) ) ;
    buf_clk cell_1205 ( .C (clk), .D (signal_1244), .Q (signal_2840) ) ;
    buf_clk cell_1206 ( .C (clk), .D (signal_1074), .Q (signal_2841) ) ;
    buf_clk cell_1207 ( .C (clk), .D (signal_1241), .Q (signal_2842) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_1075), .Q (signal_2843) ) ;
    buf_clk cell_1209 ( .C (clk), .D (signal_1238), .Q (signal_2844) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_1076), .Q (signal_2845) ) ;
    buf_clk cell_1211 ( .C (clk), .D (signal_1235), .Q (signal_2846) ) ;
    buf_clk cell_1212 ( .C (clk), .D (signal_1077), .Q (signal_2847) ) ;
    buf_clk cell_1213 ( .C (clk), .D (signal_1232), .Q (signal_2848) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_1078), .Q (signal_2849) ) ;
    buf_clk cell_1215 ( .C (clk), .D (signal_1229), .Q (signal_2850) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_1079), .Q (signal_2851) ) ;
    buf_clk cell_1217 ( .C (clk), .D (signal_1226), .Q (signal_2852) ) ;
    buf_clk cell_1218 ( .C (clk), .D (signal_1080), .Q (signal_2853) ) ;
    buf_clk cell_1219 ( .C (clk), .D (signal_1223), .Q (signal_2854) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_1081), .Q (signal_2855) ) ;
    buf_clk cell_1221 ( .C (clk), .D (signal_1220), .Q (signal_2856) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_1082), .Q (signal_2857) ) ;
    buf_clk cell_1223 ( .C (clk), .D (signal_1217), .Q (signal_2858) ) ;
    buf_clk cell_1224 ( .C (clk), .D (signal_1083), .Q (signal_2859) ) ;
    buf_clk cell_1225 ( .C (clk), .D (signal_1214), .Q (signal_2860) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_1084), .Q (signal_2861) ) ;
    buf_clk cell_1227 ( .C (clk), .D (signal_1211), .Q (signal_2862) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_1085), .Q (signal_2863) ) ;
    buf_clk cell_1229 ( .C (clk), .D (signal_1208), .Q (signal_2864) ) ;
    buf_clk cell_1230 ( .C (clk), .D (signal_1086), .Q (signal_2865) ) ;
    buf_clk cell_1231 ( .C (clk), .D (signal_1205), .Q (signal_2866) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_1087), .Q (signal_2867) ) ;
    buf_clk cell_1233 ( .C (clk), .D (signal_1202), .Q (signal_2868) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_1088), .Q (signal_2869) ) ;
    buf_clk cell_1235 ( .C (clk), .D (signal_1199), .Q (signal_2870) ) ;
    buf_clk cell_1236 ( .C (clk), .D (signal_1089), .Q (signal_2871) ) ;
    buf_clk cell_1237 ( .C (clk), .D (signal_1196), .Q (signal_2872) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_1090), .Q (signal_2873) ) ;
    buf_clk cell_1239 ( .C (clk), .D (signal_1193), .Q (signal_2874) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_1091), .Q (signal_2875) ) ;
    buf_clk cell_1241 ( .C (clk), .D (signal_1190), .Q (signal_2876) ) ;
    buf_clk cell_1242 ( .C (clk), .D (signal_1092), .Q (signal_2877) ) ;
    buf_clk cell_1243 ( .C (clk), .D (signal_1187), .Q (signal_2878) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_1093), .Q (signal_2879) ) ;
    buf_clk cell_1245 ( .C (clk), .D (signal_1184), .Q (signal_2880) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_1094), .Q (signal_2881) ) ;
    buf_clk cell_1247 ( .C (clk), .D (signal_1181), .Q (signal_2882) ) ;
    buf_clk cell_1248 ( .C (clk), .D (signal_1095), .Q (signal_2883) ) ;
    buf_clk cell_1249 ( .C (clk), .D (signal_1178), .Q (signal_2884) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_1096), .Q (signal_2885) ) ;
    buf_clk cell_1251 ( .C (clk), .D (signal_1175), .Q (signal_2886) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_1097), .Q (signal_2887) ) ;
    buf_clk cell_1253 ( .C (clk), .D (signal_1172), .Q (signal_2888) ) ;
    buf_clk cell_1254 ( .C (clk), .D (signal_1098), .Q (signal_2889) ) ;
    buf_clk cell_1255 ( .C (clk), .D (signal_1169), .Q (signal_2890) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_1099), .Q (signal_2891) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_1166), .Q (signal_2892) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_1030), .Q (signal_2893) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_1031), .Q (signal_2894) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_1032), .Q (signal_2895) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_1033), .Q (signal_2896) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_1034), .Q (signal_2897) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_1035), .Q (signal_2898) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(1)) cell_65 ( .clk (clk), .D ({signal_1611, signal_840}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_67 ( .clk (clk), .D ({signal_1609, signal_841}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_69 ( .clk (clk), .D ({signal_1607, signal_842}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_71 ( .clk (clk), .D ({signal_1605, signal_843}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_73 ( .clk (clk), .D ({signal_1603, signal_844}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_75 ( .clk (clk), .D ({signal_1601, signal_845}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_77 ( .clk (clk), .D ({signal_1599, signal_846}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_79 ( .clk (clk), .D ({signal_1597, signal_847}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_81 ( .clk (clk), .D ({signal_1595, signal_848}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_83 ( .clk (clk), .D ({signal_1593, signal_849}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_85 ( .clk (clk), .D ({signal_1591, signal_850}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_87 ( .clk (clk), .D ({signal_1589, signal_851}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_89 ( .clk (clk), .D ({signal_1587, signal_852}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_91 ( .clk (clk), .D ({signal_1585, signal_853}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_93 ( .clk (clk), .D ({signal_1583, signal_854}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_95 ( .clk (clk), .D ({signal_1581, signal_855}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_97 ( .clk (clk), .D ({signal_1579, signal_856}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_99 ( .clk (clk), .D ({signal_1577, signal_857}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_101 ( .clk (clk), .D ({signal_1575, signal_858}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_103 ( .clk (clk), .D ({signal_1573, signal_859}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_105 ( .clk (clk), .D ({signal_1571, signal_860}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_107 ( .clk (clk), .D ({signal_1569, signal_861}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_109 ( .clk (clk), .D ({signal_1567, signal_862}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_111 ( .clk (clk), .D ({signal_1565, signal_863}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_113 ( .clk (clk), .D ({signal_1563, signal_864}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_115 ( .clk (clk), .D ({signal_1561, signal_865}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_117 ( .clk (clk), .D ({signal_1559, signal_866}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_119 ( .clk (clk), .D ({signal_1557, signal_867}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_121 ( .clk (clk), .D ({signal_1555, signal_868}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_123 ( .clk (clk), .D ({signal_1553, signal_869}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_125 ( .clk (clk), .D ({signal_1551, signal_870}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_127 ( .clk (clk), .D ({signal_1549, signal_871}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_129 ( .clk (clk), .D ({signal_1547, signal_872}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_131 ( .clk (clk), .D ({signal_1545, signal_873}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_133 ( .clk (clk), .D ({signal_1543, signal_874}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_135 ( .clk (clk), .D ({signal_1541, signal_875}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_137 ( .clk (clk), .D ({signal_1539, signal_876}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_139 ( .clk (clk), .D ({signal_1537, signal_877}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_141 ( .clk (clk), .D ({signal_1535, signal_878}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_143 ( .clk (clk), .D ({signal_1533, signal_879}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_145 ( .clk (clk), .D ({signal_1531, signal_880}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_147 ( .clk (clk), .D ({signal_1529, signal_881}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_149 ( .clk (clk), .D ({signal_1527, signal_882}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_151 ( .clk (clk), .D ({signal_1525, signal_883}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_153 ( .clk (clk), .D ({signal_1523, signal_884}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_155 ( .clk (clk), .D ({signal_1521, signal_885}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_157 ( .clk (clk), .D ({signal_1519, signal_886}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_159 ( .clk (clk), .D ({signal_1517, signal_887}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_161 ( .clk (clk), .D ({signal_1515, signal_888}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_163 ( .clk (clk), .D ({signal_1513, signal_889}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_165 ( .clk (clk), .D ({signal_1511, signal_890}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_167 ( .clk (clk), .D ({signal_1509, signal_891}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_169 ( .clk (clk), .D ({signal_1507, signal_892}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_171 ( .clk (clk), .D ({signal_1505, signal_893}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_173 ( .clk (clk), .D ({signal_1503, signal_894}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_175 ( .clk (clk), .D ({signal_1501, signal_895}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_177 ( .clk (clk), .D ({signal_1499, signal_896}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_179 ( .clk (clk), .D ({signal_1497, signal_897}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_181 ( .clk (clk), .D ({signal_1495, signal_898}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_183 ( .clk (clk), .D ({signal_1493, signal_899}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_185 ( .clk (clk), .D ({signal_1491, signal_900}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_187 ( .clk (clk), .D ({signal_1489, signal_901}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_189 ( .clk (clk), .D ({signal_1487, signal_902}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_191 ( .clk (clk), .D ({signal_1485, signal_903}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_834 ( .clk (clk), .D ({signal_2766, signal_2765}), .Q ({signal_1257, signal_1132}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_836 ( .clk (clk), .D ({signal_2768, signal_2767}), .Q ({signal_1254, signal_1133}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_838 ( .clk (clk), .D ({signal_2770, signal_2769}), .Q ({signal_1251, signal_1134}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_840 ( .clk (clk), .D ({signal_2772, signal_2771}), .Q ({signal_1248, signal_1135}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_842 ( .clk (clk), .D ({signal_2774, signal_2773}), .Q ({signal_1245, signal_1136}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_844 ( .clk (clk), .D ({signal_2776, signal_2775}), .Q ({signal_1242, signal_1137}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_846 ( .clk (clk), .D ({signal_2778, signal_2777}), .Q ({signal_1239, signal_1138}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_848 ( .clk (clk), .D ({signal_2780, signal_2779}), .Q ({signal_1236, signal_1139}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_850 ( .clk (clk), .D ({signal_2782, signal_2781}), .Q ({signal_1233, signal_1140}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_852 ( .clk (clk), .D ({signal_2784, signal_2783}), .Q ({signal_1230, signal_1141}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_854 ( .clk (clk), .D ({signal_2786, signal_2785}), .Q ({signal_1227, signal_1142}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_856 ( .clk (clk), .D ({signal_2788, signal_2787}), .Q ({signal_1224, signal_1143}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_858 ( .clk (clk), .D ({signal_2790, signal_2789}), .Q ({signal_1221, signal_1144}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_860 ( .clk (clk), .D ({signal_2792, signal_2791}), .Q ({signal_1218, signal_1145}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_862 ( .clk (clk), .D ({signal_2794, signal_2793}), .Q ({signal_1215, signal_1146}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_864 ( .clk (clk), .D ({signal_2796, signal_2795}), .Q ({signal_1212, signal_1147}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_866 ( .clk (clk), .D ({signal_2798, signal_2797}), .Q ({signal_1209, signal_1148}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_868 ( .clk (clk), .D ({signal_2800, signal_2799}), .Q ({signal_1206, signal_1149}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_870 ( .clk (clk), .D ({signal_2802, signal_2801}), .Q ({signal_1203, signal_1150}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_872 ( .clk (clk), .D ({signal_2804, signal_2803}), .Q ({signal_1200, signal_1151}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_874 ( .clk (clk), .D ({signal_2806, signal_2805}), .Q ({signal_1197, signal_1152}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_876 ( .clk (clk), .D ({signal_2808, signal_2807}), .Q ({signal_1194, signal_1153}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_878 ( .clk (clk), .D ({signal_2810, signal_2809}), .Q ({signal_1191, signal_1154}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_880 ( .clk (clk), .D ({signal_2812, signal_2811}), .Q ({signal_1188, signal_1155}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_882 ( .clk (clk), .D ({signal_2814, signal_2813}), .Q ({signal_1185, signal_1156}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_884 ( .clk (clk), .D ({signal_2816, signal_2815}), .Q ({signal_1182, signal_1157}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_886 ( .clk (clk), .D ({signal_2818, signal_2817}), .Q ({signal_1179, signal_1158}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_888 ( .clk (clk), .D ({signal_2820, signal_2819}), .Q ({signal_1176, signal_1159}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_890 ( .clk (clk), .D ({signal_2822, signal_2821}), .Q ({signal_1173, signal_1160}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_892 ( .clk (clk), .D ({signal_2824, signal_2823}), .Q ({signal_1170, signal_1161}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_894 ( .clk (clk), .D ({signal_2826, signal_2825}), .Q ({signal_1167, signal_1162}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_896 ( .clk (clk), .D ({signal_2828, signal_2827}), .Q ({signal_1164, signal_1163}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_898 ( .clk (clk), .D ({signal_2830, signal_2829}), .Q ({signal_1329, signal_1108}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_900 ( .clk (clk), .D ({signal_2832, signal_2831}), .Q ({signal_1326, signal_1109}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_902 ( .clk (clk), .D ({signal_2834, signal_2833}), .Q ({signal_1323, signal_1110}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_904 ( .clk (clk), .D ({signal_2836, signal_2835}), .Q ({signal_1320, signal_1111}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_906 ( .clk (clk), .D ({signal_2838, signal_2837}), .Q ({signal_1353, signal_1100}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_908 ( .clk (clk), .D ({signal_2840, signal_2839}), .Q ({signal_1350, signal_1101}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_910 ( .clk (clk), .D ({signal_2842, signal_2841}), .Q ({signal_1347, signal_1102}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_912 ( .clk (clk), .D ({signal_2844, signal_2843}), .Q ({signal_1344, signal_1103}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_914 ( .clk (clk), .D ({signal_2846, signal_2845}), .Q ({signal_1305, signal_1116}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_916 ( .clk (clk), .D ({signal_2848, signal_2847}), .Q ({signal_1302, signal_1117}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_918 ( .clk (clk), .D ({signal_2850, signal_2849}), .Q ({signal_1299, signal_1118}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_920 ( .clk (clk), .D ({signal_2852, signal_2851}), .Q ({signal_1296, signal_1119}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_922 ( .clk (clk), .D ({signal_2854, signal_2853}), .Q ({signal_1269, signal_1128}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_924 ( .clk (clk), .D ({signal_2856, signal_2855}), .Q ({signal_1266, signal_1129}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_926 ( .clk (clk), .D ({signal_2858, signal_2857}), .Q ({signal_1263, signal_1130}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_928 ( .clk (clk), .D ({signal_2860, signal_2859}), .Q ({signal_1260, signal_1131}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_930 ( .clk (clk), .D ({signal_2862, signal_2861}), .Q ({signal_1281, signal_1124}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_932 ( .clk (clk), .D ({signal_2864, signal_2863}), .Q ({signal_1278, signal_1125}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_934 ( .clk (clk), .D ({signal_2866, signal_2865}), .Q ({signal_1275, signal_1126}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_936 ( .clk (clk), .D ({signal_2868, signal_2867}), .Q ({signal_1272, signal_1127}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_938 ( .clk (clk), .D ({signal_2870, signal_2869}), .Q ({signal_1317, signal_1112}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_940 ( .clk (clk), .D ({signal_2872, signal_2871}), .Q ({signal_1314, signal_1113}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_942 ( .clk (clk), .D ({signal_2874, signal_2873}), .Q ({signal_1311, signal_1114}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_944 ( .clk (clk), .D ({signal_2876, signal_2875}), .Q ({signal_1308, signal_1115}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_946 ( .clk (clk), .D ({signal_2878, signal_2877}), .Q ({signal_1293, signal_1120}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_948 ( .clk (clk), .D ({signal_2880, signal_2879}), .Q ({signal_1290, signal_1121}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_950 ( .clk (clk), .D ({signal_2882, signal_2881}), .Q ({signal_1287, signal_1122}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_952 ( .clk (clk), .D ({signal_2884, signal_2883}), .Q ({signal_1284, signal_1123}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_954 ( .clk (clk), .D ({signal_2886, signal_2885}), .Q ({signal_1341, signal_1104}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_956 ( .clk (clk), .D ({signal_2888, signal_2887}), .Q ({signal_1338, signal_1105}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_958 ( .clk (clk), .D ({signal_2890, signal_2889}), .Q ({signal_1335, signal_1106}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_960 ( .clk (clk), .D ({signal_2892, signal_2891}), .Q ({signal_1332, signal_1107}) ) ;
    DFF_X1 cell_968 ( .CK (clk), .D (signal_2893), .Q (signal_939), .QN () ) ;
    DFF_X1 cell_970 ( .CK (clk), .D (signal_2894), .Q (signal_940), .QN () ) ;
    DFF_X1 cell_972 ( .CK (clk), .D (signal_2895), .Q (signal_1025), .QN () ) ;
    DFF_X1 cell_974 ( .CK (clk), .D (signal_2896), .Q (signal_1026), .QN () ) ;
    DFF_X1 cell_976 ( .CK (clk), .D (signal_2897), .Q (signal_943), .QN () ) ;
    DFF_X1 cell_978 ( .CK (clk), .D (signal_2898), .Q (signal_1028), .QN () ) ;
endmodule
