/* modified netlist. Source: module SkinnyTop in file Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 26 time(s)  */

module SkinnyTop_HPC2_BDDsylvan_ClockGating_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [875:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output Synch ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_943 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2183 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2683 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2689 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2803 ;
    wire signal_2805 ;
    wire signal_2807 ;
    wire signal_2809 ;
    wire signal_2811 ;
    wire signal_2813 ;
    wire signal_2815 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2916 ;
    wire signal_2918 ;
    wire signal_2920 ;
    wire signal_2922 ;
    wire signal_2924 ;
    wire signal_2926 ;
    wire signal_2928 ;
    wire signal_2930 ;
    wire signal_2932 ;
    wire signal_2934 ;
    wire signal_2936 ;
    wire signal_2938 ;
    wire signal_2940 ;
    wire signal_2942 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3149 ;
    wire signal_3151 ;
    wire signal_3153 ;
    wire signal_3155 ;
    wire signal_3157 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3201 ;
    wire signal_3203 ;
    wire signal_3205 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3231 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3245 ;
    wire signal_3247 ;
    wire signal_3249 ;
    wire signal_3251 ;
    wire signal_3253 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_4142 ;

    /* cells in depth 0 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_769 ( .s (rst), .b ({signal_1992, signal_1163}), .a ({Key_s1[0], Key_s0[0]}), .c ({signal_1994, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_770 ( .s (rst), .b ({signal_1995, signal_1162}), .a ({Key_s1[1], Key_s0[1]}), .c ({signal_1997, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_771 ( .s (rst), .b ({signal_1998, signal_1161}), .a ({Key_s1[2], Key_s0[2]}), .c ({signal_2000, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_772 ( .s (rst), .b ({signal_2001, signal_1160}), .a ({Key_s1[3], Key_s0[3]}), .c ({signal_2003, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_773 ( .s (rst), .b ({signal_2004, signal_1159}), .a ({Key_s1[4], Key_s0[4]}), .c ({signal_2006, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_774 ( .s (rst), .b ({signal_2007, signal_1158}), .a ({Key_s1[5], Key_s0[5]}), .c ({signal_2009, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_775 ( .s (rst), .b ({signal_2010, signal_1157}), .a ({Key_s1[6], Key_s0[6]}), .c ({signal_2012, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_776 ( .s (rst), .b ({signal_2013, signal_1156}), .a ({Key_s1[7], Key_s0[7]}), .c ({signal_2015, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_777 ( .s (rst), .b ({signal_2016, signal_1155}), .a ({Key_s1[8], Key_s0[8]}), .c ({signal_2018, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_778 ( .s (rst), .b ({signal_2019, signal_1154}), .a ({Key_s1[9], Key_s0[9]}), .c ({signal_2021, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_779 ( .s (rst), .b ({signal_2022, signal_1153}), .a ({Key_s1[10], Key_s0[10]}), .c ({signal_2024, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_780 ( .s (rst), .b ({signal_2025, signal_1152}), .a ({Key_s1[11], Key_s0[11]}), .c ({signal_2027, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_781 ( .s (rst), .b ({signal_2028, signal_1151}), .a ({Key_s1[12], Key_s0[12]}), .c ({signal_2030, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_782 ( .s (rst), .b ({signal_2031, signal_1150}), .a ({Key_s1[13], Key_s0[13]}), .c ({signal_2033, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_783 ( .s (rst), .b ({signal_2034, signal_1149}), .a ({Key_s1[14], Key_s0[14]}), .c ({signal_2036, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_784 ( .s (rst), .b ({signal_2037, signal_1148}), .a ({Key_s1[15], Key_s0[15]}), .c ({signal_2039, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_785 ( .s (rst), .b ({signal_2040, signal_1147}), .a ({Key_s1[16], Key_s0[16]}), .c ({signal_2042, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_786 ( .s (rst), .b ({signal_2043, signal_1146}), .a ({Key_s1[17], Key_s0[17]}), .c ({signal_2045, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_787 ( .s (rst), .b ({signal_2046, signal_1145}), .a ({Key_s1[18], Key_s0[18]}), .c ({signal_2048, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_788 ( .s (rst), .b ({signal_2049, signal_1144}), .a ({Key_s1[19], Key_s0[19]}), .c ({signal_2051, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_789 ( .s (rst), .b ({signal_2052, signal_1143}), .a ({Key_s1[20], Key_s0[20]}), .c ({signal_2054, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_790 ( .s (rst), .b ({signal_2055, signal_1142}), .a ({Key_s1[21], Key_s0[21]}), .c ({signal_2057, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_791 ( .s (rst), .b ({signal_2058, signal_1141}), .a ({Key_s1[22], Key_s0[22]}), .c ({signal_2060, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_792 ( .s (rst), .b ({signal_2061, signal_1140}), .a ({Key_s1[23], Key_s0[23]}), .c ({signal_2063, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_793 ( .s (rst), .b ({signal_2064, signal_1139}), .a ({Key_s1[24], Key_s0[24]}), .c ({signal_2066, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_794 ( .s (rst), .b ({signal_2067, signal_1138}), .a ({Key_s1[25], Key_s0[25]}), .c ({signal_2069, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_795 ( .s (rst), .b ({signal_2070, signal_1137}), .a ({Key_s1[26], Key_s0[26]}), .c ({signal_2072, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_796 ( .s (rst), .b ({signal_2073, signal_1136}), .a ({Key_s1[27], Key_s0[27]}), .c ({signal_2075, signal_1072}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_797 ( .s (rst), .b ({signal_2076, signal_1135}), .a ({Key_s1[28], Key_s0[28]}), .c ({signal_2078, signal_1071}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_798 ( .s (rst), .b ({signal_2079, signal_1134}), .a ({Key_s1[29], Key_s0[29]}), .c ({signal_2081, signal_1070}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_799 ( .s (rst), .b ({signal_2082, signal_1133}), .a ({Key_s1[30], Key_s0[30]}), .c ({signal_2084, signal_1069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_800 ( .s (rst), .b ({signal_2085, signal_1132}), .a ({Key_s1[31], Key_s0[31]}), .c ({signal_2087, signal_1068}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_801 ( .s (rst), .b ({signal_2088, signal_1131}), .a ({Key_s1[32], Key_s0[32]}), .c ({signal_2090, signal_1067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_802 ( .s (rst), .b ({signal_2091, signal_1130}), .a ({Key_s1[33], Key_s0[33]}), .c ({signal_2093, signal_1066}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_803 ( .s (rst), .b ({signal_2094, signal_1129}), .a ({Key_s1[34], Key_s0[34]}), .c ({signal_2096, signal_1065}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_804 ( .s (rst), .b ({signal_2097, signal_1128}), .a ({Key_s1[35], Key_s0[35]}), .c ({signal_2099, signal_1064}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_805 ( .s (rst), .b ({signal_2100, signal_1127}), .a ({Key_s1[36], Key_s0[36]}), .c ({signal_2102, signal_1063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_806 ( .s (rst), .b ({signal_2103, signal_1126}), .a ({Key_s1[37], Key_s0[37]}), .c ({signal_2105, signal_1062}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_807 ( .s (rst), .b ({signal_2106, signal_1125}), .a ({Key_s1[38], Key_s0[38]}), .c ({signal_2108, signal_1061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_808 ( .s (rst), .b ({signal_2109, signal_1124}), .a ({Key_s1[39], Key_s0[39]}), .c ({signal_2111, signal_1060}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_809 ( .s (rst), .b ({signal_2112, signal_1123}), .a ({Key_s1[40], Key_s0[40]}), .c ({signal_2114, signal_1059}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_810 ( .s (rst), .b ({signal_2115, signal_1122}), .a ({Key_s1[41], Key_s0[41]}), .c ({signal_2117, signal_1058}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_811 ( .s (rst), .b ({signal_2118, signal_1121}), .a ({Key_s1[42], Key_s0[42]}), .c ({signal_2120, signal_1057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_812 ( .s (rst), .b ({signal_2121, signal_1120}), .a ({Key_s1[43], Key_s0[43]}), .c ({signal_2123, signal_1056}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_813 ( .s (rst), .b ({signal_2124, signal_1119}), .a ({Key_s1[44], Key_s0[44]}), .c ({signal_2126, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_814 ( .s (rst), .b ({signal_2127, signal_1118}), .a ({Key_s1[45], Key_s0[45]}), .c ({signal_2129, signal_1054}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_815 ( .s (rst), .b ({signal_2130, signal_1117}), .a ({Key_s1[46], Key_s0[46]}), .c ({signal_2132, signal_1053}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_816 ( .s (rst), .b ({signal_2133, signal_1116}), .a ({Key_s1[47], Key_s0[47]}), .c ({signal_2135, signal_1052}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_817 ( .s (rst), .b ({signal_2136, signal_1115}), .a ({Key_s1[48], Key_s0[48]}), .c ({signal_2138, signal_1051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_818 ( .s (rst), .b ({signal_2139, signal_1114}), .a ({Key_s1[49], Key_s0[49]}), .c ({signal_2141, signal_1050}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_819 ( .s (rst), .b ({signal_2142, signal_1113}), .a ({Key_s1[50], Key_s0[50]}), .c ({signal_2144, signal_1049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_820 ( .s (rst), .b ({signal_2145, signal_1112}), .a ({Key_s1[51], Key_s0[51]}), .c ({signal_2147, signal_1048}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_821 ( .s (rst), .b ({signal_2148, signal_1111}), .a ({Key_s1[52], Key_s0[52]}), .c ({signal_2150, signal_1047}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_822 ( .s (rst), .b ({signal_2151, signal_1110}), .a ({Key_s1[53], Key_s0[53]}), .c ({signal_2153, signal_1046}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_823 ( .s (rst), .b ({signal_2154, signal_1109}), .a ({Key_s1[54], Key_s0[54]}), .c ({signal_2156, signal_1045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_824 ( .s (rst), .b ({signal_2157, signal_1108}), .a ({Key_s1[55], Key_s0[55]}), .c ({signal_2159, signal_1044}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_825 ( .s (rst), .b ({signal_2160, signal_1107}), .a ({Key_s1[56], Key_s0[56]}), .c ({signal_2162, signal_1043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_826 ( .s (rst), .b ({signal_2163, signal_1106}), .a ({Key_s1[57], Key_s0[57]}), .c ({signal_2165, signal_1042}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_827 ( .s (rst), .b ({signal_2166, signal_1105}), .a ({Key_s1[58], Key_s0[58]}), .c ({signal_2168, signal_1041}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_828 ( .s (rst), .b ({signal_2169, signal_1104}), .a ({Key_s1[59], Key_s0[59]}), .c ({signal_2171, signal_1040}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_829 ( .s (rst), .b ({signal_2172, signal_1103}), .a ({Key_s1[60], Key_s0[60]}), .c ({signal_2174, signal_1039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_830 ( .s (rst), .b ({signal_2175, signal_1102}), .a ({Key_s1[61], Key_s0[61]}), .c ({signal_2177, signal_1038}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_831 ( .s (rst), .b ({signal_2178, signal_1101}), .a ({Key_s1[62], Key_s0[62]}), .c ({signal_2180, signal_1037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_832 ( .s (rst), .b ({signal_2181, signal_1100}), .a ({Key_s1[63], Key_s0[63]}), .c ({signal_2183, signal_1036}) ) ;
    MUX2_X1 cell_961 ( .S (rst), .A (signal_1029), .B (1'b1), .Z (signal_1035) ) ;
    MUX2_X1 cell_962 ( .S (rst), .A (signal_1028), .B (1'b0), .Z (signal_1034) ) ;
    MUX2_X1 cell_963 ( .S (rst), .A (signal_1027), .B (1'b0), .Z (signal_1033) ) ;
    MUX2_X1 cell_964 ( .S (rst), .A (signal_1026), .B (1'b0), .Z (signal_1032) ) ;
    MUX2_X1 cell_965 ( .S (rst), .A (signal_1025), .B (1'b0), .Z (signal_1031) ) ;
    MUX2_X1 cell_966 ( .S (rst), .A (signal_1024), .B (1'b0), .Z (signal_1030) ) ;
    MUX2_X1 cell_979 ( .S (signal_940), .A (signal_759), .B (signal_939), .Z (signal_1029) ) ;
    NAND2_X1 cell_980 ( .A1 (signal_939), .A2 (signal_760), .ZN (signal_759) ) ;
    NAND2_X1 cell_981 ( .A1 (signal_761), .A2 (signal_762), .ZN (signal_760) ) ;
    NOR2_X1 cell_982 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_762) ) ;
    AND2_X1 cell_983 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_761) ) ;
    AND2_X1 cell_984 ( .A1 (signal_763), .A2 (signal_943), .ZN (signal_1027) ) ;
    NAND2_X1 cell_985 ( .A1 (signal_764), .A2 (signal_939), .ZN (signal_763) ) ;
    NOR2_X1 cell_986 ( .A1 (signal_940), .A2 (signal_765), .ZN (signal_764) ) ;
    NAND2_X1 cell_987 ( .A1 (signal_1028), .A2 (signal_766), .ZN (signal_765) ) ;
    NOR2_X1 cell_988 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_766) ) ;
    OR2_X1 cell_989 ( .A1 (signal_940), .A2 (signal_767), .ZN (signal_1024) ) ;
    NOR2_X1 cell_990 ( .A1 (signal_1025), .A2 (signal_768), .ZN (signal_767) ) ;
    NAND2_X1 cell_991 ( .A1 (signal_939), .A2 (signal_769), .ZN (signal_768) ) ;
    NOR2_X1 cell_992 ( .A1 (signal_1026), .A2 (signal_770), .ZN (signal_769) ) ;
    NAND2_X1 cell_993 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_770) ) ;
    NOR2_X1 cell_994 ( .A1 (signal_771), .A2 (signal_772), .ZN (done) ) ;
    NAND2_X1 cell_995 ( .A1 (signal_940), .A2 (signal_939), .ZN (signal_772) ) ;
    NAND2_X1 cell_996 ( .A1 (signal_773), .A2 (signal_774), .ZN (signal_771) ) ;
    NOR2_X1 cell_997 ( .A1 (signal_1025), .A2 (signal_775), .ZN (signal_774) ) ;
    INV_X1 cell_998 ( .A (signal_1028), .ZN (signal_775) ) ;
    NOR2_X1 cell_999 ( .A1 (signal_943), .A2 (signal_1026), .ZN (signal_773) ) ;
    MUX2_X1 cell_1000 ( .S (1'b0), .A (1'b0), .B (1'b1), .Z (signal_1164) ) ;
    MUX2_X1 cell_1001 ( .S (1'b0), .A (1'b1), .B (1'b0), .Z (signal_1165) ) ;
    ClockGatingController #(27) cell_1892 ( .clk (clk), .rst (rst), .GatedClk (signal_4142), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1002 ( .s ({Ciphertext_s1[51], Ciphertext_s0[51]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[0]), .c ({signal_2185, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1003 ( .s ({Ciphertext_s1[51], Ciphertext_s0[51]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[1]), .c ({signal_2186, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1004 ( .s ({Ciphertext_s1[55], Ciphertext_s0[55]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[2]), .c ({signal_2188, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1005 ( .s ({Ciphertext_s1[55], Ciphertext_s0[55]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[3]), .c ({signal_2189, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1006 ( .s ({Ciphertext_s1[59], Ciphertext_s0[59]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[4]), .c ({signal_2191, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1007 ( .s ({Ciphertext_s1[59], Ciphertext_s0[59]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[5]), .c ({signal_2192, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1008 ( .s ({Ciphertext_s1[39], Ciphertext_s0[39]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[6]), .c ({signal_2194, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1009 ( .s ({Ciphertext_s1[39], Ciphertext_s0[39]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[7]), .c ({signal_2195, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1010 ( .s ({Ciphertext_s1[43], Ciphertext_s0[43]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[8]), .c ({signal_2197, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1011 ( .s ({Ciphertext_s1[43], Ciphertext_s0[43]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[9]), .c ({signal_2198, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1012 ( .s ({Ciphertext_s1[35], Ciphertext_s0[35]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[10]), .c ({signal_2200, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1013 ( .s ({Ciphertext_s1[35], Ciphertext_s0[35]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[11]), .c ({signal_2201, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1014 ( .s ({Ciphertext_s1[63], Ciphertext_s0[63]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[12]), .c ({signal_2203, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1015 ( .s ({Ciphertext_s1[63], Ciphertext_s0[63]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[13]), .c ({signal_2204, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1016 ( .s ({Ciphertext_s1[47], Ciphertext_s0[47]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[14]), .c ({signal_2206, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1017 ( .s ({Ciphertext_s1[47], Ciphertext_s0[47]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[15]), .c ({signal_2207, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1018 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[16]), .c ({signal_2209, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1019 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[17]), .c ({signal_2210, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1020 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[18]), .c ({signal_2212, signal_1184}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1021 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[19]), .c ({signal_2213, signal_1185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1022 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[20]), .c ({signal_2215, signal_1186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1023 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[21]), .c ({signal_2216, signal_1187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1024 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[22]), .c ({signal_2218, signal_1188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1025 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[23]), .c ({signal_2219, signal_1189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1026 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[24]), .c ({signal_2221, signal_1190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1027 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[25]), .c ({signal_2222, signal_1191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1028 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[26]), .c ({signal_2224, signal_1192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1029 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[27]), .c ({signal_2225, signal_1193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1030 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[28]), .c ({signal_2227, signal_1194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1031 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[29]), .c ({signal_2228, signal_1195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1032 ( .s ({Ciphertext_s1[51], Ciphertext_s0[51]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[30]), .c ({signal_2229, signal_1196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1033 ( .s ({Ciphertext_s1[51], Ciphertext_s0[51]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[31]), .c ({signal_2230, signal_1197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1034 ( .s ({Ciphertext_s1[55], Ciphertext_s0[55]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[32]), .c ({signal_2231, signal_1198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1035 ( .s ({Ciphertext_s1[55], Ciphertext_s0[55]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[33]), .c ({signal_2232, signal_1199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1036 ( .s ({Ciphertext_s1[59], Ciphertext_s0[59]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[34]), .c ({signal_2233, signal_1200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1037 ( .s ({Ciphertext_s1[59], Ciphertext_s0[59]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[35]), .c ({signal_2234, signal_1201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1064 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[36]), .c ({signal_2261, signal_1228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1065 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[37]), .c ({signal_2262, signal_1229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1066 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[38]), .c ({signal_2263, signal_1230}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1067 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[39]), .c ({signal_2264, signal_1231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1068 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[40]), .c ({signal_2265, signal_1232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1069 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[41]), .c ({signal_2266, signal_1233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .s ({Ciphertext_s1[63], Ciphertext_s0[63]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[42]), .c ({signal_2275, signal_1242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .s ({Ciphertext_s1[63], Ciphertext_s0[63]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[43]), .c ({signal_2276, signal_1243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .s ({Ciphertext_s1[47], Ciphertext_s0[47]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[44]), .c ({signal_2304, signal_1270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1107 ( .s ({Ciphertext_s1[47], Ciphertext_s0[47]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[45]), .c ({signal_2305, signal_1271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1108 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[46]), .c ({signal_2306, signal_1272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1109 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[47]), .c ({signal_2307, signal_1273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1110 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({1'b0, signal_1165}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[48]), .c ({signal_2308, signal_1274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1111 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({1'b0, signal_1164}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[49]), .c ({signal_2309, signal_1275}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1038 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2186, signal_1167}), .a ({signal_2185, signal_1166}), .clk (clk), .r (Fresh[50]), .c ({signal_2235, signal_1202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1039 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2185, signal_1166}), .a ({signal_2186, signal_1167}), .clk (clk), .r (Fresh[51]), .c ({signal_2236, signal_1203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1040 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2189, signal_1169}), .a ({signal_2188, signal_1168}), .clk (clk), .r (Fresh[52]), .c ({signal_2237, signal_1204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1041 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2188, signal_1168}), .a ({signal_2189, signal_1169}), .clk (clk), .r (Fresh[53]), .c ({signal_2238, signal_1205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1042 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2192, signal_1171}), .a ({signal_2191, signal_1170}), .clk (clk), .r (Fresh[54]), .c ({signal_2239, signal_1206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1043 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2191, signal_1170}), .a ({signal_2192, signal_1171}), .clk (clk), .r (Fresh[55]), .c ({signal_2240, signal_1207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1044 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2195, signal_1173}), .a ({signal_2194, signal_1172}), .clk (clk), .r (Fresh[56]), .c ({signal_2241, signal_1208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1045 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2194, signal_1172}), .a ({signal_2195, signal_1173}), .clk (clk), .r (Fresh[57]), .c ({signal_2242, signal_1209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1046 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2198, signal_1175}), .a ({signal_2197, signal_1174}), .clk (clk), .r (Fresh[58]), .c ({signal_2243, signal_1210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1047 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2197, signal_1174}), .a ({signal_2198, signal_1175}), .clk (clk), .r (Fresh[59]), .c ({signal_2244, signal_1211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1048 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2201, signal_1177}), .a ({signal_2200, signal_1176}), .clk (clk), .r (Fresh[60]), .c ({signal_2245, signal_1212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1049 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2200, signal_1176}), .a ({signal_2201, signal_1177}), .clk (clk), .r (Fresh[61]), .c ({signal_2246, signal_1213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1050 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2204, signal_1179}), .a ({signal_2203, signal_1178}), .clk (clk), .r (Fresh[62]), .c ({signal_2247, signal_1214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1051 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2203, signal_1178}), .a ({signal_2204, signal_1179}), .clk (clk), .r (Fresh[63]), .c ({signal_2248, signal_1215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1052 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2185, signal_1166}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[64]), .c ({signal_2249, signal_1216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1053 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2186, signal_1167}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[65]), .c ({signal_2250, signal_1217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1054 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2188, signal_1168}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[66]), .c ({signal_2251, signal_1218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1055 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2189, signal_1169}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[67]), .c ({signal_2252, signal_1219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1056 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2191, signal_1170}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[68]), .c ({signal_2253, signal_1220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1057 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2192, signal_1171}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[69]), .c ({signal_2254, signal_1221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1058 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2194, signal_1172}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[70]), .c ({signal_2255, signal_1222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1059 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2195, signal_1173}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[71]), .c ({signal_2256, signal_1223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1060 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2197, signal_1174}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[72]), .c ({signal_2257, signal_1224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1061 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2198, signal_1175}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[73]), .c ({signal_2258, signal_1225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1062 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2200, signal_1176}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[74]), .c ({signal_2259, signal_1226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1063 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2201, signal_1177}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[75]), .c ({signal_2260, signal_1227}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1070 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2203, signal_1178}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[76]), .c ({signal_2267, signal_1234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1071 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2204, signal_1179}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[77]), .c ({signal_2268, signal_1235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1072 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, 1'b1}), .a ({signal_2185, signal_1166}), .clk (clk), .r (Fresh[78]), .c ({signal_2269, signal_1236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1073 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, 1'b0}), .a ({signal_2186, signal_1167}), .clk (clk), .r (Fresh[79]), .c ({signal_2270, signal_1237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1074 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, 1'b1}), .a ({signal_2188, signal_1168}), .clk (clk), .r (Fresh[80]), .c ({signal_2271, signal_1238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, 1'b0}), .a ({signal_2189, signal_1169}), .clk (clk), .r (Fresh[81]), .c ({signal_2272, signal_1239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, 1'b1}), .a ({signal_2191, signal_1170}), .clk (clk), .r (Fresh[82]), .c ({signal_2273, signal_1240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, 1'b0}), .a ({signal_2192, signal_1171}), .clk (clk), .r (Fresh[83]), .c ({signal_2274, signal_1241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({1'b0, 1'b1}), .a ({signal_2194, signal_1172}), .clk (clk), .r (Fresh[84]), .c ({signal_2277, signal_1244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({1'b0, 1'b0}), .a ({signal_2195, signal_1173}), .clk (clk), .r (Fresh[85]), .c ({signal_2278, signal_1245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({1'b0, 1'b1}), .a ({signal_2197, signal_1174}), .clk (clk), .r (Fresh[86]), .c ({signal_2279, signal_1246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({1'b0, 1'b0}), .a ({signal_2198, signal_1175}), .clk (clk), .r (Fresh[87]), .c ({signal_2280, signal_1247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2207, signal_1181}), .a ({signal_2206, signal_1180}), .clk (clk), .r (Fresh[88]), .c ({signal_2282, signal_1248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2206, signal_1180}), .a ({signal_2207, signal_1181}), .clk (clk), .r (Fresh[89]), .c ({signal_2283, signal_1249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({1'b0, 1'b1}), .a ({signal_2200, signal_1176}), .clk (clk), .r (Fresh[90]), .c ({signal_2284, signal_1250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({1'b0, 1'b0}), .a ({signal_2201, signal_1177}), .clk (clk), .r (Fresh[91]), .c ({signal_2285, signal_1251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, 1'b1}), .a ({signal_2203, signal_1178}), .clk (clk), .r (Fresh[92]), .c ({signal_2286, signal_1252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, 1'b0}), .a ({signal_2204, signal_1179}), .clk (clk), .r (Fresh[93]), .c ({signal_2287, signal_1253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2186, signal_1167}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[94]), .c ({signal_2288, signal_1254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1091 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2185, signal_1166}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[95]), .c ({signal_2289, signal_1255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1092 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2188, signal_1168}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[96]), .c ({signal_2290, signal_1256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1093 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2189, signal_1169}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[97]), .c ({signal_2291, signal_1257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1094 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2192, signal_1171}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[98]), .c ({signal_2292, signal_1258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2191, signal_1170}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[99]), .c ({signal_2293, signal_1259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2195, signal_1173}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[100]), .c ({signal_2294, signal_1260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .s ({Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({signal_2194, signal_1172}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[101]), .c ({signal_2295, signal_1261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2197, signal_1174}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[102]), .c ({signal_2296, signal_1262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .s ({Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({signal_2198, signal_1175}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[103]), .c ({signal_2297, signal_1263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2206, signal_1180}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[104]), .c ({signal_2298, signal_1264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2207, signal_1181}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[105]), .c ({signal_2299, signal_1265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2201, signal_1177}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[106]), .c ({signal_2300, signal_1266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .s ({Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({signal_2200, signal_1176}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[107]), .c ({signal_2301, signal_1267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2204, signal_1179}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[108]), .c ({signal_2302, signal_1268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2203, signal_1178}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[109]), .c ({signal_2303, signal_1269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1112 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2230, signal_1197}), .a ({signal_2229, signal_1196}), .clk (clk), .r (Fresh[110]), .c ({signal_2310, signal_1276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1113 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2229, signal_1196}), .a ({signal_2230, signal_1197}), .clk (clk), .r (Fresh[111]), .c ({signal_2311, signal_1277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1114 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2232, signal_1199}), .a ({signal_2231, signal_1198}), .clk (clk), .r (Fresh[112]), .c ({signal_2312, signal_1278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1115 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2231, signal_1198}), .a ({signal_2232, signal_1199}), .clk (clk), .r (Fresh[113]), .c ({signal_2313, signal_1279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1116 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2234, signal_1201}), .a ({signal_2233, signal_1200}), .clk (clk), .r (Fresh[114]), .c ({signal_2314, signal_1280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1117 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2233, signal_1200}), .a ({signal_2234, signal_1201}), .clk (clk), .r (Fresh[115]), .c ({signal_2315, signal_1281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1118 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2229, signal_1196}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[116]), .c ({signal_2316, signal_1282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1119 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2230, signal_1197}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[117]), .c ({signal_2317, signal_1283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1120 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2231, signal_1198}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[118]), .c ({signal_2318, signal_1284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1121 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2232, signal_1199}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[119]), .c ({signal_2319, signal_1285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1122 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2233, signal_1200}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[120]), .c ({signal_2320, signal_1286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1123 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2234, signal_1201}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[121]), .c ({signal_2321, signal_1287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1136 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, signal_1164}), .a ({signal_2229, signal_1196}), .clk (clk), .r (Fresh[122]), .c ({signal_2340, signal_1300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1137 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({1'b0, signal_1165}), .a ({signal_2230, signal_1197}), .clk (clk), .r (Fresh[123]), .c ({signal_2341, signal_1301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1138 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, signal_1164}), .a ({signal_2231, signal_1198}), .clk (clk), .r (Fresh[124]), .c ({signal_2342, signal_1302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({1'b0, signal_1165}), .a ({signal_2232, signal_1199}), .clk (clk), .r (Fresh[125]), .c ({signal_2343, signal_1303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, signal_1164}), .a ({signal_2233, signal_1200}), .clk (clk), .r (Fresh[126]), .c ({signal_2344, signal_1304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({1'b0, signal_1165}), .a ({signal_2234, signal_1201}), .clk (clk), .r (Fresh[127]), .c ({signal_2345, signal_1305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2230, signal_1197}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[128]), .c ({signal_2367, signal_1320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .s ({Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({signal_2229, signal_1196}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[129]), .c ({signal_2368, signal_1321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2232, signal_1199}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[130]), .c ({signal_2369, signal_1322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .s ({Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({signal_2231, signal_1198}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[131]), .c ({signal_2370, signal_1323}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2234, signal_1201}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[132]), .c ({signal_2371, signal_1324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .s ({Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({signal_2233, signal_1200}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[133]), .c ({signal_2372, signal_1325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2276, signal_1243}), .a ({signal_2275, signal_1242}), .clk (clk), .r (Fresh[134]), .c ({signal_2388, signal_1340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2275, signal_1242}), .a ({signal_2276, signal_1243}), .clk (clk), .r (Fresh[135]), .c ({signal_2389, signal_1341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2275, signal_1242}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[136]), .c ({signal_2421, signal_1372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2276, signal_1243}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[137]), .c ({signal_2422, signal_1373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1228 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, signal_1164}), .a ({signal_2275, signal_1242}), .clk (clk), .r (Fresh[138]), .c ({signal_2442, signal_1392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1229 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({1'b0, signal_1165}), .a ({signal_2276, signal_1243}), .clk (clk), .r (Fresh[139]), .c ({signal_2443, signal_1393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1230 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2304, signal_1270}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[140]), .c ({signal_2444, signal_1394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1231 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({1'b0, signal_1164}), .a ({signal_2304, signal_1270}), .clk (clk), .r (Fresh[141]), .c ({signal_2445, signal_1395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1232 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2304, signal_1270}), .a ({signal_2305, signal_1271}), .clk (clk), .r (Fresh[142]), .c ({signal_2446, signal_1396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1233 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2305, signal_1271}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[143]), .c ({signal_2447, signal_1397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1234 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({1'b0, signal_1165}), .a ({signal_2305, signal_1271}), .clk (clk), .r (Fresh[144]), .c ({signal_2448, signal_1398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1235 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2305, signal_1271}), .a ({signal_2304, signal_1270}), .clk (clk), .r (Fresh[145]), .c ({signal_2449, signal_1399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1236 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2276, signal_1243}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[146]), .c ({signal_2450, signal_1400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1237 ( .s ({Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({signal_2275, signal_1242}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[147]), .c ({signal_2451, signal_1401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1238 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2305, signal_1271}), .a ({1'b0, signal_1164}), .clk (clk), .r (Fresh[148]), .c ({signal_2452, signal_1402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1239 ( .s ({Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({signal_2304, signal_1270}), .a ({1'b0, signal_1165}), .clk (clk), .r (Fresh[149]), .c ({signal_2453, signal_1403}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1124 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2235, signal_1202}), .a ({signal_2185, signal_1166}), .clk (clk), .r (Fresh[150]), .c ({signal_2323, signal_1288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1125 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2236, signal_1203}), .a ({signal_2186, signal_1167}), .clk (clk), .r (Fresh[151]), .c ({signal_2324, signal_1289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1126 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2237, signal_1204}), .a ({signal_2188, signal_1168}), .clk (clk), .r (Fresh[152]), .c ({signal_2326, signal_1290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1127 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2238, signal_1205}), .a ({signal_2189, signal_1169}), .clk (clk), .r (Fresh[153]), .c ({signal_2327, signal_1291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1128 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2239, signal_1206}), .a ({signal_2191, signal_1170}), .clk (clk), .r (Fresh[154]), .c ({signal_2329, signal_1292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1129 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2240, signal_1207}), .a ({signal_2192, signal_1171}), .clk (clk), .r (Fresh[155]), .c ({signal_2330, signal_1293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1130 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2241, signal_1208}), .a ({signal_2194, signal_1172}), .clk (clk), .r (Fresh[156]), .c ({signal_2332, signal_1294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1131 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2242, signal_1209}), .a ({signal_2195, signal_1173}), .clk (clk), .r (Fresh[157]), .c ({signal_2333, signal_1295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1132 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2243, signal_1210}), .a ({signal_2197, signal_1174}), .clk (clk), .r (Fresh[158]), .c ({signal_2335, signal_1296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1133 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2244, signal_1211}), .a ({signal_2198, signal_1175}), .clk (clk), .r (Fresh[159]), .c ({signal_2336, signal_1297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1134 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2245, signal_1212}), .a ({signal_2200, signal_1176}), .clk (clk), .r (Fresh[160]), .c ({signal_2338, signal_1298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1135 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2246, signal_1213}), .a ({signal_2201, signal_1177}), .clk (clk), .r (Fresh[161]), .c ({signal_2339, signal_1299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2247, signal_1214}), .a ({signal_2203, signal_1178}), .clk (clk), .r (Fresh[162]), .c ({signal_2347, signal_1306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2248, signal_1215}), .a ({signal_2204, signal_1179}), .clk (clk), .r (Fresh[163]), .c ({signal_2348, signal_1307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2250, signal_1217}), .a ({signal_2249, signal_1216}), .clk (clk), .r (Fresh[164]), .c ({signal_2350, signal_1308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2249, signal_1216}), .a ({signal_2250, signal_1217}), .clk (clk), .r (Fresh[165]), .c ({signal_2351, signal_1309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2252, signal_1219}), .a ({signal_2251, signal_1218}), .clk (clk), .r (Fresh[166]), .c ({signal_2353, signal_1310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2251, signal_1218}), .a ({signal_2252, signal_1219}), .clk (clk), .r (Fresh[167]), .c ({signal_2354, signal_1311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2254, signal_1221}), .a ({signal_2253, signal_1220}), .clk (clk), .r (Fresh[168]), .c ({signal_2356, signal_1312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2253, signal_1220}), .a ({signal_2254, signal_1221}), .clk (clk), .r (Fresh[169]), .c ({signal_2357, signal_1313}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2256, signal_1223}), .a ({signal_2255, signal_1222}), .clk (clk), .r (Fresh[170]), .c ({signal_2359, signal_1314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2255, signal_1222}), .a ({signal_2256, signal_1223}), .clk (clk), .r (Fresh[171]), .c ({signal_2360, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2258, signal_1225}), .a ({signal_2257, signal_1224}), .clk (clk), .r (Fresh[172]), .c ({signal_2362, signal_1316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2257, signal_1224}), .a ({signal_2258, signal_1225}), .clk (clk), .r (Fresh[173]), .c ({signal_2363, signal_1317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2260, signal_1227}), .a ({signal_2259, signal_1226}), .clk (clk), .r (Fresh[174]), .c ({signal_2365, signal_1318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2259, signal_1226}), .a ({signal_2260, signal_1227}), .clk (clk), .r (Fresh[175]), .c ({signal_2366, signal_1319}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2268, signal_1235}), .a ({signal_2267, signal_1234}), .clk (clk), .r (Fresh[176]), .c ({signal_2374, signal_1326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2267, signal_1234}), .a ({signal_2268, signal_1235}), .clk (clk), .r (Fresh[177]), .c ({signal_2375, signal_1327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({1'b0, 1'b0}), .a ({signal_2249, signal_1216}), .clk (clk), .r (Fresh[178]), .c ({signal_2376, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2236, signal_1203}), .a ({signal_2269, signal_1236}), .clk (clk), .r (Fresh[179]), .c ({signal_2377, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({1'b0, 1'b1}), .a ({signal_2250, signal_1217}), .clk (clk), .r (Fresh[180]), .c ({signal_2378, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2235, signal_1202}), .a ({signal_2270, signal_1237}), .clk (clk), .r (Fresh[181]), .c ({signal_2379, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({1'b0, 1'b0}), .a ({signal_2251, signal_1218}), .clk (clk), .r (Fresh[182]), .c ({signal_2380, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2238, signal_1205}), .a ({signal_2271, signal_1238}), .clk (clk), .r (Fresh[183]), .c ({signal_2381, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({1'b0, 1'b1}), .a ({signal_2252, signal_1219}), .clk (clk), .r (Fresh[184]), .c ({signal_2382, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2237, signal_1204}), .a ({signal_2272, signal_1239}), .clk (clk), .r (Fresh[185]), .c ({signal_2383, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({1'b0, 1'b0}), .a ({signal_2253, signal_1220}), .clk (clk), .r (Fresh[186]), .c ({signal_2384, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2240, signal_1207}), .a ({signal_2273, signal_1240}), .clk (clk), .r (Fresh[187]), .c ({signal_2385, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({1'b0, 1'b1}), .a ({signal_2254, signal_1221}), .clk (clk), .r (Fresh[188]), .c ({signal_2386, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2239, signal_1206}), .a ({signal_2274, signal_1241}), .clk (clk), .r (Fresh[189]), .c ({signal_2387, signal_1339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({1'b0, 1'b0}), .a ({signal_2255, signal_1222}), .clk (clk), .r (Fresh[190]), .c ({signal_2390, signal_1342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2242, signal_1209}), .a ({signal_2277, signal_1244}), .clk (clk), .r (Fresh[191]), .c ({signal_2391, signal_1343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({1'b0, 1'b1}), .a ({signal_2256, signal_1223}), .clk (clk), .r (Fresh[192]), .c ({signal_2392, signal_1344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2241, signal_1208}), .a ({signal_2278, signal_1245}), .clk (clk), .r (Fresh[193]), .c ({signal_2393, signal_1345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({1'b0, 1'b0}), .a ({signal_2257, signal_1224}), .clk (clk), .r (Fresh[194]), .c ({signal_2394, signal_1346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2244, signal_1211}), .a ({signal_2279, signal_1246}), .clk (clk), .r (Fresh[195]), .c ({signal_2395, signal_1347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({1'b0, 1'b1}), .a ({signal_2258, signal_1225}), .clk (clk), .r (Fresh[196]), .c ({signal_2396, signal_1348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2243, signal_1210}), .a ({signal_2280, signal_1247}), .clk (clk), .r (Fresh[197]), .c ({signal_2397, signal_1349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2282, signal_1248}), .a ({signal_2206, signal_1180}), .clk (clk), .r (Fresh[198]), .c ({signal_2399, signal_1350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2283, signal_1249}), .a ({signal_2207, signal_1181}), .clk (clk), .r (Fresh[199]), .c ({signal_2400, signal_1351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({1'b0, 1'b0}), .a ({signal_2259, signal_1226}), .clk (clk), .r (Fresh[200]), .c ({signal_2401, signal_1352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2246, signal_1213}), .a ({signal_2284, signal_1250}), .clk (clk), .r (Fresh[201]), .c ({signal_2402, signal_1353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({1'b0, 1'b1}), .a ({signal_2260, signal_1227}), .clk (clk), .r (Fresh[202]), .c ({signal_2403, signal_1354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2245, signal_1212}), .a ({signal_2285, signal_1251}), .clk (clk), .r (Fresh[203]), .c ({signal_2404, signal_1355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({1'b0, 1'b0}), .a ({signal_2267, signal_1234}), .clk (clk), .r (Fresh[204]), .c ({signal_2405, signal_1356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2248, signal_1215}), .a ({signal_2286, signal_1252}), .clk (clk), .r (Fresh[205]), .c ({signal_2406, signal_1357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({1'b0, 1'b1}), .a ({signal_2268, signal_1235}), .clk (clk), .r (Fresh[206]), .c ({signal_2407, signal_1358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2247, signal_1214}), .a ({signal_2287, signal_1253}), .clk (clk), .r (Fresh[207]), .c ({signal_2408, signal_1359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2288, signal_1254}), .a ({signal_2209, signal_1182}), .clk (clk), .r (Fresh[208]), .c ({signal_2409, signal_1360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2289, signal_1255}), .a ({signal_2209, signal_1182}), .clk (clk), .r (Fresh[209]), .c ({signal_2410, signal_1361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2289, signal_1255}), .a ({signal_2210, signal_1183}), .clk (clk), .r (Fresh[210]), .c ({signal_2411, signal_1362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2288, signal_1254}), .a ({signal_2210, signal_1183}), .clk (clk), .r (Fresh[211]), .c ({signal_2412, signal_1363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2290, signal_1256}), .a ({signal_2212, signal_1184}), .clk (clk), .r (Fresh[212]), .c ({signal_2413, signal_1364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2291, signal_1257}), .a ({signal_2212, signal_1184}), .clk (clk), .r (Fresh[213]), .c ({signal_2414, signal_1365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2291, signal_1257}), .a ({signal_2213, signal_1185}), .clk (clk), .r (Fresh[214]), .c ({signal_2415, signal_1366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2290, signal_1256}), .a ({signal_2213, signal_1185}), .clk (clk), .r (Fresh[215]), .c ({signal_2416, signal_1367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2292, signal_1258}), .a ({signal_2215, signal_1186}), .clk (clk), .r (Fresh[216]), .c ({signal_2417, signal_1368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2293, signal_1259}), .a ({signal_2215, signal_1186}), .clk (clk), .r (Fresh[217]), .c ({signal_2418, signal_1369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2293, signal_1259}), .a ({signal_2216, signal_1187}), .clk (clk), .r (Fresh[218]), .c ({signal_2419, signal_1370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2292, signal_1258}), .a ({signal_2216, signal_1187}), .clk (clk), .r (Fresh[219]), .c ({signal_2420, signal_1371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2294, signal_1260}), .a ({signal_2218, signal_1188}), .clk (clk), .r (Fresh[220]), .c ({signal_2423, signal_1374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2295, signal_1261}), .a ({signal_2218, signal_1188}), .clk (clk), .r (Fresh[221]), .c ({signal_2424, signal_1375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2295, signal_1261}), .a ({signal_2219, signal_1189}), .clk (clk), .r (Fresh[222]), .c ({signal_2425, signal_1376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .s ({Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({signal_2294, signal_1260}), .a ({signal_2219, signal_1189}), .clk (clk), .r (Fresh[223]), .c ({signal_2426, signal_1377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2296, signal_1262}), .a ({signal_2221, signal_1190}), .clk (clk), .r (Fresh[224]), .c ({signal_2427, signal_1378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2297, signal_1263}), .a ({signal_2221, signal_1190}), .clk (clk), .r (Fresh[225]), .c ({signal_2428, signal_1379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2297, signal_1263}), .a ({signal_2222, signal_1191}), .clk (clk), .r (Fresh[226]), .c ({signal_2429, signal_1380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .s ({Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({signal_2296, signal_1262}), .a ({signal_2222, signal_1191}), .clk (clk), .r (Fresh[227]), .c ({signal_2430, signal_1381}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2299, signal_1265}), .a ({signal_2298, signal_1264}), .clk (clk), .r (Fresh[228]), .c ({signal_2432, signal_1382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2298, signal_1264}), .a ({signal_2299, signal_1265}), .clk (clk), .r (Fresh[229]), .c ({signal_2433, signal_1383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2300, signal_1266}), .a ({signal_2224, signal_1192}), .clk (clk), .r (Fresh[230]), .c ({signal_2434, signal_1384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2301, signal_1267}), .a ({signal_2224, signal_1192}), .clk (clk), .r (Fresh[231]), .c ({signal_2435, signal_1385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2301, signal_1267}), .a ({signal_2225, signal_1193}), .clk (clk), .r (Fresh[232]), .c ({signal_2436, signal_1386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .s ({Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({signal_2300, signal_1266}), .a ({signal_2225, signal_1193}), .clk (clk), .r (Fresh[233]), .c ({signal_2437, signal_1387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1224 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2302, signal_1268}), .a ({signal_2227, signal_1194}), .clk (clk), .r (Fresh[234]), .c ({signal_2438, signal_1388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1225 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2303, signal_1269}), .a ({signal_2227, signal_1194}), .clk (clk), .r (Fresh[235]), .c ({signal_2439, signal_1389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1226 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2303, signal_1269}), .a ({signal_2228, signal_1195}), .clk (clk), .r (Fresh[236]), .c ({signal_2440, signal_1390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1227 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2302, signal_1268}), .a ({signal_2228, signal_1195}), .clk (clk), .r (Fresh[237]), .c ({signal_2441, signal_1391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1240 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2310, signal_1276}), .a ({signal_2229, signal_1196}), .clk (clk), .r (Fresh[238]), .c ({signal_2454, signal_1404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1241 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2311, signal_1277}), .a ({signal_2230, signal_1197}), .clk (clk), .r (Fresh[239]), .c ({signal_2455, signal_1405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1242 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2312, signal_1278}), .a ({signal_2231, signal_1198}), .clk (clk), .r (Fresh[240]), .c ({signal_2456, signal_1406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1243 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2313, signal_1279}), .a ({signal_2232, signal_1199}), .clk (clk), .r (Fresh[241]), .c ({signal_2457, signal_1407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1244 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2314, signal_1280}), .a ({signal_2233, signal_1200}), .clk (clk), .r (Fresh[242]), .c ({signal_2458, signal_1408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1245 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2315, signal_1281}), .a ({signal_2234, signal_1201}), .clk (clk), .r (Fresh[243]), .c ({signal_2459, signal_1409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1246 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2317, signal_1283}), .a ({signal_2316, signal_1282}), .clk (clk), .r (Fresh[244]), .c ({signal_2460, signal_1410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1247 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2316, signal_1282}), .a ({signal_2317, signal_1283}), .clk (clk), .r (Fresh[245]), .c ({signal_2461, signal_1411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1248 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2319, signal_1285}), .a ({signal_2318, signal_1284}), .clk (clk), .r (Fresh[246]), .c ({signal_2462, signal_1412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1249 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2318, signal_1284}), .a ({signal_2319, signal_1285}), .clk (clk), .r (Fresh[247]), .c ({signal_2463, signal_1413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1250 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2321, signal_1287}), .a ({signal_2320, signal_1286}), .clk (clk), .r (Fresh[248]), .c ({signal_2464, signal_1414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1251 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2320, signal_1286}), .a ({signal_2321, signal_1287}), .clk (clk), .r (Fresh[249]), .c ({signal_2465, signal_1415}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1264 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({1'b0, signal_1165}), .a ({signal_2316, signal_1282}), .clk (clk), .r (Fresh[250]), .c ({signal_2482, signal_1428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1265 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2311, signal_1277}), .a ({signal_2340, signal_1300}), .clk (clk), .r (Fresh[251]), .c ({signal_2483, signal_1429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1266 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({1'b0, signal_1164}), .a ({signal_2317, signal_1283}), .clk (clk), .r (Fresh[252]), .c ({signal_2484, signal_1430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2310, signal_1276}), .a ({signal_2341, signal_1301}), .clk (clk), .r (Fresh[253]), .c ({signal_2485, signal_1431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({1'b0, signal_1165}), .a ({signal_2318, signal_1284}), .clk (clk), .r (Fresh[254]), .c ({signal_2486, signal_1432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2313, signal_1279}), .a ({signal_2342, signal_1302}), .clk (clk), .r (Fresh[255]), .c ({signal_2487, signal_1433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({1'b0, signal_1164}), .a ({signal_2319, signal_1285}), .clk (clk), .r (Fresh[256]), .c ({signal_2488, signal_1434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2312, signal_1278}), .a ({signal_2343, signal_1303}), .clk (clk), .r (Fresh[257]), .c ({signal_2489, signal_1435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({1'b0, signal_1165}), .a ({signal_2320, signal_1286}), .clk (clk), .r (Fresh[258]), .c ({signal_2490, signal_1436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2315, signal_1281}), .a ({signal_2344, signal_1304}), .clk (clk), .r (Fresh[259]), .c ({signal_2491, signal_1437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({1'b0, signal_1164}), .a ({signal_2321, signal_1287}), .clk (clk), .r (Fresh[260]), .c ({signal_2492, signal_1438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2314, signal_1280}), .a ({signal_2345, signal_1305}), .clk (clk), .r (Fresh[261]), .c ({signal_2493, signal_1439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2367, signal_1320}), .a ({signal_2261, signal_1228}), .clk (clk), .r (Fresh[262]), .c ({signal_2508, signal_1454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2368, signal_1321}), .a ({signal_2261, signal_1228}), .clk (clk), .r (Fresh[263]), .c ({signal_2509, signal_1455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2368, signal_1321}), .a ({signal_2262, signal_1229}), .clk (clk), .r (Fresh[264]), .c ({signal_2510, signal_1456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .s ({Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({signal_2367, signal_1320}), .a ({signal_2262, signal_1229}), .clk (clk), .r (Fresh[265]), .c ({signal_2511, signal_1457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2369, signal_1322}), .a ({signal_2263, signal_1230}), .clk (clk), .r (Fresh[266]), .c ({signal_2512, signal_1458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2370, signal_1323}), .a ({signal_2263, signal_1230}), .clk (clk), .r (Fresh[267]), .c ({signal_2513, signal_1459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2370, signal_1323}), .a ({signal_2264, signal_1231}), .clk (clk), .r (Fresh[268]), .c ({signal_2514, signal_1460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .s ({Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({signal_2369, signal_1322}), .a ({signal_2264, signal_1231}), .clk (clk), .r (Fresh[269]), .c ({signal_2515, signal_1461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2371, signal_1324}), .a ({signal_2265, signal_1232}), .clk (clk), .r (Fresh[270]), .c ({signal_2516, signal_1462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1299 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2372, signal_1325}), .a ({signal_2265, signal_1232}), .clk (clk), .r (Fresh[271]), .c ({signal_2517, signal_1463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1300 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2372, signal_1325}), .a ({signal_2266, signal_1233}), .clk (clk), .r (Fresh[272]), .c ({signal_2518, signal_1464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1301 ( .s ({Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({signal_2371, signal_1324}), .a ({signal_2266, signal_1233}), .clk (clk), .r (Fresh[273]), .c ({signal_2519, signal_1465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1310 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2388, signal_1340}), .a ({signal_2275, signal_1242}), .clk (clk), .r (Fresh[274]), .c ({signal_2528, signal_1474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1311 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2389, signal_1341}), .a ({signal_2276, signal_1243}), .clk (clk), .r (Fresh[275]), .c ({signal_2529, signal_1475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2422, signal_1373}), .a ({signal_2421, signal_1372}), .clk (clk), .r (Fresh[276]), .c ({signal_2546, signal_1492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2421, signal_1372}), .a ({signal_2422, signal_1373}), .clk (clk), .r (Fresh[277]), .c ({signal_2547, signal_1493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1340 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({1'b0, signal_1165}), .a ({signal_2421, signal_1372}), .clk (clk), .r (Fresh[278]), .c ({signal_2558, signal_1504}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1341 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2389, signal_1341}), .a ({signal_2442, signal_1392}), .clk (clk), .r (Fresh[279]), .c ({signal_2559, signal_1505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1342 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({1'b0, signal_1164}), .a ({signal_2422, signal_1373}), .clk (clk), .r (Fresh[280]), .c ({signal_2560, signal_1506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1343 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2388, signal_1340}), .a ({signal_2443, signal_1393}), .clk (clk), .r (Fresh[281]), .c ({signal_2561, signal_1507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1344 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({1'b0, signal_1165}), .a ({signal_2444, signal_1394}), .clk (clk), .r (Fresh[282]), .c ({signal_2562, signal_1508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1345 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2446, signal_1396}), .a ({signal_2445, signal_1395}), .clk (clk), .r (Fresh[283]), .c ({signal_2563, signal_1509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1346 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({1'b0, signal_1164}), .a ({signal_2447, signal_1397}), .clk (clk), .r (Fresh[284]), .c ({signal_2564, signal_1510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1347 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2449, signal_1399}), .a ({signal_2448, signal_1398}), .clk (clk), .r (Fresh[285]), .c ({signal_2565, signal_1511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1348 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2450, signal_1400}), .a ({signal_2306, signal_1272}), .clk (clk), .r (Fresh[286]), .c ({signal_2566, signal_1512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1349 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2451, signal_1401}), .a ({signal_2306, signal_1272}), .clk (clk), .r (Fresh[287]), .c ({signal_2567, signal_1513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1350 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2451, signal_1401}), .a ({signal_2307, signal_1273}), .clk (clk), .r (Fresh[288]), .c ({signal_2568, signal_1514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1351 ( .s ({Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({signal_2450, signal_1400}), .a ({signal_2307, signal_1273}), .clk (clk), .r (Fresh[289]), .c ({signal_2569, signal_1515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1352 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2452, signal_1402}), .a ({signal_2308, signal_1274}), .clk (clk), .r (Fresh[290]), .c ({signal_2570, signal_1516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1353 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2453, signal_1403}), .a ({signal_2308, signal_1274}), .clk (clk), .r (Fresh[291]), .c ({signal_2571, signal_1517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1354 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2453, signal_1403}), .a ({signal_2309, signal_1275}), .clk (clk), .r (Fresh[292]), .c ({signal_2572, signal_1518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1355 ( .s ({Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({signal_2452, signal_1402}), .a ({signal_2309, signal_1275}), .clk (clk), .r (Fresh[293]), .c ({signal_2573, signal_1519}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_34 ( .s (rst), .b ({signal_2574, signal_805}), .a ({Plaintext_s1[34], Plaintext_s0[34]}), .c ({signal_2679, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_35 ( .s (rst), .b ({signal_2577, signal_804}), .a ({Plaintext_s1[35], Plaintext_s0[35]}), .c ({signal_2681, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_38 ( .s (rst), .b ({signal_2575, signal_801}), .a ({Plaintext_s1[38], Plaintext_s0[38]}), .c ({signal_2683, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (rst), .b ({signal_2578, signal_800}), .a ({Plaintext_s1[39], Plaintext_s0[39]}), .c ({signal_2685, signal_864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (rst), .b ({signal_2576, signal_797}), .a ({Plaintext_s1[42], Plaintext_s0[42]}), .c ({signal_2687, signal_861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (rst), .b ({signal_2579, signal_796}), .a ({Plaintext_s1[43], Plaintext_s0[43]}), .c ({signal_2689, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (rst), .b ({signal_2602, signal_793}), .a ({Plaintext_s1[46], Plaintext_s0[46]}), .c ({signal_2691, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (rst), .b ({signal_2621, signal_792}), .a ({Plaintext_s1[47], Plaintext_s0[47]}), .c ({signal_2693, signal_856}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1252 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2324, signal_1289}), .a ({signal_2323, signal_1288}), .clk (clk), .r (Fresh[294]), .c ({signal_2467, signal_1416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1253 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2323, signal_1288}), .a ({signal_2324, signal_1289}), .clk (clk), .r (Fresh[295]), .c ({signal_2468, signal_1417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1254 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2327, signal_1291}), .a ({signal_2326, signal_1290}), .clk (clk), .r (Fresh[296]), .c ({signal_2470, signal_1418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1255 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2326, signal_1290}), .a ({signal_2327, signal_1291}), .clk (clk), .r (Fresh[297]), .c ({signal_2471, signal_1419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1256 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2330, signal_1293}), .a ({signal_2329, signal_1292}), .clk (clk), .r (Fresh[298]), .c ({signal_2473, signal_1420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1257 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2329, signal_1292}), .a ({signal_2330, signal_1293}), .clk (clk), .r (Fresh[299]), .c ({signal_2474, signal_1421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1258 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2333, signal_1295}), .a ({signal_2332, signal_1294}), .clk (clk), .r (Fresh[300]), .c ({signal_2475, signal_1422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1259 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2332, signal_1294}), .a ({signal_2333, signal_1295}), .clk (clk), .r (Fresh[301]), .c ({signal_2476, signal_1423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1260 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2336, signal_1297}), .a ({signal_2335, signal_1296}), .clk (clk), .r (Fresh[302]), .c ({signal_2477, signal_1424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1261 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2335, signal_1296}), .a ({signal_2336, signal_1297}), .clk (clk), .r (Fresh[303]), .c ({signal_2478, signal_1425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1262 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2339, signal_1299}), .a ({signal_2338, signal_1298}), .clk (clk), .r (Fresh[304]), .c ({signal_2480, signal_1426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1263 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2338, signal_1298}), .a ({signal_2339, signal_1299}), .clk (clk), .r (Fresh[305]), .c ({signal_2481, signal_1427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .s ({signal_2082, signal_1133}), .b ({signal_2348, signal_1307}), .a ({signal_2347, signal_1306}), .clk (clk), .r (Fresh[306]), .c ({signal_2494, signal_1440}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .s ({signal_2082, signal_1133}), .b ({signal_2347, signal_1306}), .a ({signal_2348, signal_1307}), .clk (clk), .r (Fresh[307]), .c ({signal_2495, signal_1441}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2351, signal_1309}), .a ({signal_2350, signal_1308}), .clk (clk), .r (Fresh[308]), .c ({signal_2496, signal_1442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2350, signal_1308}), .a ({signal_2351, signal_1309}), .clk (clk), .r (Fresh[309]), .c ({signal_2497, signal_1443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2354, signal_1311}), .a ({signal_2353, signal_1310}), .clk (clk), .r (Fresh[310]), .c ({signal_2498, signal_1444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2353, signal_1310}), .a ({signal_2354, signal_1311}), .clk (clk), .r (Fresh[311]), .c ({signal_2499, signal_1445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2357, signal_1313}), .a ({signal_2356, signal_1312}), .clk (clk), .r (Fresh[312]), .c ({signal_2500, signal_1446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2356, signal_1312}), .a ({signal_2357, signal_1313}), .clk (clk), .r (Fresh[313]), .c ({signal_2501, signal_1447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2360, signal_1315}), .a ({signal_2359, signal_1314}), .clk (clk), .r (Fresh[314]), .c ({signal_2502, signal_1448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2359, signal_1314}), .a ({signal_2360, signal_1315}), .clk (clk), .r (Fresh[315]), .c ({signal_2503, signal_1449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2363, signal_1317}), .a ({signal_2362, signal_1316}), .clk (clk), .r (Fresh[316]), .c ({signal_2504, signal_1450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2362, signal_1316}), .a ({signal_2363, signal_1317}), .clk (clk), .r (Fresh[317]), .c ({signal_2505, signal_1451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2366, signal_1319}), .a ({signal_2365, signal_1318}), .clk (clk), .r (Fresh[318]), .c ({signal_2506, signal_1452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2365, signal_1318}), .a ({signal_2366, signal_1319}), .clk (clk), .r (Fresh[319]), .c ({signal_2507, signal_1453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1302 ( .s ({signal_2085, signal_1132}), .b ({signal_2375, signal_1327}), .a ({signal_2374, signal_1326}), .clk (clk), .r (Fresh[320]), .c ({signal_2520, signal_1466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1303 ( .s ({signal_2085, signal_1132}), .b ({signal_2374, signal_1326}), .a ({signal_2375, signal_1327}), .clk (clk), .r (Fresh[321]), .c ({signal_2521, signal_1467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1304 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2377, signal_1329}), .a ({signal_2376, signal_1328}), .clk (clk), .r (Fresh[322]), .c ({signal_2522, signal_1468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1305 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2379, signal_1331}), .a ({signal_2378, signal_1330}), .clk (clk), .r (Fresh[323]), .c ({signal_2523, signal_1469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1306 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2381, signal_1333}), .a ({signal_2380, signal_1332}), .clk (clk), .r (Fresh[324]), .c ({signal_2524, signal_1470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1307 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2383, signal_1335}), .a ({signal_2382, signal_1334}), .clk (clk), .r (Fresh[325]), .c ({signal_2525, signal_1471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1308 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2385, signal_1337}), .a ({signal_2384, signal_1336}), .clk (clk), .r (Fresh[326]), .c ({signal_2526, signal_1472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1309 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2387, signal_1339}), .a ({signal_2386, signal_1338}), .clk (clk), .r (Fresh[327]), .c ({signal_2527, signal_1473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1312 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2391, signal_1343}), .a ({signal_2390, signal_1342}), .clk (clk), .r (Fresh[328]), .c ({signal_2530, signal_1476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1313 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2393, signal_1345}), .a ({signal_2392, signal_1344}), .clk (clk), .r (Fresh[329]), .c ({signal_2531, signal_1477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1314 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2395, signal_1347}), .a ({signal_2394, signal_1346}), .clk (clk), .r (Fresh[330]), .c ({signal_2532, signal_1478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1315 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2397, signal_1349}), .a ({signal_2396, signal_1348}), .clk (clk), .r (Fresh[331]), .c ({signal_2533, signal_1479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1316 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2400, signal_1351}), .a ({signal_2399, signal_1350}), .clk (clk), .r (Fresh[332]), .c ({signal_2534, signal_1480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1317 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2399, signal_1350}), .a ({signal_2400, signal_1351}), .clk (clk), .r (Fresh[333]), .c ({signal_2535, signal_1481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1318 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2402, signal_1353}), .a ({signal_2401, signal_1352}), .clk (clk), .r (Fresh[334]), .c ({signal_2536, signal_1482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2404, signal_1355}), .a ({signal_2403, signal_1354}), .clk (clk), .r (Fresh[335]), .c ({signal_2537, signal_1483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2406, signal_1357}), .a ({signal_2405, signal_1356}), .clk (clk), .r (Fresh[336]), .c ({signal_2538, signal_1484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2408, signal_1359}), .a ({signal_2407, signal_1358}), .clk (clk), .r (Fresh[337]), .c ({signal_2539, signal_1485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2410, signal_1361}), .a ({signal_2409, signal_1360}), .clk (clk), .r (Fresh[338]), .c ({signal_2540, signal_1486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2412, signal_1363}), .a ({signal_2411, signal_1362}), .clk (clk), .r (Fresh[339]), .c ({signal_2541, signal_1487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2414, signal_1365}), .a ({signal_2413, signal_1364}), .clk (clk), .r (Fresh[340]), .c ({signal_2542, signal_1488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2416, signal_1367}), .a ({signal_2415, signal_1366}), .clk (clk), .r (Fresh[341]), .c ({signal_2543, signal_1489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2418, signal_1369}), .a ({signal_2417, signal_1368}), .clk (clk), .r (Fresh[342]), .c ({signal_2544, signal_1490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2420, signal_1371}), .a ({signal_2419, signal_1370}), .clk (clk), .r (Fresh[343]), .c ({signal_2545, signal_1491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2424, signal_1375}), .a ({signal_2423, signal_1374}), .clk (clk), .r (Fresh[344]), .c ({signal_2548, signal_1494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .s ({Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({signal_2426, signal_1377}), .a ({signal_2425, signal_1376}), .clk (clk), .r (Fresh[345]), .c ({signal_2549, signal_1495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2428, signal_1379}), .a ({signal_2427, signal_1378}), .clk (clk), .r (Fresh[346]), .c ({signal_2550, signal_1496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1333 ( .s ({Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({signal_2430, signal_1381}), .a ({signal_2429, signal_1380}), .clk (clk), .r (Fresh[347]), .c ({signal_2551, signal_1497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1334 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2433, signal_1383}), .a ({signal_2432, signal_1382}), .clk (clk), .r (Fresh[348]), .c ({signal_2552, signal_1498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1335 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2432, signal_1382}), .a ({signal_2433, signal_1383}), .clk (clk), .r (Fresh[349]), .c ({signal_2553, signal_1499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1336 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2435, signal_1385}), .a ({signal_2434, signal_1384}), .clk (clk), .r (Fresh[350]), .c ({signal_2554, signal_1500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1337 ( .s ({Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({signal_2437, signal_1387}), .a ({signal_2436, signal_1386}), .clk (clk), .r (Fresh[351]), .c ({signal_2555, signal_1501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1338 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2439, signal_1389}), .a ({signal_2438, signal_1388}), .clk (clk), .r (Fresh[352]), .c ({signal_2556, signal_1502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1339 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2441, signal_1391}), .a ({signal_2440, signal_1390}), .clk (clk), .r (Fresh[353]), .c ({signal_2557, signal_1503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1356 ( .s ({signal_2046, signal_1145}), .b ({signal_2455, signal_1405}), .a ({signal_2454, signal_1404}), .clk (clk), .r (Fresh[354]), .c ({signal_2574, signal_805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1357 ( .s ({signal_2058, signal_1141}), .b ({signal_2457, signal_1407}), .a ({signal_2456, signal_1406}), .clk (clk), .r (Fresh[355]), .c ({signal_2575, signal_801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1358 ( .s ({signal_2070, signal_1137}), .b ({signal_2459, signal_1409}), .a ({signal_2458, signal_1408}), .clk (clk), .r (Fresh[356]), .c ({signal_2576, signal_797}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1359 ( .s ({signal_2049, signal_1144}), .b ({signal_2461, signal_1411}), .a ({signal_2460, signal_1410}), .clk (clk), .r (Fresh[357]), .c ({signal_2577, signal_804}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1360 ( .s ({signal_2061, signal_1140}), .b ({signal_2463, signal_1413}), .a ({signal_2462, signal_1412}), .clk (clk), .r (Fresh[358]), .c ({signal_2578, signal_800}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1361 ( .s ({signal_2073, signal_1136}), .b ({signal_2465, signal_1415}), .a ({signal_2464, signal_1414}), .clk (clk), .r (Fresh[359]), .c ({signal_2579, signal_796}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1374 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2483, signal_1429}), .a ({signal_2482, signal_1428}), .clk (clk), .r (Fresh[360]), .c ({signal_2596, signal_1532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1375 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2485, signal_1431}), .a ({signal_2484, signal_1430}), .clk (clk), .r (Fresh[361]), .c ({signal_2597, signal_1533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1376 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2487, signal_1433}), .a ({signal_2486, signal_1432}), .clk (clk), .r (Fresh[362]), .c ({signal_2598, signal_1534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1377 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2489, signal_1435}), .a ({signal_2488, signal_1434}), .clk (clk), .r (Fresh[363]), .c ({signal_2599, signal_1535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1378 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2491, signal_1437}), .a ({signal_2490, signal_1436}), .clk (clk), .r (Fresh[364]), .c ({signal_2600, signal_1536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1379 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2493, signal_1439}), .a ({signal_2492, signal_1438}), .clk (clk), .r (Fresh[365]), .c ({signal_2601, signal_1537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1380 ( .s (signal_1026), .b ({signal_2495, signal_1441}), .a ({signal_2494, signal_1440}), .c ({signal_2602, signal_793}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2509, signal_1455}), .a ({signal_2508, signal_1454}), .clk (clk), .r (Fresh[366]), .c ({signal_2615, signal_1550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .s ({Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({signal_2511, signal_1457}), .a ({signal_2510, signal_1456}), .clk (clk), .r (Fresh[367]), .c ({signal_2616, signal_1551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2513, signal_1459}), .a ({signal_2512, signal_1458}), .clk (clk), .r (Fresh[368]), .c ({signal_2617, signal_1552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .s ({Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({signal_2515, signal_1461}), .a ({signal_2514, signal_1460}), .clk (clk), .r (Fresh[369]), .c ({signal_2618, signal_1553}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2517, signal_1463}), .a ({signal_2516, signal_1462}), .clk (clk), .r (Fresh[370]), .c ({signal_2619, signal_1554}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1398 ( .s ({Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({signal_2519, signal_1465}), .a ({signal_2518, signal_1464}), .clk (clk), .r (Fresh[371]), .c ({signal_2620, signal_1555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1399 ( .s (signal_1025), .b ({signal_2521, signal_1467}), .a ({signal_2520, signal_1466}), .c ({signal_2621, signal_792}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1406 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2529, signal_1475}), .a ({signal_2528, signal_1474}), .clk (clk), .r (Fresh[372]), .c ({signal_2628, signal_1562}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1407 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2528, signal_1474}), .a ({signal_2529, signal_1475}), .clk (clk), .r (Fresh[373]), .c ({signal_2629, signal_1563}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2547, signal_1493}), .a ({signal_2546, signal_1492}), .clk (clk), .r (Fresh[374]), .c ({signal_2652, signal_1586}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2546, signal_1492}), .a ({signal_2547, signal_1493}), .clk (clk), .r (Fresh[375]), .c ({signal_2653, signal_1587}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1448 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2559, signal_1505}), .a ({signal_2558, signal_1504}), .clk (clk), .r (Fresh[376]), .c ({signal_2670, signal_1604}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1449 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2561, signal_1507}), .a ({signal_2560, signal_1506}), .clk (clk), .r (Fresh[377]), .c ({signal_2671, signal_1605}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1450 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2563, signal_1509}), .a ({signal_2562, signal_1508}), .clk (clk), .r (Fresh[378]), .c ({signal_2672, signal_1606}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1451 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2565, signal_1511}), .a ({signal_2564, signal_1510}), .clk (clk), .r (Fresh[379]), .c ({signal_2673, signal_1607}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1452 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2567, signal_1513}), .a ({signal_2566, signal_1512}), .clk (clk), .r (Fresh[380]), .c ({signal_2674, signal_1608}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1453 ( .s ({Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({signal_2569, signal_1515}), .a ({signal_2568, signal_1514}), .clk (clk), .r (Fresh[381]), .c ({signal_2675, signal_1609}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1454 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2571, signal_1517}), .a ({signal_2570, signal_1516}), .clk (clk), .r (Fresh[382]), .c ({signal_2676, signal_1610}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1455 ( .s ({Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({signal_2573, signal_1519}), .a ({signal_2572, signal_1518}), .clk (clk), .r (Fresh[383]), .c ({signal_2677, signal_1611}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_32 ( .s (rst), .b ({signal_2710, signal_807}), .a ({Plaintext_s1[32], Plaintext_s0[32]}), .c ({signal_2803, signal_871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_33 ( .s (rst), .b ({signal_2729, signal_806}), .a ({Plaintext_s1[33], Plaintext_s0[33]}), .c ({signal_2805, signal_870}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_36 ( .s (rst), .b ({signal_2711, signal_803}), .a ({Plaintext_s1[36], Plaintext_s0[36]}), .c ({signal_2807, signal_867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_37 ( .s (rst), .b ({signal_2730, signal_802}), .a ({Plaintext_s1[37], Plaintext_s0[37]}), .c ({signal_2809, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (rst), .b ({signal_2712, signal_799}), .a ({Plaintext_s1[40], Plaintext_s0[40]}), .c ({signal_2811, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (rst), .b ({signal_2731, signal_798}), .a ({Plaintext_s1[41], Plaintext_s0[41]}), .c ({signal_2813, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (rst), .b ({signal_2772, signal_795}), .a ({Plaintext_s1[44], Plaintext_s0[44]}), .c ({signal_2815, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (rst), .b ({signal_2789, signal_794}), .a ({Plaintext_s1[45], Plaintext_s0[45]}), .c ({signal_2817, signal_858}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1362 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2468, signal_1417}), .a ({signal_2467, signal_1416}), .clk (clk), .r (Fresh[384]), .c ({signal_2581, signal_1520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2467, signal_1416}), .a ({signal_2468, signal_1417}), .clk (clk), .r (Fresh[385]), .c ({signal_2582, signal_1521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2471, signal_1419}), .a ({signal_2470, signal_1418}), .clk (clk), .r (Fresh[386]), .c ({signal_2584, signal_1522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2470, signal_1418}), .a ({signal_2471, signal_1419}), .clk (clk), .r (Fresh[387]), .c ({signal_2585, signal_1523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2474, signal_1421}), .a ({signal_2473, signal_1420}), .clk (clk), .r (Fresh[388]), .c ({signal_2587, signal_1524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2473, signal_1420}), .a ({signal_2474, signal_1421}), .clk (clk), .r (Fresh[389]), .c ({signal_2588, signal_1525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1368 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2476, signal_1423}), .a ({signal_2475, signal_1422}), .clk (clk), .r (Fresh[390]), .c ({signal_2589, signal_1526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1369 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2475, signal_1422}), .a ({signal_2476, signal_1423}), .clk (clk), .r (Fresh[391]), .c ({signal_2590, signal_1527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1370 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2478, signal_1425}), .a ({signal_2477, signal_1424}), .clk (clk), .r (Fresh[392]), .c ({signal_2591, signal_1528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1371 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2477, signal_1424}), .a ({signal_2478, signal_1425}), .clk (clk), .r (Fresh[393]), .c ({signal_2592, signal_1529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1372 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2481, signal_1427}), .a ({signal_2480, signal_1426}), .clk (clk), .r (Fresh[394]), .c ({signal_2594, signal_1530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1373 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2480, signal_1426}), .a ({signal_2481, signal_1427}), .clk (clk), .r (Fresh[395]), .c ({signal_2595, signal_1531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1381 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2496, signal_1442}), .a ({signal_2350, signal_1308}), .clk (clk), .r (Fresh[396]), .c ({signal_2603, signal_1538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1382 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2497, signal_1443}), .a ({signal_2351, signal_1309}), .clk (clk), .r (Fresh[397]), .c ({signal_2604, signal_1539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1383 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2498, signal_1444}), .a ({signal_2353, signal_1310}), .clk (clk), .r (Fresh[398]), .c ({signal_2605, signal_1540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2499, signal_1445}), .a ({signal_2354, signal_1311}), .clk (clk), .r (Fresh[399]), .c ({signal_2606, signal_1541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2500, signal_1446}), .a ({signal_2356, signal_1312}), .clk (clk), .r (Fresh[400]), .c ({signal_2607, signal_1542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2501, signal_1447}), .a ({signal_2357, signal_1313}), .clk (clk), .r (Fresh[401]), .c ({signal_2608, signal_1543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2502, signal_1448}), .a ({signal_2359, signal_1314}), .clk (clk), .r (Fresh[402]), .c ({signal_2609, signal_1544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2503, signal_1449}), .a ({signal_2360, signal_1315}), .clk (clk), .r (Fresh[403]), .c ({signal_2610, signal_1545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2504, signal_1450}), .a ({signal_2362, signal_1316}), .clk (clk), .r (Fresh[404]), .c ({signal_2611, signal_1546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2505, signal_1451}), .a ({signal_2363, signal_1317}), .clk (clk), .r (Fresh[405]), .c ({signal_2612, signal_1547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2506, signal_1452}), .a ({signal_2365, signal_1318}), .clk (clk), .r (Fresh[406]), .c ({signal_2613, signal_1548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2507, signal_1453}), .a ({signal_2366, signal_1319}), .clk (clk), .r (Fresh[407]), .c ({signal_2614, signal_1549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1400 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2523, signal_1469}), .a ({signal_2522, signal_1468}), .clk (clk), .r (Fresh[408]), .c ({signal_2622, signal_1556}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1401 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2522, signal_1468}), .a ({signal_2523, signal_1469}), .clk (clk), .r (Fresh[409]), .c ({signal_2623, signal_1557}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1402 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2525, signal_1471}), .a ({signal_2524, signal_1470}), .clk (clk), .r (Fresh[410]), .c ({signal_2624, signal_1558}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1403 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2524, signal_1470}), .a ({signal_2525, signal_1471}), .clk (clk), .r (Fresh[411]), .c ({signal_2625, signal_1559}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1404 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2527, signal_1473}), .a ({signal_2526, signal_1472}), .clk (clk), .r (Fresh[412]), .c ({signal_2626, signal_1560}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1405 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2526, signal_1472}), .a ({signal_2527, signal_1473}), .clk (clk), .r (Fresh[413]), .c ({signal_2627, signal_1561}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1408 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2531, signal_1477}), .a ({signal_2530, signal_1476}), .clk (clk), .r (Fresh[414]), .c ({signal_2630, signal_1564}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1409 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2530, signal_1476}), .a ({signal_2531, signal_1477}), .clk (clk), .r (Fresh[415]), .c ({signal_2631, signal_1565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1410 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2533, signal_1479}), .a ({signal_2532, signal_1478}), .clk (clk), .r (Fresh[416]), .c ({signal_2632, signal_1566}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1411 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2532, signal_1478}), .a ({signal_2533, signal_1479}), .clk (clk), .r (Fresh[417]), .c ({signal_2633, signal_1567}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1412 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2535, signal_1481}), .a ({signal_2534, signal_1480}), .clk (clk), .r (Fresh[418]), .c ({signal_2634, signal_1568}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1413 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2534, signal_1480}), .a ({signal_2535, signal_1481}), .clk (clk), .r (Fresh[419]), .c ({signal_2635, signal_1569}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1414 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2537, signal_1483}), .a ({signal_2536, signal_1482}), .clk (clk), .r (Fresh[420]), .c ({signal_2636, signal_1570}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1415 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2536, signal_1482}), .a ({signal_2537, signal_1483}), .clk (clk), .r (Fresh[421]), .c ({signal_2637, signal_1571}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .s ({signal_2076, signal_1135}), .b ({signal_2539, signal_1485}), .a ({signal_2538, signal_1484}), .clk (clk), .r (Fresh[422]), .c ({signal_2638, signal_1572}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .s ({signal_2076, signal_1135}), .b ({signal_2538, signal_1484}), .a ({signal_2539, signal_1485}), .clk (clk), .r (Fresh[423]), .c ({signal_2639, signal_1573}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2541, signal_1487}), .a ({signal_2540, signal_1486}), .clk (clk), .r (Fresh[424]), .c ({signal_2640, signal_1574}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2540, signal_1486}), .a ({signal_2541, signal_1487}), .clk (clk), .r (Fresh[425]), .c ({signal_2641, signal_1575}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2541, signal_1487}), .a ({signal_2540, signal_1486}), .clk (clk), .r (Fresh[426]), .c ({signal_2642, signal_1576}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2540, signal_1486}), .a ({signal_2541, signal_1487}), .clk (clk), .r (Fresh[427]), .c ({signal_2643, signal_1577}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2543, signal_1489}), .a ({signal_2542, signal_1488}), .clk (clk), .r (Fresh[428]), .c ({signal_2644, signal_1578}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2542, signal_1488}), .a ({signal_2543, signal_1489}), .clk (clk), .r (Fresh[429]), .c ({signal_2645, signal_1579}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2543, signal_1489}), .a ({signal_2542, signal_1488}), .clk (clk), .r (Fresh[430]), .c ({signal_2646, signal_1580}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2542, signal_1488}), .a ({signal_2543, signal_1489}), .clk (clk), .r (Fresh[431]), .c ({signal_2647, signal_1581}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2545, signal_1491}), .a ({signal_2544, signal_1490}), .clk (clk), .r (Fresh[432]), .c ({signal_2648, signal_1582}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2544, signal_1490}), .a ({signal_2545, signal_1491}), .clk (clk), .r (Fresh[433]), .c ({signal_2649, signal_1583}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2545, signal_1491}), .a ({signal_2544, signal_1490}), .clk (clk), .r (Fresh[434]), .c ({signal_2650, signal_1584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2544, signal_1490}), .a ({signal_2545, signal_1491}), .clk (clk), .r (Fresh[435]), .c ({signal_2651, signal_1585}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2549, signal_1495}), .a ({signal_2548, signal_1494}), .clk (clk), .r (Fresh[436]), .c ({signal_2654, signal_1588}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2548, signal_1494}), .a ({signal_2549, signal_1495}), .clk (clk), .r (Fresh[437]), .c ({signal_2655, signal_1589}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .s ({Ciphertext_s1[27], Ciphertext_s0[27]}), .b ({signal_2549, signal_1495}), .a ({signal_2548, signal_1494}), .clk (clk), .r (Fresh[438]), .c ({signal_2656, signal_1590}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2548, signal_1494}), .a ({signal_2549, signal_1495}), .clk (clk), .r (Fresh[439]), .c ({signal_2657, signal_1591}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2551, signal_1497}), .a ({signal_2550, signal_1496}), .clk (clk), .r (Fresh[440]), .c ({signal_2658, signal_1592}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2550, signal_1496}), .a ({signal_2551, signal_1497}), .clk (clk), .r (Fresh[441]), .c ({signal_2659, signal_1593}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .s ({Ciphertext_s1[31], Ciphertext_s0[31]}), .b ({signal_2551, signal_1497}), .a ({signal_2550, signal_1496}), .clk (clk), .r (Fresh[442]), .c ({signal_2660, signal_1594}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2550, signal_1496}), .a ({signal_2551, signal_1497}), .clk (clk), .r (Fresh[443]), .c ({signal_2661, signal_1595}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2552, signal_1498}), .a ({signal_2432, signal_1382}), .clk (clk), .r (Fresh[444]), .c ({signal_2662, signal_1596}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2553, signal_1499}), .a ({signal_2433, signal_1383}), .clk (clk), .r (Fresh[445]), .c ({signal_2663, signal_1597}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2555, signal_1501}), .a ({signal_2554, signal_1500}), .clk (clk), .r (Fresh[446]), .c ({signal_2664, signal_1598}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2554, signal_1500}), .a ({signal_2555, signal_1501}), .clk (clk), .r (Fresh[447]), .c ({signal_2665, signal_1599}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2555, signal_1501}), .a ({signal_2554, signal_1500}), .clk (clk), .r (Fresh[448]), .c ({signal_2666, signal_1600}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2554, signal_1500}), .a ({signal_2555, signal_1501}), .clk (clk), .r (Fresh[449]), .c ({signal_2667, signal_1601}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .s ({signal_2079, signal_1134}), .b ({signal_2557, signal_1503}), .a ({signal_2556, signal_1502}), .clk (clk), .r (Fresh[450]), .c ({signal_2668, signal_1602}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1447 ( .s ({signal_2079, signal_1134}), .b ({signal_2556, signal_1502}), .a ({signal_2557, signal_1503}), .clk (clk), .r (Fresh[451]), .c ({signal_2669, signal_1603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1468 ( .s ({signal_2040, signal_1147}), .b ({signal_2597, signal_1533}), .a ({signal_2596, signal_1532}), .clk (clk), .r (Fresh[452]), .c ({signal_2710, signal_807}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1469 ( .s ({signal_2052, signal_1143}), .b ({signal_2599, signal_1535}), .a ({signal_2598, signal_1534}), .clk (clk), .r (Fresh[453]), .c ({signal_2711, signal_803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1470 ( .s ({signal_2064, signal_1139}), .b ({signal_2601, signal_1537}), .a ({signal_2600, signal_1536}), .clk (clk), .r (Fresh[454]), .c ({signal_2712, signal_799}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1483 ( .s ({signal_2043, signal_1146}), .b ({signal_2616, signal_1551}), .a ({signal_2615, signal_1550}), .clk (clk), .r (Fresh[455]), .c ({signal_2729, signal_806}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1484 ( .s ({signal_2055, signal_1142}), .b ({signal_2618, signal_1553}), .a ({signal_2617, signal_1552}), .clk (clk), .r (Fresh[456]), .c ({signal_2730, signal_802}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1485 ( .s ({signal_2067, signal_1138}), .b ({signal_2620, signal_1555}), .a ({signal_2619, signal_1554}), .clk (clk), .r (Fresh[457]), .c ({signal_2731, signal_798}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1504 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2629, signal_1563}), .a ({signal_2628, signal_1562}), .clk (clk), .r (Fresh[458]), .c ({signal_2750, signal_1654}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1505 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2628, signal_1562}), .a ({signal_2629, signal_1563}), .clk (clk), .r (Fresh[459]), .c ({signal_2751, signal_1655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1526 ( .s (signal_1028), .b ({signal_2639, signal_1573}), .a ({signal_2638, signal_1572}), .c ({signal_2772, signal_795}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1533 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2652, signal_1586}), .a ({signal_2546, signal_1492}), .clk (clk), .r (Fresh[460]), .c ({signal_2779, signal_1682}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1534 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2653, signal_1587}), .a ({signal_2547, signal_1493}), .clk (clk), .r (Fresh[461]), .c ({signal_2780, signal_1683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1543 ( .s (signal_943), .b ({signal_2669, signal_1603}), .a ({signal_2668, signal_1602}), .c ({signal_2789, signal_794}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1544 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2671, signal_1605}), .a ({signal_2670, signal_1604}), .clk (clk), .r (Fresh[462]), .c ({signal_2790, signal_1692}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1545 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2670, signal_1604}), .a ({signal_2671, signal_1605}), .clk (clk), .r (Fresh[463]), .c ({signal_2791, signal_1693}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1546 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2673, signal_1607}), .a ({signal_2672, signal_1606}), .clk (clk), .r (Fresh[464]), .c ({signal_2792, signal_1694}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1547 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2672, signal_1606}), .a ({signal_2673, signal_1607}), .clk (clk), .r (Fresh[465]), .c ({signal_2793, signal_1695}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1548 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2675, signal_1609}), .a ({signal_2674, signal_1608}), .clk (clk), .r (Fresh[466]), .c ({signal_2794, signal_1696}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1549 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2674, signal_1608}), .a ({signal_2675, signal_1609}), .clk (clk), .r (Fresh[467]), .c ({signal_2795, signal_1697}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1550 ( .s ({Ciphertext_s1[23], Ciphertext_s0[23]}), .b ({signal_2675, signal_1609}), .a ({signal_2674, signal_1608}), .clk (clk), .r (Fresh[468]), .c ({signal_2796, signal_1698}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1551 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2674, signal_1608}), .a ({signal_2675, signal_1609}), .clk (clk), .r (Fresh[469]), .c ({signal_2797, signal_1699}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1552 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2677, signal_1611}), .a ({signal_2676, signal_1610}), .clk (clk), .r (Fresh[470]), .c ({signal_2798, signal_1700}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1553 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2676, signal_1610}), .a ({signal_2677, signal_1611}), .clk (clk), .r (Fresh[471]), .c ({signal_2799, signal_1701}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1554 ( .s ({Ciphertext_s1[19], Ciphertext_s0[19]}), .b ({signal_2677, signal_1611}), .a ({signal_2676, signal_1610}), .clk (clk), .r (Fresh[472]), .c ({signal_2800, signal_1702}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1555 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2676, signal_1610}), .a ({signal_2677, signal_1611}), .clk (clk), .r (Fresh[473]), .c ({signal_2801, signal_1703}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1456 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2581, signal_1520}), .a ({signal_2467, signal_1416}), .clk (clk), .r (Fresh[474]), .c ({signal_2695, signal_1612}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1457 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2582, signal_1521}), .a ({signal_2468, signal_1417}), .clk (clk), .r (Fresh[475]), .c ({signal_2696, signal_1613}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1458 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2584, signal_1522}), .a ({signal_2470, signal_1418}), .clk (clk), .r (Fresh[476]), .c ({signal_2698, signal_1614}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1459 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2585, signal_1523}), .a ({signal_2471, signal_1419}), .clk (clk), .r (Fresh[477]), .c ({signal_2699, signal_1615}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1460 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2587, signal_1524}), .a ({signal_2473, signal_1420}), .clk (clk), .r (Fresh[478]), .c ({signal_2701, signal_1616}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1461 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2588, signal_1525}), .a ({signal_2474, signal_1421}), .clk (clk), .r (Fresh[479]), .c ({signal_2702, signal_1617}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1462 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2589, signal_1526}), .a ({signal_2475, signal_1422}), .clk (clk), .r (Fresh[480]), .c ({signal_2703, signal_1618}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1463 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2590, signal_1527}), .a ({signal_2476, signal_1423}), .clk (clk), .r (Fresh[481]), .c ({signal_2704, signal_1619}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1464 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2591, signal_1528}), .a ({signal_2477, signal_1424}), .clk (clk), .r (Fresh[482]), .c ({signal_2705, signal_1620}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1465 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2592, signal_1529}), .a ({signal_2478, signal_1425}), .clk (clk), .r (Fresh[483]), .c ({signal_2706, signal_1621}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1466 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2594, signal_1530}), .a ({signal_2480, signal_1426}), .clk (clk), .r (Fresh[484]), .c ({signal_2708, signal_1622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1467 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2595, signal_1531}), .a ({signal_2481, signal_1427}), .clk (clk), .r (Fresh[485]), .c ({signal_2709, signal_1623}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1471 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2604, signal_1539}), .a ({signal_2603, signal_1538}), .clk (clk), .r (Fresh[486]), .c ({signal_2714, signal_1624}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1472 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2603, signal_1538}), .a ({signal_2604, signal_1539}), .clk (clk), .r (Fresh[487]), .c ({signal_2715, signal_1625}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1473 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2606, signal_1541}), .a ({signal_2605, signal_1540}), .clk (clk), .r (Fresh[488]), .c ({signal_2717, signal_1626}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1474 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2605, signal_1540}), .a ({signal_2606, signal_1541}), .clk (clk), .r (Fresh[489]), .c ({signal_2718, signal_1627}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1475 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2608, signal_1543}), .a ({signal_2607, signal_1542}), .clk (clk), .r (Fresh[490]), .c ({signal_2720, signal_1628}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1476 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2607, signal_1542}), .a ({signal_2608, signal_1543}), .clk (clk), .r (Fresh[491]), .c ({signal_2721, signal_1629}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1477 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2610, signal_1545}), .a ({signal_2609, signal_1544}), .clk (clk), .r (Fresh[492]), .c ({signal_2722, signal_1630}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1478 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2609, signal_1544}), .a ({signal_2610, signal_1545}), .clk (clk), .r (Fresh[493]), .c ({signal_2723, signal_1631}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1479 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2612, signal_1547}), .a ({signal_2611, signal_1546}), .clk (clk), .r (Fresh[494]), .c ({signal_2724, signal_1632}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1480 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2611, signal_1546}), .a ({signal_2612, signal_1547}), .clk (clk), .r (Fresh[495]), .c ({signal_2725, signal_1633}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1481 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2614, signal_1549}), .a ({signal_2613, signal_1548}), .clk (clk), .r (Fresh[496]), .c ({signal_2727, signal_1634}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1482 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2613, signal_1548}), .a ({signal_2614, signal_1549}), .clk (clk), .r (Fresh[497]), .c ({signal_2728, signal_1635}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1486 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2622, signal_1556}), .a ({signal_2522, signal_1468}), .clk (clk), .r (Fresh[498]), .c ({signal_2732, signal_1636}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1487 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2522, signal_1468}), .a ({signal_2622, signal_1556}), .clk (clk), .r (Fresh[499]), .c ({signal_2733, signal_1637}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1488 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2622, signal_1556}), .a ({signal_2623, signal_1557}), .clk (clk), .r (Fresh[500]), .c ({signal_2734, signal_1638}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1489 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2623, signal_1557}), .a ({signal_2523, signal_1469}), .clk (clk), .r (Fresh[501]), .c ({signal_2735, signal_1639}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1490 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2523, signal_1469}), .a ({signal_2623, signal_1557}), .clk (clk), .r (Fresh[502]), .c ({signal_2736, signal_1640}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1491 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2623, signal_1557}), .a ({signal_2622, signal_1556}), .clk (clk), .r (Fresh[503]), .c ({signal_2737, signal_1641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1492 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2624, signal_1558}), .a ({signal_2524, signal_1470}), .clk (clk), .r (Fresh[504]), .c ({signal_2738, signal_1642}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1493 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2524, signal_1470}), .a ({signal_2624, signal_1558}), .clk (clk), .r (Fresh[505]), .c ({signal_2739, signal_1643}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1494 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2624, signal_1558}), .a ({signal_2625, signal_1559}), .clk (clk), .r (Fresh[506]), .c ({signal_2740, signal_1644}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1495 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2625, signal_1559}), .a ({signal_2525, signal_1471}), .clk (clk), .r (Fresh[507]), .c ({signal_2741, signal_1645}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1496 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2525, signal_1471}), .a ({signal_2625, signal_1559}), .clk (clk), .r (Fresh[508]), .c ({signal_2742, signal_1646}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1497 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2625, signal_1559}), .a ({signal_2624, signal_1558}), .clk (clk), .r (Fresh[509]), .c ({signal_2743, signal_1647}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1498 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2626, signal_1560}), .a ({signal_2526, signal_1472}), .clk (clk), .r (Fresh[510]), .c ({signal_2744, signal_1648}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1499 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2526, signal_1472}), .a ({signal_2626, signal_1560}), .clk (clk), .r (Fresh[511]), .c ({signal_2745, signal_1649}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1500 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2626, signal_1560}), .a ({signal_2627, signal_1561}), .clk (clk), .r (Fresh[512]), .c ({signal_2746, signal_1650}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1501 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2627, signal_1561}), .a ({signal_2527, signal_1473}), .clk (clk), .r (Fresh[513]), .c ({signal_2747, signal_1651}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1502 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2527, signal_1473}), .a ({signal_2627, signal_1561}), .clk (clk), .r (Fresh[514]), .c ({signal_2748, signal_1652}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1503 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2627, signal_1561}), .a ({signal_2626, signal_1560}), .clk (clk), .r (Fresh[515]), .c ({signal_2749, signal_1653}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1506 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2630, signal_1564}), .a ({signal_2530, signal_1476}), .clk (clk), .r (Fresh[516]), .c ({signal_2752, signal_1656}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1507 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2530, signal_1476}), .a ({signal_2630, signal_1564}), .clk (clk), .r (Fresh[517]), .c ({signal_2753, signal_1657}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1508 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2630, signal_1564}), .a ({signal_2631, signal_1565}), .clk (clk), .r (Fresh[518]), .c ({signal_2754, signal_1658}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1509 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2631, signal_1565}), .a ({signal_2531, signal_1477}), .clk (clk), .r (Fresh[519]), .c ({signal_2755, signal_1659}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1510 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2531, signal_1477}), .a ({signal_2631, signal_1565}), .clk (clk), .r (Fresh[520]), .c ({signal_2756, signal_1660}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1511 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2631, signal_1565}), .a ({signal_2630, signal_1564}), .clk (clk), .r (Fresh[521]), .c ({signal_2757, signal_1661}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1512 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2632, signal_1566}), .a ({signal_2532, signal_1478}), .clk (clk), .r (Fresh[522]), .c ({signal_2758, signal_1662}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1513 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2532, signal_1478}), .a ({signal_2632, signal_1566}), .clk (clk), .r (Fresh[523]), .c ({signal_2759, signal_1663}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1514 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2632, signal_1566}), .a ({signal_2633, signal_1567}), .clk (clk), .r (Fresh[524]), .c ({signal_2760, signal_1664}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1515 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2633, signal_1567}), .a ({signal_2533, signal_1479}), .clk (clk), .r (Fresh[525]), .c ({signal_2761, signal_1665}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1516 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2533, signal_1479}), .a ({signal_2633, signal_1567}), .clk (clk), .r (Fresh[526]), .c ({signal_2762, signal_1666}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1517 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2633, signal_1567}), .a ({signal_2632, signal_1566}), .clk (clk), .r (Fresh[527]), .c ({signal_2763, signal_1667}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1518 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2634, signal_1568}), .a ({signal_2534, signal_1480}), .clk (clk), .r (Fresh[528]), .c ({signal_2764, signal_1668}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1519 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2635, signal_1569}), .a ({signal_2535, signal_1481}), .clk (clk), .r (Fresh[529]), .c ({signal_2765, signal_1669}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1520 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2636, signal_1570}), .a ({signal_2536, signal_1482}), .clk (clk), .r (Fresh[530]), .c ({signal_2766, signal_1670}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1521 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2536, signal_1482}), .a ({signal_2636, signal_1570}), .clk (clk), .r (Fresh[531]), .c ({signal_2767, signal_1671}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1522 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2636, signal_1570}), .a ({signal_2637, signal_1571}), .clk (clk), .r (Fresh[532]), .c ({signal_2768, signal_1672}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1523 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2637, signal_1571}), .a ({signal_2537, signal_1483}), .clk (clk), .r (Fresh[533]), .c ({signal_2769, signal_1673}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1524 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2537, signal_1483}), .a ({signal_2637, signal_1571}), .clk (clk), .r (Fresh[534]), .c ({signal_2770, signal_1674}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1525 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2637, signal_1571}), .a ({signal_2636, signal_1570}), .clk (clk), .r (Fresh[535]), .c ({signal_2771, signal_1675}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1527 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2641, signal_1575}), .a ({signal_2540, signal_1486}), .clk (clk), .r (Fresh[536]), .c ({signal_2773, signal_1676}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1528 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2642, signal_1576}), .a ({signal_2541, signal_1487}), .clk (clk), .r (Fresh[537]), .c ({signal_2774, signal_1677}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1529 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2645, signal_1579}), .a ({signal_2542, signal_1488}), .clk (clk), .r (Fresh[538]), .c ({signal_2775, signal_1678}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1530 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2646, signal_1580}), .a ({signal_2543, signal_1489}), .clk (clk), .r (Fresh[539]), .c ({signal_2776, signal_1679}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1531 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2649, signal_1583}), .a ({signal_2544, signal_1490}), .clk (clk), .r (Fresh[540]), .c ({signal_2777, signal_1680}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1532 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2650, signal_1584}), .a ({signal_2545, signal_1491}), .clk (clk), .r (Fresh[541]), .c ({signal_2778, signal_1681}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1535 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2655, signal_1589}), .a ({signal_2548, signal_1494}), .clk (clk), .r (Fresh[542]), .c ({signal_2781, signal_1684}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1536 ( .s ({Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({signal_2656, signal_1590}), .a ({signal_2549, signal_1495}), .clk (clk), .r (Fresh[543]), .c ({signal_2782, signal_1685}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1537 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2659, signal_1593}), .a ({signal_2550, signal_1496}), .clk (clk), .r (Fresh[544]), .c ({signal_2783, signal_1686}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1538 ( .s ({Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({signal_2660, signal_1594}), .a ({signal_2551, signal_1497}), .clk (clk), .r (Fresh[545]), .c ({signal_2784, signal_1687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1539 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2663, signal_1597}), .a ({signal_2662, signal_1596}), .clk (clk), .r (Fresh[546]), .c ({signal_2785, signal_1688}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1540 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2662, signal_1596}), .a ({signal_2663, signal_1597}), .clk (clk), .r (Fresh[547]), .c ({signal_2786, signal_1689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1541 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2665, signal_1599}), .a ({signal_2554, signal_1500}), .clk (clk), .r (Fresh[548]), .c ({signal_2787, signal_1690}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1542 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2666, signal_1600}), .a ({signal_2555, signal_1501}), .clk (clk), .r (Fresh[549]), .c ({signal_2788, signal_1691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1592 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2750, signal_1654}), .a ({signal_2628, signal_1562}), .clk (clk), .r (Fresh[550]), .c ({signal_2857, signal_1728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1593 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2751, signal_1655}), .a ({signal_2629, signal_1563}), .clk (clk), .r (Fresh[551]), .c ({signal_2858, signal_1729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1619 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2780, signal_1683}), .a ({signal_2779, signal_1682}), .clk (clk), .r (Fresh[552]), .c ({signal_2884, signal_1754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1620 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2779, signal_1682}), .a ({signal_2780, signal_1683}), .clk (clk), .r (Fresh[553]), .c ({signal_2885, signal_1755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1634 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2790, signal_1692}), .a ({signal_2670, signal_1604}), .clk (clk), .r (Fresh[554]), .c ({signal_2899, signal_1768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1635 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2670, signal_1604}), .a ({signal_2790, signal_1692}), .clk (clk), .r (Fresh[555]), .c ({signal_2900, signal_1769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1636 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2790, signal_1692}), .a ({signal_2791, signal_1693}), .clk (clk), .r (Fresh[556]), .c ({signal_2901, signal_1770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1637 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2791, signal_1693}), .a ({signal_2671, signal_1605}), .clk (clk), .r (Fresh[557]), .c ({signal_2902, signal_1771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1638 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2671, signal_1605}), .a ({signal_2791, signal_1693}), .clk (clk), .r (Fresh[558]), .c ({signal_2903, signal_1772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1639 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2791, signal_1693}), .a ({signal_2790, signal_1692}), .clk (clk), .r (Fresh[559]), .c ({signal_2904, signal_1773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1640 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2792, signal_1694}), .a ({signal_2672, signal_1606}), .clk (clk), .r (Fresh[560]), .c ({signal_2905, signal_1774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1641 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2672, signal_1606}), .a ({signal_2792, signal_1694}), .clk (clk), .r (Fresh[561]), .c ({signal_2906, signal_1775}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1642 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2792, signal_1694}), .a ({signal_2793, signal_1695}), .clk (clk), .r (Fresh[562]), .c ({signal_2907, signal_1776}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1643 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2793, signal_1695}), .a ({signal_2673, signal_1607}), .clk (clk), .r (Fresh[563]), .c ({signal_2908, signal_1777}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1644 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2673, signal_1607}), .a ({signal_2793, signal_1695}), .clk (clk), .r (Fresh[564]), .c ({signal_2909, signal_1778}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1645 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2793, signal_1695}), .a ({signal_2792, signal_1694}), .clk (clk), .r (Fresh[565]), .c ({signal_2910, signal_1779}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1646 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2795, signal_1697}), .a ({signal_2674, signal_1608}), .clk (clk), .r (Fresh[566]), .c ({signal_2911, signal_1780}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1647 ( .s ({Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({signal_2796, signal_1698}), .a ({signal_2675, signal_1609}), .clk (clk), .r (Fresh[567]), .c ({signal_2912, signal_1781}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1648 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2799, signal_1701}), .a ({signal_2676, signal_1610}), .clk (clk), .r (Fresh[568]), .c ({signal_2913, signal_1782}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1649 ( .s ({Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({signal_2800, signal_1702}), .a ({signal_2677, signal_1611}), .clk (clk), .r (Fresh[569]), .c ({signal_2914, signal_1783}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_2 ( .s (rst), .b ({signal_2818, signal_837}), .a ({Plaintext_s1[2], Plaintext_s0[2]}), .c ({signal_2916, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3 ( .s (rst), .b ({signal_2833, signal_836}), .a ({Plaintext_s1[3], Plaintext_s0[3]}), .c ({signal_2918, signal_900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_6 ( .s (rst), .b ({signal_2819, signal_833}), .a ({Plaintext_s1[6], Plaintext_s0[6]}), .c ({signal_2920, signal_897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_7 ( .s (rst), .b ({signal_2834, signal_832}), .a ({Plaintext_s1[7], Plaintext_s0[7]}), .c ({signal_2922, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_10 ( .s (rst), .b ({signal_2820, signal_829}), .a ({Plaintext_s1[10], Plaintext_s0[10]}), .c ({signal_2924, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_11 ( .s (rst), .b ({signal_2835, signal_828}), .a ({Plaintext_s1[11], Plaintext_s0[11]}), .c ({signal_2926, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_14 ( .s (rst), .b ({signal_3028, signal_825}), .a ({Plaintext_s1[14], Plaintext_s0[14]}), .c ({signal_3083, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_15 ( .s (rst), .b ({signal_3044, signal_824}), .a ({Plaintext_s1[15], Plaintext_s0[15]}), .c ({signal_3085, signal_888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_18 ( .s (rst), .b ({signal_2821, signal_821}), .a ({Plaintext_s1[18], Plaintext_s0[18]}), .c ({signal_2928, signal_885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_19 ( .s (rst), .b ({signal_2836, signal_820}), .a ({Plaintext_s1[19], Plaintext_s0[19]}), .c ({signal_2930, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_22 ( .s (rst), .b ({signal_2822, signal_817}), .a ({Plaintext_s1[22], Plaintext_s0[22]}), .c ({signal_2932, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_23 ( .s (rst), .b ({signal_2837, signal_816}), .a ({Plaintext_s1[23], Plaintext_s0[23]}), .c ({signal_2934, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_26 ( .s (rst), .b ({signal_2867, signal_813}), .a ({Plaintext_s1[26], Plaintext_s0[26]}), .c ({signal_2936, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_27 ( .s (rst), .b ({signal_2894, signal_812}), .a ({Plaintext_s1[27], Plaintext_s0[27]}), .c ({signal_2938, signal_876}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_30 ( .s (rst), .b ({signal_2823, signal_809}), .a ({Plaintext_s1[30], Plaintext_s0[30]}), .c ({signal_2940, signal_873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_31 ( .s (rst), .b ({signal_2838, signal_808}), .a ({Plaintext_s1[31], Plaintext_s0[31]}), .c ({signal_2942, signal_872}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1556 ( .s ({signal_2046, signal_1145}), .b ({signal_2696, signal_1613}), .a ({signal_2695, signal_1612}), .clk (clk), .r (Fresh[570]), .c ({signal_2818, signal_837}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1557 ( .s ({signal_2058, signal_1141}), .b ({signal_2699, signal_1615}), .a ({signal_2698, signal_1614}), .clk (clk), .r (Fresh[571]), .c ({signal_2819, signal_833}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1558 ( .s ({signal_2070, signal_1137}), .b ({signal_2702, signal_1617}), .a ({signal_2701, signal_1616}), .clk (clk), .r (Fresh[572]), .c ({signal_2820, signal_829}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1559 ( .s ({signal_2010, signal_1157}), .b ({signal_2704, signal_1619}), .a ({signal_2703, signal_1618}), .clk (clk), .r (Fresh[573]), .c ({signal_2821, signal_821}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1560 ( .s ({signal_2022, signal_1153}), .b ({signal_2706, signal_1621}), .a ({signal_2705, signal_1620}), .clk (clk), .r (Fresh[574]), .c ({signal_2822, signal_817}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1561 ( .s ({signal_1998, signal_1161}), .b ({signal_2709, signal_1623}), .a ({signal_2708, signal_1622}), .clk (clk), .r (Fresh[575]), .c ({signal_2823, signal_809}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1562 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2695, signal_1612}), .a ({signal_2696, signal_1613}), .clk (clk), .r (Fresh[576]), .c ({signal_2825, signal_1704}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1563 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2696, signal_1613}), .a ({signal_2695, signal_1612}), .clk (clk), .r (Fresh[577]), .c ({signal_2826, signal_1705}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1564 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2698, signal_1614}), .a ({signal_2699, signal_1615}), .clk (clk), .r (Fresh[578]), .c ({signal_2828, signal_1706}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1565 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2699, signal_1615}), .a ({signal_2698, signal_1614}), .clk (clk), .r (Fresh[579]), .c ({signal_2829, signal_1707}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1566 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2701, signal_1616}), .a ({signal_2702, signal_1617}), .clk (clk), .r (Fresh[580]), .c ({signal_2831, signal_1708}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1567 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2702, signal_1617}), .a ({signal_2701, signal_1616}), .clk (clk), .r (Fresh[581]), .c ({signal_2832, signal_1709}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1568 ( .s ({signal_2049, signal_1144}), .b ({signal_2715, signal_1625}), .a ({signal_2714, signal_1624}), .clk (clk), .r (Fresh[582]), .c ({signal_2833, signal_836}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1569 ( .s ({signal_2061, signal_1140}), .b ({signal_2718, signal_1627}), .a ({signal_2717, signal_1626}), .clk (clk), .r (Fresh[583]), .c ({signal_2834, signal_832}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1570 ( .s ({signal_2073, signal_1136}), .b ({signal_2721, signal_1629}), .a ({signal_2720, signal_1628}), .clk (clk), .r (Fresh[584]), .c ({signal_2835, signal_828}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1571 ( .s ({signal_2013, signal_1156}), .b ({signal_2723, signal_1631}), .a ({signal_2722, signal_1630}), .clk (clk), .r (Fresh[585]), .c ({signal_2836, signal_820}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1572 ( .s ({signal_2025, signal_1152}), .b ({signal_2725, signal_1633}), .a ({signal_2724, signal_1632}), .clk (clk), .r (Fresh[586]), .c ({signal_2837, signal_816}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1573 ( .s ({signal_2001, signal_1160}), .b ({signal_2728, signal_1635}), .a ({signal_2727, signal_1634}), .clk (clk), .r (Fresh[587]), .c ({signal_2838, signal_808}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1574 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2714, signal_1624}), .a ({signal_2715, signal_1625}), .clk (clk), .r (Fresh[588]), .c ({signal_2839, signal_1710}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1575 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2715, signal_1625}), .a ({signal_2714, signal_1624}), .clk (clk), .r (Fresh[589]), .c ({signal_2840, signal_1711}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1576 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2717, signal_1626}), .a ({signal_2718, signal_1627}), .clk (clk), .r (Fresh[590]), .c ({signal_2841, signal_1712}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1577 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2718, signal_1627}), .a ({signal_2717, signal_1626}), .clk (clk), .r (Fresh[591]), .c ({signal_2842, signal_1713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1578 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2720, signal_1628}), .a ({signal_2721, signal_1629}), .clk (clk), .r (Fresh[592]), .c ({signal_2843, signal_1714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1579 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2721, signal_1629}), .a ({signal_2720, signal_1628}), .clk (clk), .r (Fresh[593]), .c ({signal_2844, signal_1715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1580 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2523, signal_1469}), .a ({signal_2732, signal_1636}), .clk (clk), .r (Fresh[594]), .c ({signal_2845, signal_1716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1581 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2734, signal_1638}), .a ({signal_2733, signal_1637}), .clk (clk), .r (Fresh[595]), .c ({signal_2846, signal_1717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1582 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2522, signal_1468}), .a ({signal_2735, signal_1639}), .clk (clk), .r (Fresh[596]), .c ({signal_2847, signal_1718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1583 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2737, signal_1641}), .a ({signal_2736, signal_1640}), .clk (clk), .r (Fresh[597]), .c ({signal_2848, signal_1719}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1584 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2525, signal_1471}), .a ({signal_2738, signal_1642}), .clk (clk), .r (Fresh[598]), .c ({signal_2849, signal_1720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1585 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2740, signal_1644}), .a ({signal_2739, signal_1643}), .clk (clk), .r (Fresh[599]), .c ({signal_2850, signal_1721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1586 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2524, signal_1470}), .a ({signal_2741, signal_1645}), .clk (clk), .r (Fresh[600]), .c ({signal_2851, signal_1722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1587 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2743, signal_1647}), .a ({signal_2742, signal_1646}), .clk (clk), .r (Fresh[601]), .c ({signal_2852, signal_1723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1588 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2527, signal_1473}), .a ({signal_2744, signal_1648}), .clk (clk), .r (Fresh[602]), .c ({signal_2853, signal_1724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1589 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2746, signal_1650}), .a ({signal_2745, signal_1649}), .clk (clk), .r (Fresh[603]), .c ({signal_2854, signal_1725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1590 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2526, signal_1472}), .a ({signal_2747, signal_1651}), .clk (clk), .r (Fresh[604]), .c ({signal_2855, signal_1726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1591 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2749, signal_1653}), .a ({signal_2748, signal_1652}), .clk (clk), .r (Fresh[605]), .c ({signal_2856, signal_1727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1594 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2531, signal_1477}), .a ({signal_2752, signal_1656}), .clk (clk), .r (Fresh[606]), .c ({signal_2859, signal_1730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1595 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2754, signal_1658}), .a ({signal_2753, signal_1657}), .clk (clk), .r (Fresh[607]), .c ({signal_2860, signal_1731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1596 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2530, signal_1476}), .a ({signal_2755, signal_1659}), .clk (clk), .r (Fresh[608]), .c ({signal_2861, signal_1732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1597 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2757, signal_1661}), .a ({signal_2756, signal_1660}), .clk (clk), .r (Fresh[609]), .c ({signal_2862, signal_1733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1598 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2533, signal_1479}), .a ({signal_2758, signal_1662}), .clk (clk), .r (Fresh[610]), .c ({signal_2863, signal_1734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1599 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2760, signal_1664}), .a ({signal_2759, signal_1663}), .clk (clk), .r (Fresh[611]), .c ({signal_2864, signal_1735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1600 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2532, signal_1478}), .a ({signal_2761, signal_1665}), .clk (clk), .r (Fresh[612]), .c ({signal_2865, signal_1736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1601 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2763, signal_1667}), .a ({signal_2762, signal_1666}), .clk (clk), .r (Fresh[613]), .c ({signal_2866, signal_1737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1602 ( .s ({signal_2034, signal_1149}), .b ({signal_2765, signal_1669}), .a ({signal_2764, signal_1668}), .clk (clk), .r (Fresh[614]), .c ({signal_2867, signal_813}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1603 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2537, signal_1483}), .a ({signal_2766, signal_1670}), .clk (clk), .r (Fresh[615]), .c ({signal_2868, signal_1738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1604 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2768, signal_1672}), .a ({signal_2767, signal_1671}), .clk (clk), .r (Fresh[616]), .c ({signal_2869, signal_1739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1605 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2536, signal_1482}), .a ({signal_2769, signal_1673}), .clk (clk), .r (Fresh[617]), .c ({signal_2870, signal_1740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1606 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2771, signal_1675}), .a ({signal_2770, signal_1674}), .clk (clk), .r (Fresh[618]), .c ({signal_2871, signal_1741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1607 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2773, signal_1676}), .a ({signal_2640, signal_1574}), .clk (clk), .r (Fresh[619]), .c ({signal_2872, signal_1742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1608 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2774, signal_1677}), .a ({signal_2640, signal_1574}), .clk (clk), .r (Fresh[620]), .c ({signal_2873, signal_1743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1609 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2774, signal_1677}), .a ({signal_2643, signal_1577}), .clk (clk), .r (Fresh[621]), .c ({signal_2874, signal_1744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1610 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2773, signal_1676}), .a ({signal_2643, signal_1577}), .clk (clk), .r (Fresh[622]), .c ({signal_2875, signal_1745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1611 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2775, signal_1678}), .a ({signal_2644, signal_1578}), .clk (clk), .r (Fresh[623]), .c ({signal_2876, signal_1746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1612 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2776, signal_1679}), .a ({signal_2644, signal_1578}), .clk (clk), .r (Fresh[624]), .c ({signal_2877, signal_1747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1613 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2776, signal_1679}), .a ({signal_2647, signal_1581}), .clk (clk), .r (Fresh[625]), .c ({signal_2878, signal_1748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1614 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2775, signal_1678}), .a ({signal_2647, signal_1581}), .clk (clk), .r (Fresh[626]), .c ({signal_2879, signal_1749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1615 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2777, signal_1680}), .a ({signal_2648, signal_1582}), .clk (clk), .r (Fresh[627]), .c ({signal_2880, signal_1750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1616 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2778, signal_1681}), .a ({signal_2648, signal_1582}), .clk (clk), .r (Fresh[628]), .c ({signal_2881, signal_1751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1617 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2778, signal_1681}), .a ({signal_2651, signal_1585}), .clk (clk), .r (Fresh[629]), .c ({signal_2882, signal_1752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1618 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2777, signal_1680}), .a ({signal_2651, signal_1585}), .clk (clk), .r (Fresh[630]), .c ({signal_2883, signal_1753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1621 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2781, signal_1684}), .a ({signal_2654, signal_1588}), .clk (clk), .r (Fresh[631]), .c ({signal_2886, signal_1756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1622 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2782, signal_1685}), .a ({signal_2654, signal_1588}), .clk (clk), .r (Fresh[632]), .c ({signal_2887, signal_1757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1623 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2782, signal_1685}), .a ({signal_2657, signal_1591}), .clk (clk), .r (Fresh[633]), .c ({signal_2888, signal_1758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1624 ( .s ({Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({signal_2781, signal_1684}), .a ({signal_2657, signal_1591}), .clk (clk), .r (Fresh[634]), .c ({signal_2889, signal_1759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1625 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2783, signal_1686}), .a ({signal_2658, signal_1592}), .clk (clk), .r (Fresh[635]), .c ({signal_2890, signal_1760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1626 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2784, signal_1687}), .a ({signal_2658, signal_1592}), .clk (clk), .r (Fresh[636]), .c ({signal_2891, signal_1761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1627 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2784, signal_1687}), .a ({signal_2661, signal_1595}), .clk (clk), .r (Fresh[637]), .c ({signal_2892, signal_1762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1628 ( .s ({Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({signal_2783, signal_1686}), .a ({signal_2661, signal_1595}), .clk (clk), .r (Fresh[638]), .c ({signal_2893, signal_1763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1629 ( .s ({signal_2037, signal_1148}), .b ({signal_2786, signal_1689}), .a ({signal_2785, signal_1688}), .clk (clk), .r (Fresh[639]), .c ({signal_2894, signal_812}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1630 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2787, signal_1690}), .a ({signal_2664, signal_1598}), .clk (clk), .r (Fresh[640]), .c ({signal_2895, signal_1764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1631 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2788, signal_1691}), .a ({signal_2664, signal_1598}), .clk (clk), .r (Fresh[641]), .c ({signal_2896, signal_1765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1632 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2788, signal_1691}), .a ({signal_2667, signal_1601}), .clk (clk), .r (Fresh[642]), .c ({signal_2897, signal_1766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1633 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2787, signal_1690}), .a ({signal_2667, signal_1601}), .clk (clk), .r (Fresh[643]), .c ({signal_2898, signal_1767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1668 ( .s ({signal_2082, signal_1133}), .b ({signal_2858, signal_1729}), .a ({signal_2857, signal_1728}), .clk (clk), .r (Fresh[644]), .c ({signal_2964, signal_1802}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1669 ( .s ({signal_2082, signal_1133}), .b ({signal_2857, signal_1728}), .a ({signal_2858, signal_1729}), .clk (clk), .r (Fresh[645]), .c ({signal_2965, signal_1803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1676 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_2857, signal_1728}), .a ({signal_2858, signal_1729}), .clk (clk), .r (Fresh[646]), .c ({signal_2973, signal_1810}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1677 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_2858, signal_1729}), .a ({signal_2857, signal_1728}), .clk (clk), .r (Fresh[647]), .c ({signal_2974, signal_1811}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1684 ( .s ({signal_2085, signal_1132}), .b ({signal_2885, signal_1755}), .a ({signal_2884, signal_1754}), .clk (clk), .r (Fresh[648]), .c ({signal_2981, signal_1818}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1685 ( .s ({signal_2085, signal_1132}), .b ({signal_2884, signal_1754}), .a ({signal_2885, signal_1755}), .clk (clk), .r (Fresh[649]), .c ({signal_2982, signal_1819}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1692 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_2884, signal_1754}), .a ({signal_2885, signal_1755}), .clk (clk), .r (Fresh[650]), .c ({signal_2989, signal_1826}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1693 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_2885, signal_1755}), .a ({signal_2884, signal_1754}), .clk (clk), .r (Fresh[651]), .c ({signal_2990, signal_1827}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1694 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2671, signal_1605}), .a ({signal_2899, signal_1768}), .clk (clk), .r (Fresh[652]), .c ({signal_2991, signal_1828}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1695 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2901, signal_1770}), .a ({signal_2900, signal_1769}), .clk (clk), .r (Fresh[653]), .c ({signal_2992, signal_1829}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1696 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2670, signal_1604}), .a ({signal_2902, signal_1771}), .clk (clk), .r (Fresh[654]), .c ({signal_2993, signal_1830}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1697 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2904, signal_1773}), .a ({signal_2903, signal_1772}), .clk (clk), .r (Fresh[655]), .c ({signal_2994, signal_1831}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1698 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2673, signal_1607}), .a ({signal_2905, signal_1774}), .clk (clk), .r (Fresh[656]), .c ({signal_2995, signal_1832}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1699 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2907, signal_1776}), .a ({signal_2906, signal_1775}), .clk (clk), .r (Fresh[657]), .c ({signal_2996, signal_1833}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1700 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2672, signal_1606}), .a ({signal_2908, signal_1777}), .clk (clk), .r (Fresh[658]), .c ({signal_2997, signal_1834}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1701 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2910, signal_1779}), .a ({signal_2909, signal_1778}), .clk (clk), .r (Fresh[659]), .c ({signal_2998, signal_1835}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1702 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2911, signal_1780}), .a ({signal_2794, signal_1696}), .clk (clk), .r (Fresh[660]), .c ({signal_2999, signal_1836}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1703 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2912, signal_1781}), .a ({signal_2794, signal_1696}), .clk (clk), .r (Fresh[661]), .c ({signal_3000, signal_1837}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1704 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2912, signal_1781}), .a ({signal_2797, signal_1699}), .clk (clk), .r (Fresh[662]), .c ({signal_3001, signal_1838}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1705 ( .s ({Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({signal_2911, signal_1780}), .a ({signal_2797, signal_1699}), .clk (clk), .r (Fresh[663]), .c ({signal_3002, signal_1839}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1706 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2913, signal_1782}), .a ({signal_2798, signal_1700}), .clk (clk), .r (Fresh[664]), .c ({signal_3003, signal_1840}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1707 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2914, signal_1783}), .a ({signal_2798, signal_1700}), .clk (clk), .r (Fresh[665]), .c ({signal_3004, signal_1841}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1708 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2914, signal_1783}), .a ({signal_2801, signal_1703}), .clk (clk), .r (Fresh[666]), .c ({signal_3005, signal_1842}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1709 ( .s ({Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({signal_2913, signal_1782}), .a ({signal_2801, signal_1703}), .clk (clk), .r (Fresh[667]), .c ({signal_3006, signal_1843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1725 ( .s (signal_1026), .b ({signal_2965, signal_1803}), .a ({signal_2964, signal_1802}), .c ({signal_3028, signal_825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1740 ( .s (signal_1025), .b ({signal_2982, signal_1819}), .a ({signal_2981, signal_1818}), .c ({signal_3044, signal_824}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1650 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2826, signal_1705}), .a ({signal_2825, signal_1704}), .clk (clk), .r (Fresh[668]), .c ({signal_2944, signal_1784}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1651 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2825, signal_1704}), .a ({signal_2826, signal_1705}), .clk (clk), .r (Fresh[669]), .c ({signal_2945, signal_1785}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1652 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2829, signal_1707}), .a ({signal_2828, signal_1706}), .clk (clk), .r (Fresh[670]), .c ({signal_2947, signal_1786}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1653 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2828, signal_1706}), .a ({signal_2829, signal_1707}), .clk (clk), .r (Fresh[671]), .c ({signal_2948, signal_1787}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1654 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2832, signal_1709}), .a ({signal_2831, signal_1708}), .clk (clk), .r (Fresh[672]), .c ({signal_2950, signal_1788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1655 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2831, signal_1708}), .a ({signal_2832, signal_1709}), .clk (clk), .r (Fresh[673]), .c ({signal_2951, signal_1789}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1656 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2839, signal_1710}), .a ({signal_2715, signal_1625}), .clk (clk), .r (Fresh[674]), .c ({signal_2952, signal_1790}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1657 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2840, signal_1711}), .a ({signal_2714, signal_1624}), .clk (clk), .r (Fresh[675]), .c ({signal_2953, signal_1791}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1658 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2841, signal_1712}), .a ({signal_2718, signal_1627}), .clk (clk), .r (Fresh[676]), .c ({signal_2954, signal_1792}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1659 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2842, signal_1713}), .a ({signal_2717, signal_1626}), .clk (clk), .r (Fresh[677]), .c ({signal_2955, signal_1793}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1660 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2843, signal_1714}), .a ({signal_2721, signal_1629}), .clk (clk), .r (Fresh[678]), .c ({signal_2956, signal_1794}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1661 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2844, signal_1715}), .a ({signal_2720, signal_1628}), .clk (clk), .r (Fresh[679]), .c ({signal_2957, signal_1795}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1662 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2846, signal_1717}), .a ({signal_2845, signal_1716}), .clk (clk), .r (Fresh[680]), .c ({signal_2958, signal_1796}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1663 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2848, signal_1719}), .a ({signal_2847, signal_1718}), .clk (clk), .r (Fresh[681]), .c ({signal_2959, signal_1797}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1664 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2850, signal_1721}), .a ({signal_2849, signal_1720}), .clk (clk), .r (Fresh[682]), .c ({signal_2960, signal_1798}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1665 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2852, signal_1723}), .a ({signal_2851, signal_1722}), .clk (clk), .r (Fresh[683]), .c ({signal_2961, signal_1799}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1666 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2854, signal_1725}), .a ({signal_2853, signal_1724}), .clk (clk), .r (Fresh[684]), .c ({signal_2962, signal_1800}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1667 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2856, signal_1727}), .a ({signal_2855, signal_1726}), .clk (clk), .r (Fresh[685]), .c ({signal_2963, signal_1801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1670 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2860, signal_1731}), .a ({signal_2859, signal_1730}), .clk (clk), .r (Fresh[686]), .c ({signal_2966, signal_1804}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1671 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2862, signal_1733}), .a ({signal_2861, signal_1732}), .clk (clk), .r (Fresh[687]), .c ({signal_2967, signal_1805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1672 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2864, signal_1735}), .a ({signal_2863, signal_1734}), .clk (clk), .r (Fresh[688]), .c ({signal_2968, signal_1806}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1673 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2866, signal_1737}), .a ({signal_2865, signal_1736}), .clk (clk), .r (Fresh[689]), .c ({signal_2969, signal_1807}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1674 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2869, signal_1739}), .a ({signal_2868, signal_1738}), .clk (clk), .r (Fresh[690]), .c ({signal_2970, signal_1808}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1675 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2871, signal_1741}), .a ({signal_2870, signal_1740}), .clk (clk), .r (Fresh[691]), .c ({signal_2971, signal_1809}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1678 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2873, signal_1743}), .a ({signal_2872, signal_1742}), .clk (clk), .r (Fresh[692]), .c ({signal_2975, signal_1812}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1679 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2875, signal_1745}), .a ({signal_2874, signal_1744}), .clk (clk), .r (Fresh[693]), .c ({signal_2976, signal_1813}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1680 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2877, signal_1747}), .a ({signal_2876, signal_1746}), .clk (clk), .r (Fresh[694]), .c ({signal_2977, signal_1814}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1681 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2879, signal_1749}), .a ({signal_2878, signal_1748}), .clk (clk), .r (Fresh[695]), .c ({signal_2978, signal_1815}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1682 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2881, signal_1751}), .a ({signal_2880, signal_1750}), .clk (clk), .r (Fresh[696]), .c ({signal_2979, signal_1816}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1683 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2883, signal_1753}), .a ({signal_2882, signal_1752}), .clk (clk), .r (Fresh[697]), .c ({signal_2980, signal_1817}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1686 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2887, signal_1757}), .a ({signal_2886, signal_1756}), .clk (clk), .r (Fresh[698]), .c ({signal_2983, signal_1820}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1687 ( .s ({Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({signal_2889, signal_1759}), .a ({signal_2888, signal_1758}), .clk (clk), .r (Fresh[699]), .c ({signal_2984, signal_1821}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1688 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2891, signal_1761}), .a ({signal_2890, signal_1760}), .clk (clk), .r (Fresh[700]), .c ({signal_2985, signal_1822}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1689 ( .s ({Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({signal_2893, signal_1763}), .a ({signal_2892, signal_1762}), .clk (clk), .r (Fresh[701]), .c ({signal_2986, signal_1823}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1690 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2896, signal_1765}), .a ({signal_2895, signal_1764}), .clk (clk), .r (Fresh[702]), .c ({signal_2987, signal_1824}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1691 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2898, signal_1767}), .a ({signal_2897, signal_1766}), .clk (clk), .r (Fresh[703]), .c ({signal_2988, signal_1825}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1735 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_2974, signal_1811}), .a ({signal_2973, signal_1810}), .clk (clk), .r (Fresh[704]), .c ({signal_3039, signal_1862}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1736 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_2973, signal_1810}), .a ({signal_2974, signal_1811}), .clk (clk), .r (Fresh[705]), .c ({signal_3040, signal_1863}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1756 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_2989, signal_1826}), .a ({signal_2885, signal_1755}), .clk (clk), .r (Fresh[706]), .c ({signal_3060, signal_1876}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1757 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_2990, signal_1827}), .a ({signal_2884, signal_1754}), .clk (clk), .r (Fresh[707]), .c ({signal_3061, signal_1877}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1758 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2992, signal_1829}), .a ({signal_2991, signal_1828}), .clk (clk), .r (Fresh[708]), .c ({signal_3062, signal_1878}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1759 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_2994, signal_1831}), .a ({signal_2993, signal_1830}), .clk (clk), .r (Fresh[709]), .c ({signal_3063, signal_1879}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1760 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2996, signal_1833}), .a ({signal_2995, signal_1832}), .clk (clk), .r (Fresh[710]), .c ({signal_3064, signal_1880}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1761 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_2998, signal_1835}), .a ({signal_2997, signal_1834}), .clk (clk), .r (Fresh[711]), .c ({signal_3065, signal_1881}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1762 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_3000, signal_1837}), .a ({signal_2999, signal_1836}), .clk (clk), .r (Fresh[712]), .c ({signal_3066, signal_1882}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1763 ( .s ({Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({signal_3002, signal_1839}), .a ({signal_3001, signal_1838}), .clk (clk), .r (Fresh[713]), .c ({signal_3067, signal_1883}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1764 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_3004, signal_1841}), .a ({signal_3003, signal_1840}), .clk (clk), .r (Fresh[714]), .c ({signal_3068, signal_1884}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1765 ( .s ({Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({signal_3006, signal_1843}), .a ({signal_3005, signal_1842}), .clk (clk), .r (Fresh[715]), .c ({signal_3069, signal_1885}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_0 ( .s (rst), .b ({signal_3025, signal_839}), .a ({Plaintext_s1[0], Plaintext_s0[0]}), .c ({signal_3071, signal_903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1 ( .s (rst), .b ({signal_3041, signal_838}), .a ({Plaintext_s1[1], Plaintext_s0[1]}), .c ({signal_3073, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_4 ( .s (rst), .b ({signal_3026, signal_835}), .a ({Plaintext_s1[4], Plaintext_s0[4]}), .c ({signal_3075, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_5 ( .s (rst), .b ({signal_3042, signal_834}), .a ({Plaintext_s1[5], Plaintext_s0[5]}), .c ({signal_3077, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_8 ( .s (rst), .b ({signal_3027, signal_831}), .a ({Plaintext_s1[8], Plaintext_s0[8]}), .c ({signal_3079, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_9 ( .s (rst), .b ({signal_3043, signal_830}), .a ({Plaintext_s1[9], Plaintext_s0[9]}), .c ({signal_3081, signal_894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_12 ( .s (rst), .b ({signal_3188, signal_827}), .a ({Plaintext_s1[12], Plaintext_s0[12]}), .c ({signal_3201, signal_891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_13 ( .s (rst), .b ({signal_3196, signal_826}), .a ({Plaintext_s1[13], Plaintext_s0[13]}), .c ({signal_3203, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_16 ( .s (rst), .b ({signal_3029, signal_823}), .a ({Plaintext_s1[16], Plaintext_s0[16]}), .c ({signal_3087, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_17 ( .s (rst), .b ({signal_3045, signal_822}), .a ({Plaintext_s1[17], Plaintext_s0[17]}), .c ({signal_3089, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_20 ( .s (rst), .b ({signal_3030, signal_819}), .a ({Plaintext_s1[20], Plaintext_s0[20]}), .c ({signal_3091, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_21 ( .s (rst), .b ({signal_3046, signal_818}), .a ({Plaintext_s1[21], Plaintext_s0[21]}), .c ({signal_3093, signal_882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_24 ( .s (rst), .b ({signal_3189, signal_815}), .a ({Plaintext_s1[24], Plaintext_s0[24]}), .c ({signal_3205, signal_879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_25 ( .s (rst), .b ({signal_3197, signal_814}), .a ({Plaintext_s1[25], Plaintext_s0[25]}), .c ({signal_3207, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_28 ( .s (rst), .b ({signal_3031, signal_811}), .a ({Plaintext_s1[28], Plaintext_s0[28]}), .c ({signal_3095, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_29 ( .s (rst), .b ({signal_3047, signal_810}), .a ({Plaintext_s1[29], Plaintext_s0[29]}), .c ({signal_3097, signal_874}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1710 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_2944, signal_1784}), .a ({signal_2825, signal_1704}), .clk (clk), .r (Fresh[716]), .c ({signal_3008, signal_1844}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1711 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_2945, signal_1785}), .a ({signal_2826, signal_1705}), .clk (clk), .r (Fresh[717]), .c ({signal_3009, signal_1845}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1712 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_2947, signal_1786}), .a ({signal_2828, signal_1706}), .clk (clk), .r (Fresh[718]), .c ({signal_3011, signal_1846}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1713 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_2948, signal_1787}), .a ({signal_2829, signal_1707}), .clk (clk), .r (Fresh[719]), .c ({signal_3012, signal_1847}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1714 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_2950, signal_1788}), .a ({signal_2831, signal_1708}), .clk (clk), .r (Fresh[720]), .c ({signal_3014, signal_1848}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1715 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_2951, signal_1789}), .a ({signal_2832, signal_1709}), .clk (clk), .r (Fresh[721]), .c ({signal_3015, signal_1849}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1716 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_2953, signal_1791}), .a ({signal_2952, signal_1790}), .clk (clk), .r (Fresh[722]), .c ({signal_3017, signal_1850}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1717 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_2952, signal_1790}), .a ({signal_2953, signal_1791}), .clk (clk), .r (Fresh[723]), .c ({signal_3018, signal_1851}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1718 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_2955, signal_1793}), .a ({signal_2954, signal_1792}), .clk (clk), .r (Fresh[724]), .c ({signal_3020, signal_1852}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1719 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_2954, signal_1792}), .a ({signal_2955, signal_1793}), .clk (clk), .r (Fresh[725]), .c ({signal_3021, signal_1853}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1720 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_2957, signal_1795}), .a ({signal_2956, signal_1794}), .clk (clk), .r (Fresh[726]), .c ({signal_3023, signal_1854}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1721 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_2956, signal_1794}), .a ({signal_2957, signal_1795}), .clk (clk), .r (Fresh[727]), .c ({signal_3024, signal_1855}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1722 ( .s ({signal_2040, signal_1147}), .b ({signal_2959, signal_1797}), .a ({signal_2958, signal_1796}), .clk (clk), .r (Fresh[728]), .c ({signal_3025, signal_839}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1723 ( .s ({signal_2052, signal_1143}), .b ({signal_2961, signal_1799}), .a ({signal_2960, signal_1798}), .clk (clk), .r (Fresh[729]), .c ({signal_3026, signal_835}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1724 ( .s ({signal_2064, signal_1139}), .b ({signal_2963, signal_1801}), .a ({signal_2962, signal_1800}), .clk (clk), .r (Fresh[730]), .c ({signal_3027, signal_831}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1726 ( .s ({signal_2004, signal_1159}), .b ({signal_2967, signal_1805}), .a ({signal_2966, signal_1804}), .clk (clk), .r (Fresh[731]), .c ({signal_3029, signal_823}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1727 ( .s ({signal_2016, signal_1155}), .b ({signal_2969, signal_1807}), .a ({signal_2968, signal_1806}), .clk (clk), .r (Fresh[732]), .c ({signal_3030, signal_819}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1728 ( .s ({signal_1992, signal_1163}), .b ({signal_2971, signal_1809}), .a ({signal_2970, signal_1808}), .clk (clk), .r (Fresh[733]), .c ({signal_3031, signal_811}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1729 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2958, signal_1796}), .a ({signal_2959, signal_1797}), .clk (clk), .r (Fresh[734]), .c ({signal_3032, signal_1856}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1730 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2959, signal_1797}), .a ({signal_2958, signal_1796}), .clk (clk), .r (Fresh[735]), .c ({signal_3033, signal_1857}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1731 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2960, signal_1798}), .a ({signal_2961, signal_1799}), .clk (clk), .r (Fresh[736]), .c ({signal_3034, signal_1858}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1732 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2961, signal_1799}), .a ({signal_2960, signal_1798}), .clk (clk), .r (Fresh[737]), .c ({signal_3035, signal_1859}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1733 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2962, signal_1800}), .a ({signal_2963, signal_1801}), .clk (clk), .r (Fresh[738]), .c ({signal_3036, signal_1860}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1734 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2963, signal_1801}), .a ({signal_2962, signal_1800}), .clk (clk), .r (Fresh[739]), .c ({signal_3037, signal_1861}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1737 ( .s ({signal_2043, signal_1146}), .b ({signal_2976, signal_1813}), .a ({signal_2975, signal_1812}), .clk (clk), .r (Fresh[740]), .c ({signal_3041, signal_838}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1738 ( .s ({signal_2055, signal_1142}), .b ({signal_2978, signal_1815}), .a ({signal_2977, signal_1814}), .clk (clk), .r (Fresh[741]), .c ({signal_3042, signal_834}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1739 ( .s ({signal_2067, signal_1138}), .b ({signal_2980, signal_1817}), .a ({signal_2979, signal_1816}), .clk (clk), .r (Fresh[742]), .c ({signal_3043, signal_830}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1741 ( .s ({signal_2007, signal_1158}), .b ({signal_2984, signal_1821}), .a ({signal_2983, signal_1820}), .clk (clk), .r (Fresh[743]), .c ({signal_3045, signal_822}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1742 ( .s ({signal_2019, signal_1154}), .b ({signal_2986, signal_1823}), .a ({signal_2985, signal_1822}), .clk (clk), .r (Fresh[744]), .c ({signal_3046, signal_818}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1743 ( .s ({signal_1995, signal_1162}), .b ({signal_2988, signal_1825}), .a ({signal_2987, signal_1824}), .clk (clk), .r (Fresh[745]), .c ({signal_3047, signal_810}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1744 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2975, signal_1812}), .a ({signal_2976, signal_1813}), .clk (clk), .r (Fresh[746]), .c ({signal_3048, signal_1864}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1745 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2976, signal_1813}), .a ({signal_2975, signal_1812}), .clk (clk), .r (Fresh[747]), .c ({signal_3049, signal_1865}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1746 ( .s ({Ciphertext_s1[15], Ciphertext_s0[15]}), .b ({signal_2975, signal_1812}), .a ({signal_2976, signal_1813}), .clk (clk), .r (Fresh[748]), .c ({signal_3050, signal_1866}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1747 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2976, signal_1813}), .a ({signal_2975, signal_1812}), .clk (clk), .r (Fresh[749]), .c ({signal_3051, signal_1867}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1748 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2977, signal_1814}), .a ({signal_2978, signal_1815}), .clk (clk), .r (Fresh[750]), .c ({signal_3052, signal_1868}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1749 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2978, signal_1815}), .a ({signal_2977, signal_1814}), .clk (clk), .r (Fresh[751]), .c ({signal_3053, signal_1869}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1750 ( .s ({Ciphertext_s1[3], Ciphertext_s0[3]}), .b ({signal_2977, signal_1814}), .a ({signal_2978, signal_1815}), .clk (clk), .r (Fresh[752]), .c ({signal_3054, signal_1870}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1751 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2978, signal_1815}), .a ({signal_2977, signal_1814}), .clk (clk), .r (Fresh[753]), .c ({signal_3055, signal_1871}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1752 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2979, signal_1816}), .a ({signal_2980, signal_1817}), .clk (clk), .r (Fresh[754]), .c ({signal_3056, signal_1872}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1753 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2980, signal_1817}), .a ({signal_2979, signal_1816}), .clk (clk), .r (Fresh[755]), .c ({signal_3057, signal_1873}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1754 ( .s ({Ciphertext_s1[7], Ciphertext_s0[7]}), .b ({signal_2979, signal_1816}), .a ({signal_2980, signal_1817}), .clk (clk), .r (Fresh[756]), .c ({signal_3058, signal_1874}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1755 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2980, signal_1817}), .a ({signal_2979, signal_1816}), .clk (clk), .r (Fresh[757]), .c ({signal_3059, signal_1875}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1790 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3039, signal_1862}), .a ({signal_2973, signal_1810}), .clk (clk), .r (Fresh[758]), .c ({signal_3123, signal_1904}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1791 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3040, signal_1863}), .a ({signal_2974, signal_1811}), .clk (clk), .r (Fresh[759]), .c ({signal_3124, signal_1905}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1798 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3061, signal_1877}), .a ({signal_3060, signal_1876}), .clk (clk), .r (Fresh[760]), .c ({signal_3132, signal_1912}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1799 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3060, signal_1876}), .a ({signal_3061, signal_1877}), .clk (clk), .r (Fresh[761]), .c ({signal_3133, signal_1913}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1800 ( .s ({signal_2076, signal_1135}), .b ({signal_3063, signal_1879}), .a ({signal_3062, signal_1878}), .clk (clk), .r (Fresh[762]), .c ({signal_3134, signal_1914}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1801 ( .s ({signal_2076, signal_1135}), .b ({signal_3062, signal_1878}), .a ({signal_3063, signal_1879}), .clk (clk), .r (Fresh[763]), .c ({signal_3135, signal_1915}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1802 ( .s ({signal_2028, signal_1151}), .b ({signal_3065, signal_1881}), .a ({signal_3064, signal_1880}), .clk (clk), .r (Fresh[764]), .c ({signal_3136, signal_1916}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1803 ( .s ({signal_2028, signal_1151}), .b ({signal_3064, signal_1880}), .a ({signal_3065, signal_1881}), .clk (clk), .r (Fresh[765]), .c ({signal_3137, signal_1917}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1804 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_3062, signal_1878}), .a ({signal_3063, signal_1879}), .clk (clk), .r (Fresh[766]), .c ({signal_3138, signal_1918}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1805 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_3063, signal_1879}), .a ({signal_3062, signal_1878}), .clk (clk), .r (Fresh[767]), .c ({signal_3139, signal_1919}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1806 ( .s ({signal_2079, signal_1134}), .b ({signal_3067, signal_1883}), .a ({signal_3066, signal_1882}), .clk (clk), .r (Fresh[768]), .c ({signal_3140, signal_1920}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1807 ( .s ({signal_2079, signal_1134}), .b ({signal_3066, signal_1882}), .a ({signal_3067, signal_1883}), .clk (clk), .r (Fresh[769]), .c ({signal_3141, signal_1921}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1808 ( .s ({signal_2031, signal_1150}), .b ({signal_3069, signal_1885}), .a ({signal_3068, signal_1884}), .clk (clk), .r (Fresh[770]), .c ({signal_3142, signal_1922}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1809 ( .s ({signal_2031, signal_1150}), .b ({signal_3068, signal_1884}), .a ({signal_3069, signal_1885}), .clk (clk), .r (Fresh[771]), .c ({signal_3143, signal_1923}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1810 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3066, signal_1882}), .a ({signal_3067, signal_1883}), .clk (clk), .r (Fresh[772]), .c ({signal_3144, signal_1924}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1811 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_3067, signal_1883}), .a ({signal_3066, signal_1882}), .clk (clk), .r (Fresh[773]), .c ({signal_3145, signal_1925}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1812 ( .s ({Ciphertext_s1[11], Ciphertext_s0[11]}), .b ({signal_3066, signal_1882}), .a ({signal_3067, signal_1883}), .clk (clk), .r (Fresh[774]), .c ({signal_3146, signal_1926}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1813 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3067, signal_1883}), .a ({signal_3066, signal_1882}), .clk (clk), .r (Fresh[775]), .c ({signal_3147, signal_1927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1842 ( .s (signal_1028), .b ({signal_3135, signal_1915}), .a ({signal_3134, signal_1914}), .c ({signal_3188, signal_827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1843 ( .s (signal_940), .b ({signal_3137, signal_1917}), .a ({signal_3136, signal_1916}), .c ({signal_3189, signal_815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1850 ( .s (signal_943), .b ({signal_3141, signal_1921}), .a ({signal_3140, signal_1920}), .c ({signal_3196, signal_826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1851 ( .s (signal_939), .b ({signal_3143, signal_1923}), .a ({signal_3142, signal_1922}), .c ({signal_3197, signal_814}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (rst), .b ({signal_3098, signal_789}), .a ({Plaintext_s1[50], Plaintext_s0[50]}), .c ({signal_3149, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (rst), .b ({signal_3101, signal_788}), .a ({Plaintext_s1[51], Plaintext_s0[51]}), .c ({signal_3151, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (rst), .b ({signal_3099, signal_785}), .a ({Plaintext_s1[54], Plaintext_s0[54]}), .c ({signal_3153, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (rst), .b ({signal_3102, signal_784}), .a ({Plaintext_s1[55], Plaintext_s0[55]}), .c ({signal_3155, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (rst), .b ({signal_3100, signal_781}), .a ({Plaintext_s1[58], Plaintext_s0[58]}), .c ({signal_3157, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (rst), .b ({signal_3103, signal_780}), .a ({Plaintext_s1[59], Plaintext_s0[59]}), .c ({signal_3159, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (rst), .b ({signal_3214, signal_777}), .a ({Plaintext_s1[62], Plaintext_s0[62]}), .c ({signal_3231, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (rst), .b ({signal_3221, signal_776}), .a ({Plaintext_s1[63], Plaintext_s0[63]}), .c ({signal_3233, signal_840}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1766 ( .s ({signal_2046, signal_1145}), .b ({signal_3009, signal_1845}), .a ({signal_3008, signal_1844}), .clk (clk), .r (Fresh[776]), .c ({signal_3098, signal_789}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1767 ( .s ({signal_2058, signal_1141}), .b ({signal_3012, signal_1847}), .a ({signal_3011, signal_1846}), .clk (clk), .r (Fresh[777]), .c ({signal_3099, signal_785}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1768 ( .s ({signal_2070, signal_1137}), .b ({signal_3015, signal_1849}), .a ({signal_3014, signal_1848}), .clk (clk), .r (Fresh[778]), .c ({signal_3100, signal_781}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1769 ( .s ({signal_2049, signal_1144}), .b ({signal_3018, signal_1851}), .a ({signal_3017, signal_1850}), .clk (clk), .r (Fresh[779]), .c ({signal_3101, signal_788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1770 ( .s ({signal_2061, signal_1140}), .b ({signal_3021, signal_1853}), .a ({signal_3020, signal_1852}), .clk (clk), .r (Fresh[780]), .c ({signal_3102, signal_784}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1771 ( .s ({signal_2073, signal_1136}), .b ({signal_3024, signal_1855}), .a ({signal_3023, signal_1854}), .clk (clk), .r (Fresh[781]), .c ({signal_3103, signal_780}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1772 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3032, signal_1856}), .a ({signal_2959, signal_1797}), .clk (clk), .r (Fresh[782]), .c ({signal_3104, signal_1886}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1773 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2959, signal_1797}), .a ({signal_3032, signal_1856}), .clk (clk), .r (Fresh[783]), .c ({signal_3105, signal_1887}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1774 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3032, signal_1856}), .a ({signal_3033, signal_1857}), .clk (clk), .r (Fresh[784]), .c ({signal_3106, signal_1888}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1775 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3033, signal_1857}), .a ({signal_2958, signal_1796}), .clk (clk), .r (Fresh[785]), .c ({signal_3107, signal_1889}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1776 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_2958, signal_1796}), .a ({signal_3033, signal_1857}), .clk (clk), .r (Fresh[786]), .c ({signal_3108, signal_1890}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1777 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3033, signal_1857}), .a ({signal_3032, signal_1856}), .clk (clk), .r (Fresh[787]), .c ({signal_3109, signal_1891}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1778 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3034, signal_1858}), .a ({signal_2961, signal_1799}), .clk (clk), .r (Fresh[788]), .c ({signal_3110, signal_1892}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1779 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2961, signal_1799}), .a ({signal_3034, signal_1858}), .clk (clk), .r (Fresh[789]), .c ({signal_3111, signal_1893}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1780 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3034, signal_1858}), .a ({signal_3035, signal_1859}), .clk (clk), .r (Fresh[790]), .c ({signal_3112, signal_1894}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1781 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3035, signal_1859}), .a ({signal_2960, signal_1798}), .clk (clk), .r (Fresh[791]), .c ({signal_3113, signal_1895}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1782 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_2960, signal_1798}), .a ({signal_3035, signal_1859}), .clk (clk), .r (Fresh[792]), .c ({signal_3114, signal_1896}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1783 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3035, signal_1859}), .a ({signal_3034, signal_1858}), .clk (clk), .r (Fresh[793]), .c ({signal_3115, signal_1897}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1784 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3036, signal_1860}), .a ({signal_2963, signal_1801}), .clk (clk), .r (Fresh[794]), .c ({signal_3116, signal_1898}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1785 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2963, signal_1801}), .a ({signal_3036, signal_1860}), .clk (clk), .r (Fresh[795]), .c ({signal_3117, signal_1899}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1786 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3036, signal_1860}), .a ({signal_3037, signal_1861}), .clk (clk), .r (Fresh[796]), .c ({signal_3118, signal_1900}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1787 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3037, signal_1861}), .a ({signal_2962, signal_1800}), .clk (clk), .r (Fresh[797]), .c ({signal_3119, signal_1901}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1788 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_2962, signal_1800}), .a ({signal_3037, signal_1861}), .clk (clk), .r (Fresh[798]), .c ({signal_3120, signal_1902}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1789 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3037, signal_1861}), .a ({signal_3036, signal_1860}), .clk (clk), .r (Fresh[799]), .c ({signal_3121, signal_1903}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1792 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3049, signal_1865}), .a ({signal_2976, signal_1813}), .clk (clk), .r (Fresh[800]), .c ({signal_3125, signal_1906}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1793 ( .s ({Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({signal_3050, signal_1866}), .a ({signal_2975, signal_1812}), .clk (clk), .r (Fresh[801]), .c ({signal_3126, signal_1907}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1794 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3053, signal_1869}), .a ({signal_2978, signal_1815}), .clk (clk), .r (Fresh[802]), .c ({signal_3127, signal_1908}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1795 ( .s ({Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({signal_3054, signal_1870}), .a ({signal_2977, signal_1814}), .clk (clk), .r (Fresh[803]), .c ({signal_3128, signal_1909}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1796 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3057, signal_1873}), .a ({signal_2980, signal_1817}), .clk (clk), .r (Fresh[804]), .c ({signal_3129, signal_1910}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1797 ( .s ({Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({signal_3058, signal_1874}), .a ({signal_2979, signal_1816}), .clk (clk), .r (Fresh[805]), .c ({signal_3130, signal_1911}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1826 ( .s ({signal_2082, signal_1133}), .b ({signal_3124, signal_1905}), .a ({signal_3123, signal_1904}), .clk (clk), .r (Fresh[806]), .c ({signal_3172, signal_1940}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1827 ( .s ({signal_2082, signal_1133}), .b ({signal_3123, signal_1904}), .a ({signal_3124, signal_1905}), .clk (clk), .r (Fresh[807]), .c ({signal_3173, signal_1941}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1840 ( .s ({signal_2085, signal_1132}), .b ({signal_3133, signal_1913}), .a ({signal_3132, signal_1912}), .clk (clk), .r (Fresh[808]), .c ({signal_3186, signal_1954}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1841 ( .s ({signal_2085, signal_1132}), .b ({signal_3132, signal_1912}), .a ({signal_3133, signal_1913}), .clk (clk), .r (Fresh[809]), .c ({signal_3187, signal_1955}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1844 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3138, signal_1918}), .a ({signal_3063, signal_1879}), .clk (clk), .r (Fresh[810]), .c ({signal_3190, signal_1956}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1845 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3063, signal_1879}), .a ({signal_3138, signal_1918}), .clk (clk), .r (Fresh[811]), .c ({signal_3191, signal_1957}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1846 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3138, signal_1918}), .a ({signal_3139, signal_1919}), .clk (clk), .r (Fresh[812]), .c ({signal_3192, signal_1958}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1847 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3139, signal_1919}), .a ({signal_3062, signal_1878}), .clk (clk), .r (Fresh[813]), .c ({signal_3193, signal_1959}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1848 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3062, signal_1878}), .a ({signal_3139, signal_1919}), .clk (clk), .r (Fresh[814]), .c ({signal_3194, signal_1960}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1849 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3139, signal_1919}), .a ({signal_3138, signal_1918}), .clk (clk), .r (Fresh[815]), .c ({signal_3195, signal_1961}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1852 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3145, signal_1925}), .a ({signal_3067, signal_1883}), .clk (clk), .r (Fresh[816]), .c ({signal_3198, signal_1962}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1853 ( .s ({Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({signal_3146, signal_1926}), .a ({signal_3066, signal_1882}), .clk (clk), .r (Fresh[817]), .c ({signal_3199, signal_1963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1860 ( .s (signal_1026), .b ({signal_3173, signal_1941}), .a ({signal_3172, signal_1940}), .c ({signal_3214, signal_777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1867 ( .s (signal_1025), .b ({signal_3187, signal_1955}), .a ({signal_3186, signal_1954}), .c ({signal_3221, signal_776}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1814 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_2958, signal_1796}), .a ({signal_3104, signal_1886}), .clk (clk), .r (Fresh[818]), .c ({signal_3160, signal_1928}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1815 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3106, signal_1888}), .a ({signal_3105, signal_1887}), .clk (clk), .r (Fresh[819]), .c ({signal_3161, signal_1929}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1816 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_2959, signal_1797}), .a ({signal_3107, signal_1889}), .clk (clk), .r (Fresh[820]), .c ({signal_3162, signal_1930}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1817 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3109, signal_1891}), .a ({signal_3108, signal_1890}), .clk (clk), .r (Fresh[821]), .c ({signal_3163, signal_1931}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1818 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_2960, signal_1798}), .a ({signal_3110, signal_1892}), .clk (clk), .r (Fresh[822]), .c ({signal_3164, signal_1932}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1819 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3112, signal_1894}), .a ({signal_3111, signal_1893}), .clk (clk), .r (Fresh[823]), .c ({signal_3165, signal_1933}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1820 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_2961, signal_1799}), .a ({signal_3113, signal_1895}), .clk (clk), .r (Fresh[824]), .c ({signal_3166, signal_1934}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1821 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3115, signal_1897}), .a ({signal_3114, signal_1896}), .clk (clk), .r (Fresh[825]), .c ({signal_3167, signal_1935}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1822 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_2962, signal_1800}), .a ({signal_3116, signal_1898}), .clk (clk), .r (Fresh[826]), .c ({signal_3168, signal_1936}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1823 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3118, signal_1900}), .a ({signal_3117, signal_1899}), .clk (clk), .r (Fresh[827]), .c ({signal_3169, signal_1937}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1824 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_2963, signal_1801}), .a ({signal_3119, signal_1901}), .clk (clk), .r (Fresh[828]), .c ({signal_3170, signal_1938}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1825 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3121, signal_1903}), .a ({signal_3120, signal_1902}), .clk (clk), .r (Fresh[829]), .c ({signal_3171, signal_1939}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1828 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3125, signal_1906}), .a ({signal_3048, signal_1864}), .clk (clk), .r (Fresh[830]), .c ({signal_3174, signal_1942}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1829 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3126, signal_1907}), .a ({signal_3048, signal_1864}), .clk (clk), .r (Fresh[831]), .c ({signal_3175, signal_1943}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1830 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3126, signal_1907}), .a ({signal_3051, signal_1867}), .clk (clk), .r (Fresh[832]), .c ({signal_3176, signal_1944}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1831 ( .s ({Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({signal_3125, signal_1906}), .a ({signal_3051, signal_1867}), .clk (clk), .r (Fresh[833]), .c ({signal_3177, signal_1945}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1832 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3127, signal_1908}), .a ({signal_3052, signal_1868}), .clk (clk), .r (Fresh[834]), .c ({signal_3178, signal_1946}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1833 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3128, signal_1909}), .a ({signal_3052, signal_1868}), .clk (clk), .r (Fresh[835]), .c ({signal_3179, signal_1947}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1834 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3128, signal_1909}), .a ({signal_3055, signal_1871}), .clk (clk), .r (Fresh[836]), .c ({signal_3180, signal_1948}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1835 ( .s ({Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({signal_3127, signal_1908}), .a ({signal_3055, signal_1871}), .clk (clk), .r (Fresh[837]), .c ({signal_3181, signal_1949}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1836 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3129, signal_1910}), .a ({signal_3056, signal_1872}), .clk (clk), .r (Fresh[838]), .c ({signal_3182, signal_1950}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1837 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3130, signal_1911}), .a ({signal_3056, signal_1872}), .clk (clk), .r (Fresh[839]), .c ({signal_3183, signal_1951}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1838 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3130, signal_1911}), .a ({signal_3059, signal_1875}), .clk (clk), .r (Fresh[840]), .c ({signal_3184, signal_1952}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1839 ( .s ({Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({signal_3129, signal_1910}), .a ({signal_3059, signal_1875}), .clk (clk), .r (Fresh[841]), .c ({signal_3185, signal_1953}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1868 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3062, signal_1878}), .a ({signal_3190, signal_1956}), .clk (clk), .r (Fresh[842]), .c ({signal_3222, signal_1976}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1869 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3192, signal_1958}), .a ({signal_3191, signal_1957}), .clk (clk), .r (Fresh[843]), .c ({signal_3223, signal_1977}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1870 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3063, signal_1879}), .a ({signal_3193, signal_1959}), .clk (clk), .r (Fresh[844]), .c ({signal_3224, signal_1978}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1871 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3195, signal_1961}), .a ({signal_3194, signal_1960}), .clk (clk), .r (Fresh[845]), .c ({signal_3225, signal_1979}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1872 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3198, signal_1962}), .a ({signal_3144, signal_1924}), .clk (clk), .r (Fresh[846]), .c ({signal_3226, signal_1980}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1873 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3199, signal_1963}), .a ({signal_3144, signal_1924}), .clk (clk), .r (Fresh[847]), .c ({signal_3227, signal_1981}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1874 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3199, signal_1963}), .a ({signal_3147, signal_1927}), .clk (clk), .r (Fresh[848]), .c ({signal_3228, signal_1982}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1875 ( .s ({Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({signal_3198, signal_1962}), .a ({signal_3147, signal_1927}), .clk (clk), .r (Fresh[849]), .c ({signal_3229, signal_1983}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1854 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_3161, signal_1929}), .a ({signal_3160, signal_1928}), .clk (clk), .r (Fresh[850]), .c ({signal_3208, signal_1964}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1855 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_3163, signal_1931}), .a ({signal_3162, signal_1930}), .clk (clk), .r (Fresh[851]), .c ({signal_3209, signal_1965}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1856 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_3165, signal_1933}), .a ({signal_3164, signal_1932}), .clk (clk), .r (Fresh[852]), .c ({signal_3210, signal_1966}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1857 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_3167, signal_1935}), .a ({signal_3166, signal_1934}), .clk (clk), .r (Fresh[853]), .c ({signal_3211, signal_1967}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1858 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_3169, signal_1937}), .a ({signal_3168, signal_1936}), .clk (clk), .r (Fresh[854]), .c ({signal_3212, signal_1968}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1859 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_3171, signal_1939}), .a ({signal_3170, signal_1938}), .clk (clk), .r (Fresh[855]), .c ({signal_3213, signal_1969}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1861 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_3175, signal_1943}), .a ({signal_3174, signal_1942}), .clk (clk), .r (Fresh[856]), .c ({signal_3215, signal_1970}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1862 ( .s ({Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({signal_3177, signal_1945}), .a ({signal_3176, signal_1944}), .clk (clk), .r (Fresh[857]), .c ({signal_3216, signal_1971}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1863 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_3179, signal_1947}), .a ({signal_3178, signal_1946}), .clk (clk), .r (Fresh[858]), .c ({signal_3217, signal_1972}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1864 ( .s ({Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({signal_3181, signal_1949}), .a ({signal_3180, signal_1948}), .clk (clk), .r (Fresh[859]), .c ({signal_3218, signal_1973}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1865 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_3183, signal_1951}), .a ({signal_3182, signal_1950}), .clk (clk), .r (Fresh[860]), .c ({signal_3219, signal_1974}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1866 ( .s ({Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({signal_3185, signal_1953}), .a ({signal_3184, signal_1952}), .clk (clk), .r (Fresh[861]), .c ({signal_3220, signal_1975}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1882 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3223, signal_1977}), .a ({signal_3222, signal_1976}), .clk (clk), .r (Fresh[862]), .c ({signal_3240, signal_1984}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1883 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3225, signal_1979}), .a ({signal_3224, signal_1978}), .clk (clk), .r (Fresh[863]), .c ({signal_3241, signal_1985}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1884 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3227, signal_1981}), .a ({signal_3226, signal_1980}), .clk (clk), .r (Fresh[864]), .c ({signal_3242, signal_1986}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1885 ( .s ({Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({signal_3229, signal_1983}), .a ({signal_3228, signal_1982}), .clk (clk), .r (Fresh[865]), .c ({signal_3243, signal_1987}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (rst), .b ({signal_3234, signal_791}), .a ({Plaintext_s1[48], Plaintext_s0[48]}), .c ({signal_3245, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (rst), .b ({signal_3237, signal_790}), .a ({Plaintext_s1[49], Plaintext_s0[49]}), .c ({signal_3247, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (rst), .b ({signal_3235, signal_787}), .a ({Plaintext_s1[52], Plaintext_s0[52]}), .c ({signal_3249, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (rst), .b ({signal_3238, signal_786}), .a ({Plaintext_s1[53], Plaintext_s0[53]}), .c ({signal_3251, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (rst), .b ({signal_3236, signal_783}), .a ({Plaintext_s1[56], Plaintext_s0[56]}), .c ({signal_3253, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (rst), .b ({signal_3239, signal_782}), .a ({Plaintext_s1[57], Plaintext_s0[57]}), .c ({signal_3255, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (rst), .b ({signal_3260, signal_779}), .a ({Plaintext_s1[60], Plaintext_s0[60]}), .c ({signal_3263, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (rst), .b ({signal_3261, signal_778}), .a ({Plaintext_s1[61], Plaintext_s0[61]}), .c ({signal_3265, signal_842}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1876 ( .s ({signal_2040, signal_1147}), .b ({signal_3209, signal_1965}), .a ({signal_3208, signal_1964}), .clk (clk), .r (Fresh[866]), .c ({signal_3234, signal_791}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1877 ( .s ({signal_2052, signal_1143}), .b ({signal_3211, signal_1967}), .a ({signal_3210, signal_1966}), .clk (clk), .r (Fresh[867]), .c ({signal_3235, signal_787}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1878 ( .s ({signal_2064, signal_1139}), .b ({signal_3213, signal_1969}), .a ({signal_3212, signal_1968}), .clk (clk), .r (Fresh[868]), .c ({signal_3236, signal_783}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1879 ( .s ({signal_2043, signal_1146}), .b ({signal_3216, signal_1971}), .a ({signal_3215, signal_1970}), .clk (clk), .r (Fresh[869]), .c ({signal_3237, signal_790}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1880 ( .s ({signal_2055, signal_1142}), .b ({signal_3218, signal_1973}), .a ({signal_3217, signal_1972}), .clk (clk), .r (Fresh[870]), .c ({signal_3238, signal_786}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1881 ( .s ({signal_2067, signal_1138}), .b ({signal_3220, signal_1975}), .a ({signal_3219, signal_1974}), .clk (clk), .r (Fresh[871]), .c ({signal_3239, signal_782}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1886 ( .s ({signal_2076, signal_1135}), .b ({signal_3241, signal_1985}), .a ({signal_3240, signal_1984}), .clk (clk), .r (Fresh[872]), .c ({signal_3256, signal_1988}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1887 ( .s ({signal_2076, signal_1135}), .b ({signal_3240, signal_1984}), .a ({signal_3241, signal_1985}), .clk (clk), .r (Fresh[873]), .c ({signal_3257, signal_1989}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1888 ( .s ({signal_2079, signal_1134}), .b ({signal_3243, signal_1987}), .a ({signal_3242, signal_1986}), .clk (clk), .r (Fresh[874]), .c ({signal_3258, signal_1990}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1889 ( .s ({signal_2079, signal_1134}), .b ({signal_3242, signal_1986}), .a ({signal_3243, signal_1987}), .clk (clk), .r (Fresh[875]), .c ({signal_3259, signal_1991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1890 ( .s (signal_1028), .b ({signal_3257, signal_1989}), .a ({signal_3256, signal_1988}), .c ({signal_3260, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_1891 ( .s (signal_943), .b ({signal_3259, signal_1991}), .a ({signal_3258, signal_1990}), .c ({signal_3261, signal_778}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_65 ( .clk (signal_4142), .D ({signal_3233, signal_840}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_67 ( .clk (signal_4142), .D ({signal_3231, signal_841}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_69 ( .clk (signal_4142), .D ({signal_3265, signal_842}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_71 ( .clk (signal_4142), .D ({signal_3263, signal_843}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_73 ( .clk (signal_4142), .D ({signal_3159, signal_844}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_75 ( .clk (signal_4142), .D ({signal_3157, signal_845}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_77 ( .clk (signal_4142), .D ({signal_3255, signal_846}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_79 ( .clk (signal_4142), .D ({signal_3253, signal_847}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_81 ( .clk (signal_4142), .D ({signal_3155, signal_848}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_83 ( .clk (signal_4142), .D ({signal_3153, signal_849}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_85 ( .clk (signal_4142), .D ({signal_3251, signal_850}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_87 ( .clk (signal_4142), .D ({signal_3249, signal_851}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_89 ( .clk (signal_4142), .D ({signal_3151, signal_852}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_91 ( .clk (signal_4142), .D ({signal_3149, signal_853}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_93 ( .clk (signal_4142), .D ({signal_3247, signal_854}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_95 ( .clk (signal_4142), .D ({signal_3245, signal_855}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_97 ( .clk (signal_4142), .D ({signal_2693, signal_856}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_99 ( .clk (signal_4142), .D ({signal_2691, signal_857}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_101 ( .clk (signal_4142), .D ({signal_2817, signal_858}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_103 ( .clk (signal_4142), .D ({signal_2815, signal_859}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_105 ( .clk (signal_4142), .D ({signal_2689, signal_860}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_107 ( .clk (signal_4142), .D ({signal_2687, signal_861}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_109 ( .clk (signal_4142), .D ({signal_2813, signal_862}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_111 ( .clk (signal_4142), .D ({signal_2811, signal_863}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_113 ( .clk (signal_4142), .D ({signal_2685, signal_864}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_115 ( .clk (signal_4142), .D ({signal_2683, signal_865}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_117 ( .clk (signal_4142), .D ({signal_2809, signal_866}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_119 ( .clk (signal_4142), .D ({signal_2807, signal_867}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_121 ( .clk (signal_4142), .D ({signal_2681, signal_868}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_123 ( .clk (signal_4142), .D ({signal_2679, signal_869}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_125 ( .clk (signal_4142), .D ({signal_2805, signal_870}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_127 ( .clk (signal_4142), .D ({signal_2803, signal_871}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_129 ( .clk (signal_4142), .D ({signal_2942, signal_872}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_131 ( .clk (signal_4142), .D ({signal_2940, signal_873}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_133 ( .clk (signal_4142), .D ({signal_3097, signal_874}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_135 ( .clk (signal_4142), .D ({signal_3095, signal_875}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_137 ( .clk (signal_4142), .D ({signal_2938, signal_876}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_139 ( .clk (signal_4142), .D ({signal_2936, signal_877}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_141 ( .clk (signal_4142), .D ({signal_3207, signal_878}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_143 ( .clk (signal_4142), .D ({signal_3205, signal_879}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_145 ( .clk (signal_4142), .D ({signal_2934, signal_880}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_147 ( .clk (signal_4142), .D ({signal_2932, signal_881}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_149 ( .clk (signal_4142), .D ({signal_3093, signal_882}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_151 ( .clk (signal_4142), .D ({signal_3091, signal_883}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_153 ( .clk (signal_4142), .D ({signal_2930, signal_884}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_155 ( .clk (signal_4142), .D ({signal_2928, signal_885}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_157 ( .clk (signal_4142), .D ({signal_3089, signal_886}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_159 ( .clk (signal_4142), .D ({signal_3087, signal_887}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_161 ( .clk (signal_4142), .D ({signal_3085, signal_888}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_163 ( .clk (signal_4142), .D ({signal_3083, signal_889}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_165 ( .clk (signal_4142), .D ({signal_3203, signal_890}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_167 ( .clk (signal_4142), .D ({signal_3201, signal_891}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_169 ( .clk (signal_4142), .D ({signal_2926, signal_892}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_171 ( .clk (signal_4142), .D ({signal_2924, signal_893}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_173 ( .clk (signal_4142), .D ({signal_3081, signal_894}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_175 ( .clk (signal_4142), .D ({signal_3079, signal_895}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_177 ( .clk (signal_4142), .D ({signal_2922, signal_896}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_179 ( .clk (signal_4142), .D ({signal_2920, signal_897}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_181 ( .clk (signal_4142), .D ({signal_3077, signal_898}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_183 ( .clk (signal_4142), .D ({signal_3075, signal_899}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_185 ( .clk (signal_4142), .D ({signal_2918, signal_900}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_187 ( .clk (signal_4142), .D ({signal_2916, signal_901}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_189 ( .clk (signal_4142), .D ({signal_3073, signal_902}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_191 ( .clk (signal_4142), .D ({signal_3071, signal_903}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_834 ( .clk (signal_4142), .D ({signal_2183, signal_1036}), .Q ({signal_2085, signal_1132}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_836 ( .clk (signal_4142), .D ({signal_2180, signal_1037}), .Q ({signal_2082, signal_1133}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_838 ( .clk (signal_4142), .D ({signal_2177, signal_1038}), .Q ({signal_2079, signal_1134}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_840 ( .clk (signal_4142), .D ({signal_2174, signal_1039}), .Q ({signal_2076, signal_1135}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_842 ( .clk (signal_4142), .D ({signal_2171, signal_1040}), .Q ({signal_2073, signal_1136}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_844 ( .clk (signal_4142), .D ({signal_2168, signal_1041}), .Q ({signal_2070, signal_1137}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_846 ( .clk (signal_4142), .D ({signal_2165, signal_1042}), .Q ({signal_2067, signal_1138}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_848 ( .clk (signal_4142), .D ({signal_2162, signal_1043}), .Q ({signal_2064, signal_1139}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_850 ( .clk (signal_4142), .D ({signal_2159, signal_1044}), .Q ({signal_2061, signal_1140}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_852 ( .clk (signal_4142), .D ({signal_2156, signal_1045}), .Q ({signal_2058, signal_1141}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_854 ( .clk (signal_4142), .D ({signal_2153, signal_1046}), .Q ({signal_2055, signal_1142}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_856 ( .clk (signal_4142), .D ({signal_2150, signal_1047}), .Q ({signal_2052, signal_1143}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_858 ( .clk (signal_4142), .D ({signal_2147, signal_1048}), .Q ({signal_2049, signal_1144}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_860 ( .clk (signal_4142), .D ({signal_2144, signal_1049}), .Q ({signal_2046, signal_1145}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_862 ( .clk (signal_4142), .D ({signal_2141, signal_1050}), .Q ({signal_2043, signal_1146}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_864 ( .clk (signal_4142), .D ({signal_2138, signal_1051}), .Q ({signal_2040, signal_1147}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_866 ( .clk (signal_4142), .D ({signal_2135, signal_1052}), .Q ({signal_2037, signal_1148}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_868 ( .clk (signal_4142), .D ({signal_2132, signal_1053}), .Q ({signal_2034, signal_1149}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_870 ( .clk (signal_4142), .D ({signal_2129, signal_1054}), .Q ({signal_2031, signal_1150}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_872 ( .clk (signal_4142), .D ({signal_2126, signal_1055}), .Q ({signal_2028, signal_1151}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_874 ( .clk (signal_4142), .D ({signal_2123, signal_1056}), .Q ({signal_2025, signal_1152}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_876 ( .clk (signal_4142), .D ({signal_2120, signal_1057}), .Q ({signal_2022, signal_1153}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_878 ( .clk (signal_4142), .D ({signal_2117, signal_1058}), .Q ({signal_2019, signal_1154}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_880 ( .clk (signal_4142), .D ({signal_2114, signal_1059}), .Q ({signal_2016, signal_1155}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_882 ( .clk (signal_4142), .D ({signal_2111, signal_1060}), .Q ({signal_2013, signal_1156}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_884 ( .clk (signal_4142), .D ({signal_2108, signal_1061}), .Q ({signal_2010, signal_1157}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_886 ( .clk (signal_4142), .D ({signal_2105, signal_1062}), .Q ({signal_2007, signal_1158}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_888 ( .clk (signal_4142), .D ({signal_2102, signal_1063}), .Q ({signal_2004, signal_1159}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_890 ( .clk (signal_4142), .D ({signal_2099, signal_1064}), .Q ({signal_2001, signal_1160}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_892 ( .clk (signal_4142), .D ({signal_2096, signal_1065}), .Q ({signal_1998, signal_1161}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_894 ( .clk (signal_4142), .D ({signal_2093, signal_1066}), .Q ({signal_1995, signal_1162}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_896 ( .clk (signal_4142), .D ({signal_2090, signal_1067}), .Q ({signal_1992, signal_1163}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_898 ( .clk (signal_4142), .D ({signal_2087, signal_1068}), .Q ({signal_2157, signal_1108}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_900 ( .clk (signal_4142), .D ({signal_2084, signal_1069}), .Q ({signal_2154, signal_1109}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_902 ( .clk (signal_4142), .D ({signal_2081, signal_1070}), .Q ({signal_2151, signal_1110}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_904 ( .clk (signal_4142), .D ({signal_2078, signal_1071}), .Q ({signal_2148, signal_1111}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_906 ( .clk (signal_4142), .D ({signal_2075, signal_1072}), .Q ({signal_2181, signal_1100}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_908 ( .clk (signal_4142), .D ({signal_2072, signal_1073}), .Q ({signal_2178, signal_1101}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_910 ( .clk (signal_4142), .D ({signal_2069, signal_1074}), .Q ({signal_2175, signal_1102}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_912 ( .clk (signal_4142), .D ({signal_2066, signal_1075}), .Q ({signal_2172, signal_1103}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_914 ( .clk (signal_4142), .D ({signal_2063, signal_1076}), .Q ({signal_2133, signal_1116}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_916 ( .clk (signal_4142), .D ({signal_2060, signal_1077}), .Q ({signal_2130, signal_1117}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_918 ( .clk (signal_4142), .D ({signal_2057, signal_1078}), .Q ({signal_2127, signal_1118}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_920 ( .clk (signal_4142), .D ({signal_2054, signal_1079}), .Q ({signal_2124, signal_1119}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_922 ( .clk (signal_4142), .D ({signal_2051, signal_1080}), .Q ({signal_2097, signal_1128}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_924 ( .clk (signal_4142), .D ({signal_2048, signal_1081}), .Q ({signal_2094, signal_1129}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_926 ( .clk (signal_4142), .D ({signal_2045, signal_1082}), .Q ({signal_2091, signal_1130}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_928 ( .clk (signal_4142), .D ({signal_2042, signal_1083}), .Q ({signal_2088, signal_1131}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_930 ( .clk (signal_4142), .D ({signal_2039, signal_1084}), .Q ({signal_2109, signal_1124}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_932 ( .clk (signal_4142), .D ({signal_2036, signal_1085}), .Q ({signal_2106, signal_1125}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_934 ( .clk (signal_4142), .D ({signal_2033, signal_1086}), .Q ({signal_2103, signal_1126}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_936 ( .clk (signal_4142), .D ({signal_2030, signal_1087}), .Q ({signal_2100, signal_1127}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_938 ( .clk (signal_4142), .D ({signal_2027, signal_1088}), .Q ({signal_2145, signal_1112}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_940 ( .clk (signal_4142), .D ({signal_2024, signal_1089}), .Q ({signal_2142, signal_1113}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_942 ( .clk (signal_4142), .D ({signal_2021, signal_1090}), .Q ({signal_2139, signal_1114}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_944 ( .clk (signal_4142), .D ({signal_2018, signal_1091}), .Q ({signal_2136, signal_1115}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_946 ( .clk (signal_4142), .D ({signal_2015, signal_1092}), .Q ({signal_2121, signal_1120}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_948 ( .clk (signal_4142), .D ({signal_2012, signal_1093}), .Q ({signal_2118, signal_1121}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_950 ( .clk (signal_4142), .D ({signal_2009, signal_1094}), .Q ({signal_2115, signal_1122}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_952 ( .clk (signal_4142), .D ({signal_2006, signal_1095}), .Q ({signal_2112, signal_1123}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_954 ( .clk (signal_4142), .D ({signal_2003, signal_1096}), .Q ({signal_2169, signal_1104}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_956 ( .clk (signal_4142), .D ({signal_2000, signal_1097}), .Q ({signal_2166, signal_1105}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_958 ( .clk (signal_4142), .D ({signal_1997, signal_1098}), .Q ({signal_2163, signal_1106}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_960 ( .clk (signal_4142), .D ({signal_1994, signal_1099}), .Q ({signal_2160, signal_1107}) ) ;
    DFF_X1 cell_968 ( .CK (signal_4142), .D (signal_1030), .Q (signal_939), .QN () ) ;
    DFF_X1 cell_970 ( .CK (signal_4142), .D (signal_1031), .Q (signal_940), .QN () ) ;
    DFF_X1 cell_972 ( .CK (signal_4142), .D (signal_1032), .Q (signal_1025), .QN () ) ;
    DFF_X1 cell_974 ( .CK (signal_4142), .D (signal_1033), .Q (signal_1026), .QN () ) ;
    DFF_X1 cell_976 ( .CK (signal_4142), .D (signal_1034), .Q (signal_943), .QN () ) ;
    DFF_X1 cell_978 ( .CK (signal_4142), .D (signal_1035), .Q (signal_1028), .QN () ) ;
endmodule
