/* modified netlist. Source: module PRESENT in file /PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module PRESENT_HPC2_ClockGating_d1 (data_in_s0, key_s0, clk, reset, data_in_s1, key_s1, Fresh, data_out_s0, done, data_out_s1, Synch);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [3:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    output Synch ;
    wire selSbox ;
    wire ctrlData_0_ ;
    wire intDone ;
    wire fsm_n15 ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n4 ;
    wire fsm_n2 ;
    wire fsm_n5 ;
    wire fsm_n20 ;
    wire fsm_ps_state_0_ ;
    wire fsm_ps_state_1_ ;
    wire fsm_n21 ;
    wire fsm_n3 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_cnt_rnd_n33 ;
    wire fsm_cnt_rnd_n32 ;
    wire fsm_cnt_rnd_n31 ;
    wire fsm_cnt_rnd_n30 ;
    wire fsm_cnt_rnd_n29 ;
    wire fsm_cnt_rnd_n28 ;
    wire fsm_cnt_rnd_n27 ;
    wire fsm_cnt_rnd_n26 ;
    wire fsm_cnt_rnd_n23 ;
    wire fsm_cnt_rnd_n22 ;
    wire fsm_cnt_rnd_n21 ;
    wire fsm_cnt_rnd_n20 ;
    wire fsm_cnt_rnd_n19 ;
    wire fsm_cnt_rnd_n17 ;
    wire fsm_cnt_rnd_n15 ;
    wire fsm_cnt_rnd_n13 ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n11 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_rnd_n24 ;
    wire fsm_cnt_rnd_n41 ;
    wire fsm_cnt_rnd_n25 ;
    wire fsm_cnt_rnd_n1 ;
    wire fsm_cnt_rnd_n18 ;
    wire fsm_cnt_rnd_n16 ;
    wire fsm_cnt_rnd_n14 ;
    wire fsm_cnt_ser_n10 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n8 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n2 ;
    wire fsm_cnt_ser_n20 ;
    wire fsm_cnt_ser_n28 ;
    wire fsm_cnt_ser_n26 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n1 ;
    wire stateFF_state_n7 ;
    wire stateFF_state_n6 ;
    wire stateFF_state_n5 ;
    wire keyFF_keystate_n8 ;
    wire keyFF_keystate_n7 ;
    wire keyFF_keystate_n6 ;
    wire sboxInst_n3 ;
    wire sboxInst_n2 ;
    wire sboxInst_n1 ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [3:0] stateFF_state_gff_1_s_next_state ;
    wire [3:0] stateFF_state_gff_2_s_next_state ;
    wire [3:0] stateFF_state_gff_3_s_next_state ;
    wire [3:0] stateFF_state_gff_4_s_next_state ;
    wire [3:0] stateFF_state_gff_5_s_next_state ;
    wire [3:0] stateFF_state_gff_6_s_next_state ;
    wire [3:0] stateFF_state_gff_7_s_next_state ;
    wire [3:0] stateFF_state_gff_8_s_next_state ;
    wire [3:0] stateFF_state_gff_9_s_next_state ;
    wire [3:0] stateFF_state_gff_10_s_next_state ;
    wire [3:0] stateFF_state_gff_11_s_next_state ;
    wire [3:0] stateFF_state_gff_12_s_next_state ;
    wire [3:0] stateFF_state_gff_13_s_next_state ;
    wire [3:0] stateFF_state_gff_14_s_next_state ;
    wire [3:0] stateFF_state_gff_15_s_next_state ;
    wire [3:0] stateFF_state_gff_16_s_next_state ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;
    wire [3:0] keyFF_keystate_gff_1_s_next_state ;
    wire [3:0] keyFF_keystate_gff_2_s_next_state ;
    wire [3:0] keyFF_keystate_gff_3_s_next_state ;
    wire [3:0] keyFF_keystate_gff_4_s_next_state ;
    wire [3:0] keyFF_keystate_gff_5_s_next_state ;
    wire [3:0] keyFF_keystate_gff_6_s_next_state ;
    wire [3:0] keyFF_keystate_gff_7_s_next_state ;
    wire [3:0] keyFF_keystate_gff_8_s_next_state ;
    wire [3:0] keyFF_keystate_gff_9_s_next_state ;
    wire [3:0] keyFF_keystate_gff_10_s_next_state ;
    wire [3:0] keyFF_keystate_gff_11_s_next_state ;
    wire [3:0] keyFF_keystate_gff_12_s_next_state ;
    wire [3:0] keyFF_keystate_gff_13_s_next_state ;
    wire [3:0] keyFF_keystate_gff_14_s_next_state ;
    wire [3:0] keyFF_keystate_gff_15_s_next_state ;
    wire [3:0] keyFF_keystate_gff_16_s_next_state ;
    wire [3:0] keyFF_keystate_gff_17_s_next_state ;
    wire [3:0] keyFF_keystate_gff_18_s_next_state ;
    wire [3:0] keyFF_keystate_gff_19_s_next_state ;
    wire [3:0] keyFF_keystate_gff_20_s_next_state ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U9 ( .a ({new_AGEMA_signal_856, roundkey[0]}), .b ({data_out_s1[60], data_out_s0[60]}), .c ({new_AGEMA_signal_858, stateXORroundkey[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U10 ( .a ({new_AGEMA_signal_859, roundkey[1]}), .b ({data_out_s1[61], data_out_s0[61]}), .c ({new_AGEMA_signal_861, stateXORroundkey[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U11 ( .a ({new_AGEMA_signal_862, roundkey[2]}), .b ({data_out_s1[62], data_out_s0[62]}), .c ({new_AGEMA_signal_864, stateXORroundkey[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U12 ( .a ({new_AGEMA_signal_865, roundkey[3]}), .b ({data_out_s1[63], data_out_s0[63]}), .c ({new_AGEMA_signal_867, stateXORroundkey[3]}) ) ;
    NOR2_X1 fsm_U20 ( .A1 (reset), .A2 (fsm_n15), .ZN (fsm_n21) ) ;
    NOR2_X1 fsm_U19 ( .A1 (fsm_n14), .A2 (done), .ZN (fsm_n15) ) ;
    NOR2_X1 fsm_U18 ( .A1 (reset), .A2 (fsm_n13), .ZN (fsm_n20) ) ;
    NOR2_X1 fsm_U17 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n12), .ZN (fsm_n13) ) ;
    NOR2_X1 fsm_U16 ( .A1 (fsm_n11), .A2 (fsm_n10), .ZN (fsm_n12) ) ;
    NAND2_X1 fsm_U15 ( .A1 (counter[3]), .A2 (counter[1]), .ZN (fsm_n10) ) ;
    OR2_X1 fsm_U14 ( .A1 (fsm_n9), .A2 (fsm_n8), .ZN (fsm_n11) ) ;
    NAND2_X1 fsm_U13 ( .A1 (counter[0]), .A2 (counter[4]), .ZN (fsm_n8) ) ;
    NAND2_X1 fsm_U12 ( .A1 (counter[2]), .A2 (fsm_ps_state_0_), .ZN (fsm_n9) ) ;
    NOR2_X1 fsm_U11 ( .A1 (fsm_n3), .A2 (fsm_n5), .ZN (done) ) ;
    AND2_X1 fsm_U10 ( .A1 (fsm_n14), .A2 (fsm_n5), .ZN (fsm_en_countRound) ) ;
    AND2_X1 fsm_U9 ( .A1 (fsm_countSerial[2]), .A2 (fsm_n7), .ZN (fsm_n14) ) ;
    NOR2_X1 fsm_U8 ( .A1 (fsm_n6), .A2 (fsm_n4), .ZN (fsm_n7) ) ;
    NAND2_X1 fsm_U7 ( .A1 (fsm_countSerial[1]), .A2 (fsm_countSerial[0]), .ZN (fsm_n4) ) ;
    NAND2_X1 fsm_U6 ( .A1 (fsm_n3), .A2 (fsm_countSerial[3]), .ZN (fsm_n6) ) ;
    NOR2_X1 fsm_U5 ( .A1 (fsm_ps_state_0_), .A2 (fsm_n5), .ZN (intDone) ) ;
    NOR2_X1 fsm_U4 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n3), .ZN (selSbox) ) ;
    NOR2_X1 fsm_U3 ( .A1 (reset), .A2 (selSbox), .ZN (fsm_rst_countSerial) ) ;
    INV_X1 fsm_U2 ( .A (reset), .ZN (fsm_n2) ) ;
    INV_X1 fsm_U1 ( .A (fsm_rst_countSerial), .ZN (ctrlData_0_) ) ;
    NAND2_X1 fsm_cnt_rnd_U28 ( .A1 (fsm_cnt_rnd_n33), .A2 (fsm_cnt_rnd_n32), .ZN (fsm_cnt_rnd_n41) ) ;
    NAND2_X1 fsm_cnt_rnd_U27 ( .A1 (fsm_cnt_rnd_n31), .A2 (counter[1]), .ZN (fsm_cnt_rnd_n32) ) ;
    NAND2_X1 fsm_cnt_rnd_U26 ( .A1 (fsm_cnt_rnd_n30), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n33) ) ;
    NAND2_X1 fsm_cnt_rnd_U25 ( .A1 (fsm_cnt_rnd_n29), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n30) ) ;
    NAND2_X1 fsm_cnt_rnd_U24 ( .A1 (fsm_cnt_rnd_n28), .A2 (fsm_cnt_rnd_n27), .ZN (fsm_cnt_rnd_n18) ) ;
    NAND2_X1 fsm_cnt_rnd_U23 ( .A1 (fsm_cnt_rnd_n26), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n27) ) ;
    MUX2_X1 fsm_cnt_rnd_U22 ( .S (fsm_cnt_rnd_n5), .A (fsm_cnt_rnd_n23), .B (fsm_cnt_rnd_n22), .Z (fsm_cnt_rnd_n16) ) ;
    NAND2_X1 fsm_cnt_rnd_U21 ( .A1 (fsm_cnt_rnd_n31), .A2 (fsm_cnt_rnd_n21), .ZN (fsm_cnt_rnd_n23) ) ;
    NAND2_X1 fsm_cnt_rnd_U20 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n21) ) ;
    NOR2_X1 fsm_cnt_rnd_U19 ( .A1 (fsm_cnt_rnd_n20), .A2 (fsm_cnt_rnd_n26), .ZN (fsm_cnt_rnd_n31) ) ;
    NOR2_X1 fsm_cnt_rnd_U18 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n6), .ZN (fsm_cnt_rnd_n26) ) ;
    INV_X1 fsm_cnt_rnd_U17 ( .A (fsm_cnt_rnd_n28), .ZN (fsm_cnt_rnd_n20) ) ;
    NAND2_X1 fsm_cnt_rnd_U16 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n28) ) ;
    MUX2_X1 fsm_cnt_rnd_U15 ( .S (counter[4]), .A (fsm_cnt_rnd_n19), .B (fsm_cnt_rnd_n17), .Z (fsm_cnt_rnd_n14) ) ;
    NAND2_X1 fsm_cnt_rnd_U14 ( .A1 (fsm_cnt_rnd_n15), .A2 (fsm_cnt_rnd_n13), .ZN (fsm_cnt_rnd_n17) ) ;
    NAND2_X1 fsm_cnt_rnd_U13 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n25), .ZN (fsm_cnt_rnd_n15) ) ;
    INV_X1 fsm_cnt_rnd_U12 ( .A (fsm_cnt_rnd_n12), .ZN (fsm_cnt_rnd_n29) ) ;
    NOR2_X1 fsm_cnt_rnd_U11 ( .A1 (fsm_cnt_rnd_n25), .A2 (fsm_cnt_rnd_n11), .ZN (fsm_cnt_rnd_n19) ) ;
    INV_X1 fsm_cnt_rnd_U10 ( .A (fsm_cnt_rnd_n10), .ZN (fsm_cnt_rnd_n1) ) ;
    MUX2_X1 fsm_cnt_rnd_U9 ( .S (fsm_cnt_rnd_n25), .A (fsm_cnt_rnd_n13), .B (fsm_cnt_rnd_n11), .Z (fsm_cnt_rnd_n10) ) ;
    NAND2_X1 fsm_cnt_rnd_U8 ( .A1 (counter[2]), .A2 (fsm_cnt_rnd_n22), .ZN (fsm_cnt_rnd_n11) ) ;
    NOR2_X1 fsm_cnt_rnd_U7 ( .A1 (fsm_cnt_rnd_n12), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n22) ) ;
    NAND2_X1 fsm_cnt_rnd_U6 ( .A1 (fsm_en_countRound), .A2 (fsm_n2), .ZN (fsm_cnt_rnd_n12) ) ;
    NAND2_X1 fsm_cnt_rnd_U5 ( .A1 (fsm_n2), .A2 (fsm_cnt_rnd_n8), .ZN (fsm_cnt_rnd_n13) ) ;
    NAND2_X1 fsm_cnt_rnd_U4 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n7), .ZN (fsm_cnt_rnd_n8) ) ;
    NOR2_X1 fsm_cnt_rnd_U3 ( .A1 (fsm_cnt_rnd_n5), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n7) ) ;
    OR2_X1 fsm_cnt_rnd_U2 ( .A1 (fsm_cnt_rnd_n24), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n9) ) ;
    INV_X1 fsm_cnt_rnd_U1 ( .A (fsm_n2), .ZN (fsm_cnt_rnd_n6) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_2__U1 ( .A (counter[2]), .ZN (fsm_cnt_rnd_n5) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_0__U1 ( .A (counter[0]), .ZN (fsm_cnt_rnd_n3) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_3__U1 ( .A (counter[3]), .ZN (fsm_cnt_rnd_n25) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_1__U1 ( .A (fsm_cnt_rnd_n24), .ZN (counter[1]) ) ;
    NOR2_X1 fsm_cnt_ser_U12 ( .A1 (fsm_cnt_ser_n10), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n3) ) ;
    XNOR2_X1 fsm_cnt_ser_U11 ( .A (fsm_n3), .B (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n10) ) ;
    NOR2_X1 fsm_cnt_ser_U10 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n8), .ZN (fsm_cnt_ser_n28) ) ;
    XOR2_X1 fsm_cnt_ser_U9 ( .A (fsm_countSerial[1]), .B (fsm_cnt_ser_n7), .Z (fsm_cnt_ser_n8) ) ;
    NOR2_X1 fsm_cnt_ser_U8 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n6), .ZN (fsm_cnt_ser_n26) ) ;
    XOR2_X1 fsm_cnt_ser_U7 ( .A (fsm_countSerial[3]), .B (fsm_cnt_ser_n5), .Z (fsm_cnt_ser_n6) ) ;
    NAND2_X1 fsm_cnt_ser_U6 ( .A1 (fsm_cnt_ser_n4), .A2 (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n5) ) ;
    NOR2_X1 fsm_cnt_ser_U5 ( .A1 (fsm_cnt_ser_n2), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n1) ) ;
    INV_X1 fsm_cnt_ser_U4 ( .A (fsm_rst_countSerial), .ZN (fsm_cnt_ser_n9) ) ;
    XNOR2_X1 fsm_cnt_ser_U3 ( .A (fsm_cnt_ser_n4), .B (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n2) ) ;
    NOR2_X1 fsm_cnt_ser_U2 ( .A1 (fsm_cnt_ser_n20), .A2 (fsm_cnt_ser_n7), .ZN (fsm_cnt_ser_n4) ) ;
    NAND2_X1 fsm_cnt_ser_U1 ( .A1 (fsm_n3), .A2 (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n7) ) ;
    INV_X1 fsm_cnt_ser_count_reg_reg_1__U1 ( .A (fsm_countSerial[1]), .ZN (fsm_cnt_ser_n20) ) ;
    INV_X1 fsm_ps_state_reg_0__U1 ( .A (fsm_ps_state_0_), .ZN (fsm_n3) ) ;
    INV_X1 fsm_ps_state_reg_1__U1 ( .A (fsm_ps_state_1_), .ZN (fsm_n5) ) ;
    INV_X1 stateFF_state_U3 ( .A (stateFF_state_n7), .ZN (stateFF_state_n6) ) ;
    INV_X1 stateFF_state_U2 ( .A (stateFF_state_n7), .ZN (stateFF_state_n5) ) ;
    INV_X1 stateFF_state_U1 ( .A (ctrlData_0_), .ZN (stateFF_state_n7) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({data_out_s1[0], data_out_s0[0]}), .a ({new_AGEMA_signal_882, stateFF_inputPar[4]}), .c ({new_AGEMA_signal_1299, stateFF_state_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({data_out_s1[1], data_out_s0[1]}), .a ({new_AGEMA_signal_885, stateFF_inputPar[5]}), .c ({new_AGEMA_signal_1300, stateFF_state_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({data_out_s1[2], data_out_s0[2]}), .a ({new_AGEMA_signal_888, stateFF_inputPar[6]}), .c ({new_AGEMA_signal_1301, stateFF_state_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({data_out_s1[3], data_out_s0[3]}), .a ({new_AGEMA_signal_891, stateFF_inputPar[7]}), .c ({new_AGEMA_signal_1302, stateFF_state_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[4], data_out_s0[4]}), .a ({new_AGEMA_signal_894, stateFF_inputPar[8]}), .c ({new_AGEMA_signal_1318, stateFF_state_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[5], data_out_s0[5]}), .a ({new_AGEMA_signal_897, stateFF_inputPar[9]}), .c ({new_AGEMA_signal_1319, stateFF_state_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[6], data_out_s0[6]}), .a ({new_AGEMA_signal_900, stateFF_inputPar[10]}), .c ({new_AGEMA_signal_1320, stateFF_state_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[7], data_out_s0[7]}), .a ({new_AGEMA_signal_903, stateFF_inputPar[11]}), .c ({new_AGEMA_signal_1321, stateFF_state_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[8], data_out_s0[8]}), .a ({new_AGEMA_signal_906, stateFF_inputPar[12]}), .c ({new_AGEMA_signal_1322, stateFF_state_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[9], data_out_s0[9]}), .a ({new_AGEMA_signal_909, stateFF_inputPar[13]}), .c ({new_AGEMA_signal_1323, stateFF_state_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[10], data_out_s0[10]}), .a ({new_AGEMA_signal_912, stateFF_inputPar[14]}), .c ({new_AGEMA_signal_1324, stateFF_state_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[11], data_out_s0[11]}), .a ({new_AGEMA_signal_914, stateFF_inputPar[15]}), .c ({new_AGEMA_signal_1325, stateFF_state_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[12], data_out_s0[12]}), .a ({new_AGEMA_signal_917, stateFF_inputPar[16]}), .c ({new_AGEMA_signal_1326, stateFF_state_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[13], data_out_s0[13]}), .a ({new_AGEMA_signal_920, stateFF_inputPar[17]}), .c ({new_AGEMA_signal_1327, stateFF_state_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[14], data_out_s0[14]}), .a ({new_AGEMA_signal_923, stateFF_inputPar[18]}), .c ({new_AGEMA_signal_1328, stateFF_state_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[15], data_out_s0[15]}), .a ({new_AGEMA_signal_926, stateFF_inputPar[19]}), .c ({new_AGEMA_signal_1329, stateFF_state_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[16], data_out_s0[16]}), .a ({new_AGEMA_signal_929, stateFF_inputPar[20]}), .c ({new_AGEMA_signal_1330, stateFF_state_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[17], data_out_s0[17]}), .a ({new_AGEMA_signal_932, stateFF_inputPar[21]}), .c ({new_AGEMA_signal_1331, stateFF_state_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[18], data_out_s0[18]}), .a ({new_AGEMA_signal_935, stateFF_inputPar[22]}), .c ({new_AGEMA_signal_1332, stateFF_state_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[19], data_out_s0[19]}), .a ({new_AGEMA_signal_938, stateFF_inputPar[23]}), .c ({new_AGEMA_signal_1333, stateFF_state_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[20], data_out_s0[20]}), .a ({new_AGEMA_signal_941, stateFF_inputPar[24]}), .c ({new_AGEMA_signal_1334, stateFF_state_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[21], data_out_s0[21]}), .a ({new_AGEMA_signal_944, stateFF_inputPar[25]}), .c ({new_AGEMA_signal_1335, stateFF_state_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[22], data_out_s0[22]}), .a ({new_AGEMA_signal_947, stateFF_inputPar[26]}), .c ({new_AGEMA_signal_1336, stateFF_state_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[23], data_out_s0[23]}), .a ({new_AGEMA_signal_950, stateFF_inputPar[27]}), .c ({new_AGEMA_signal_1337, stateFF_state_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[24], data_out_s0[24]}), .a ({new_AGEMA_signal_953, stateFF_inputPar[28]}), .c ({new_AGEMA_signal_1338, stateFF_state_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[25], data_out_s0[25]}), .a ({new_AGEMA_signal_956, stateFF_inputPar[29]}), .c ({new_AGEMA_signal_1339, stateFF_state_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[26], data_out_s0[26]}), .a ({new_AGEMA_signal_959, stateFF_inputPar[30]}), .c ({new_AGEMA_signal_1340, stateFF_state_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[27], data_out_s0[27]}), .a ({new_AGEMA_signal_961, stateFF_inputPar[31]}), .c ({new_AGEMA_signal_1341, stateFF_state_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[28], data_out_s0[28]}), .a ({new_AGEMA_signal_964, stateFF_inputPar[32]}), .c ({new_AGEMA_signal_1342, stateFF_state_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[29], data_out_s0[29]}), .a ({new_AGEMA_signal_967, stateFF_inputPar[33]}), .c ({new_AGEMA_signal_1343, stateFF_state_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[30], data_out_s0[30]}), .a ({new_AGEMA_signal_970, stateFF_inputPar[34]}), .c ({new_AGEMA_signal_1344, stateFF_state_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[31], data_out_s0[31]}), .a ({new_AGEMA_signal_973, stateFF_inputPar[35]}), .c ({new_AGEMA_signal_1345, stateFF_state_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[32], data_out_s0[32]}), .a ({new_AGEMA_signal_976, stateFF_inputPar[36]}), .c ({new_AGEMA_signal_1346, stateFF_state_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[33], data_out_s0[33]}), .a ({new_AGEMA_signal_979, stateFF_inputPar[37]}), .c ({new_AGEMA_signal_1347, stateFF_state_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[34], data_out_s0[34]}), .a ({new_AGEMA_signal_982, stateFF_inputPar[38]}), .c ({new_AGEMA_signal_1348, stateFF_state_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[35], data_out_s0[35]}), .a ({new_AGEMA_signal_985, stateFF_inputPar[39]}), .c ({new_AGEMA_signal_1349, stateFF_state_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[36], data_out_s0[36]}), .a ({new_AGEMA_signal_988, stateFF_inputPar[40]}), .c ({new_AGEMA_signal_1350, stateFF_state_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[37], data_out_s0[37]}), .a ({new_AGEMA_signal_991, stateFF_inputPar[41]}), .c ({new_AGEMA_signal_1351, stateFF_state_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[38], data_out_s0[38]}), .a ({new_AGEMA_signal_994, stateFF_inputPar[42]}), .c ({new_AGEMA_signal_1352, stateFF_state_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[39], data_out_s0[39]}), .a ({new_AGEMA_signal_997, stateFF_inputPar[43]}), .c ({new_AGEMA_signal_1353, stateFF_state_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[40], data_out_s0[40]}), .a ({new_AGEMA_signal_1000, stateFF_inputPar[44]}), .c ({new_AGEMA_signal_1354, stateFF_state_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[41], data_out_s0[41]}), .a ({new_AGEMA_signal_1003, stateFF_inputPar[45]}), .c ({new_AGEMA_signal_1355, stateFF_state_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[42], data_out_s0[42]}), .a ({new_AGEMA_signal_1006, stateFF_inputPar[46]}), .c ({new_AGEMA_signal_1356, stateFF_state_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[43], data_out_s0[43]}), .a ({new_AGEMA_signal_1008, stateFF_inputPar[47]}), .c ({new_AGEMA_signal_1357, stateFF_state_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[44], data_out_s0[44]}), .a ({new_AGEMA_signal_1011, stateFF_inputPar[48]}), .c ({new_AGEMA_signal_1358, stateFF_state_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[45], data_out_s0[45]}), .a ({new_AGEMA_signal_1014, stateFF_inputPar[49]}), .c ({new_AGEMA_signal_1359, stateFF_state_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[46], data_out_s0[46]}), .a ({new_AGEMA_signal_1017, stateFF_inputPar[50]}), .c ({new_AGEMA_signal_1360, stateFF_state_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[47], data_out_s0[47]}), .a ({new_AGEMA_signal_1020, stateFF_inputPar[51]}), .c ({new_AGEMA_signal_1361, stateFF_state_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[48], data_out_s0[48]}), .a ({new_AGEMA_signal_1023, stateFF_inputPar[52]}), .c ({new_AGEMA_signal_1362, stateFF_state_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[49], data_out_s0[49]}), .a ({new_AGEMA_signal_1026, stateFF_inputPar[53]}), .c ({new_AGEMA_signal_1363, stateFF_state_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[50], data_out_s0[50]}), .a ({new_AGEMA_signal_1029, stateFF_inputPar[54]}), .c ({new_AGEMA_signal_1364, stateFF_state_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[51], data_out_s0[51]}), .a ({new_AGEMA_signal_1032, stateFF_inputPar[55]}), .c ({new_AGEMA_signal_1365, stateFF_state_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[52], data_out_s0[52]}), .a ({new_AGEMA_signal_1035, stateFF_inputPar[56]}), .c ({new_AGEMA_signal_1366, stateFF_state_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[53], data_out_s0[53]}), .a ({new_AGEMA_signal_1038, stateFF_inputPar[57]}), .c ({new_AGEMA_signal_1367, stateFF_state_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[54], data_out_s0[54]}), .a ({new_AGEMA_signal_1041, stateFF_inputPar[58]}), .c ({new_AGEMA_signal_1368, stateFF_state_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[55], data_out_s0[55]}), .a ({new_AGEMA_signal_1044, stateFF_inputPar[59]}), .c ({new_AGEMA_signal_1369, stateFF_state_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[56], data_out_s0[56]}), .a ({new_AGEMA_signal_1047, stateFF_inputPar[60]}), .c ({new_AGEMA_signal_1370, stateFF_state_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[57], data_out_s0[57]}), .a ({new_AGEMA_signal_1050, stateFF_inputPar[61]}), .c ({new_AGEMA_signal_1371, stateFF_state_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[58], data_out_s0[58]}), .a ({new_AGEMA_signal_1053, stateFF_inputPar[62]}), .c ({new_AGEMA_signal_1372, stateFF_state_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[59], data_out_s0[59]}), .a ({new_AGEMA_signal_1055, stateFF_inputPar[63]}), .c ({new_AGEMA_signal_1373, stateFF_state_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({data_out_s1[0], data_out_s0[0]}), .a ({data_in_s1[0], data_in_s0[0]}), .c ({new_AGEMA_signal_870, stateFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({data_out_s1[4], data_out_s0[4]}), .a ({data_in_s1[1], data_in_s0[1]}), .c ({new_AGEMA_signal_873, stateFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({data_out_s1[8], data_out_s0[8]}), .a ({data_in_s1[2], data_in_s0[2]}), .c ({new_AGEMA_signal_876, stateFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({data_out_s1[12], data_out_s0[12]}), .a ({data_in_s1[3], data_in_s0[3]}), .c ({new_AGEMA_signal_879, stateFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({data_out_s1[16], data_out_s0[16]}), .a ({data_in_s1[4], data_in_s0[4]}), .c ({new_AGEMA_signal_882, stateFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({data_out_s1[20], data_out_s0[20]}), .a ({data_in_s1[5], data_in_s0[5]}), .c ({new_AGEMA_signal_885, stateFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({data_out_s1[24], data_out_s0[24]}), .a ({data_in_s1[6], data_in_s0[6]}), .c ({new_AGEMA_signal_888, stateFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({data_out_s1[28], data_out_s0[28]}), .a ({data_in_s1[7], data_in_s0[7]}), .c ({new_AGEMA_signal_891, stateFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({data_out_s1[32], data_out_s0[32]}), .a ({data_in_s1[8], data_in_s0[8]}), .c ({new_AGEMA_signal_894, stateFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({data_out_s1[36], data_out_s0[36]}), .a ({data_in_s1[9], data_in_s0[9]}), .c ({new_AGEMA_signal_897, stateFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({data_out_s1[40], data_out_s0[40]}), .a ({data_in_s1[10], data_in_s0[10]}), .c ({new_AGEMA_signal_900, stateFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({data_out_s1[44], data_out_s0[44]}), .a ({data_in_s1[11], data_in_s0[11]}), .c ({new_AGEMA_signal_903, stateFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({data_out_s1[48], data_out_s0[48]}), .a ({data_in_s1[12], data_in_s0[12]}), .c ({new_AGEMA_signal_906, stateFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({data_out_s1[52], data_out_s0[52]}), .a ({data_in_s1[13], data_in_s0[13]}), .c ({new_AGEMA_signal_909, stateFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({data_out_s1[56], data_out_s0[56]}), .a ({data_in_s1[14], data_in_s0[14]}), .c ({new_AGEMA_signal_912, stateFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({data_out_s1[60], data_out_s0[60]}), .a ({data_in_s1[15], data_in_s0[15]}), .c ({new_AGEMA_signal_914, stateFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({data_out_s1[1], data_out_s0[1]}), .a ({data_in_s1[16], data_in_s0[16]}), .c ({new_AGEMA_signal_917, stateFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({data_out_s1[5], data_out_s0[5]}), .a ({data_in_s1[17], data_in_s0[17]}), .c ({new_AGEMA_signal_920, stateFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({data_out_s1[9], data_out_s0[9]}), .a ({data_in_s1[18], data_in_s0[18]}), .c ({new_AGEMA_signal_923, stateFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({data_out_s1[13], data_out_s0[13]}), .a ({data_in_s1[19], data_in_s0[19]}), .c ({new_AGEMA_signal_926, stateFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({data_out_s1[17], data_out_s0[17]}), .a ({data_in_s1[20], data_in_s0[20]}), .c ({new_AGEMA_signal_929, stateFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({data_out_s1[21], data_out_s0[21]}), .a ({data_in_s1[21], data_in_s0[21]}), .c ({new_AGEMA_signal_932, stateFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({data_out_s1[25], data_out_s0[25]}), .a ({data_in_s1[22], data_in_s0[22]}), .c ({new_AGEMA_signal_935, stateFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({data_out_s1[29], data_out_s0[29]}), .a ({data_in_s1[23], data_in_s0[23]}), .c ({new_AGEMA_signal_938, stateFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({data_out_s1[33], data_out_s0[33]}), .a ({data_in_s1[24], data_in_s0[24]}), .c ({new_AGEMA_signal_941, stateFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({data_out_s1[37], data_out_s0[37]}), .a ({data_in_s1[25], data_in_s0[25]}), .c ({new_AGEMA_signal_944, stateFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({data_out_s1[41], data_out_s0[41]}), .a ({data_in_s1[26], data_in_s0[26]}), .c ({new_AGEMA_signal_947, stateFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({data_out_s1[45], data_out_s0[45]}), .a ({data_in_s1[27], data_in_s0[27]}), .c ({new_AGEMA_signal_950, stateFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({data_out_s1[49], data_out_s0[49]}), .a ({data_in_s1[28], data_in_s0[28]}), .c ({new_AGEMA_signal_953, stateFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({data_out_s1[53], data_out_s0[53]}), .a ({data_in_s1[29], data_in_s0[29]}), .c ({new_AGEMA_signal_956, stateFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({data_out_s1[57], data_out_s0[57]}), .a ({data_in_s1[30], data_in_s0[30]}), .c ({new_AGEMA_signal_959, stateFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({data_out_s1[61], data_out_s0[61]}), .a ({data_in_s1[31], data_in_s0[31]}), .c ({new_AGEMA_signal_961, stateFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({data_out_s1[2], data_out_s0[2]}), .a ({data_in_s1[32], data_in_s0[32]}), .c ({new_AGEMA_signal_964, stateFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({data_out_s1[6], data_out_s0[6]}), .a ({data_in_s1[33], data_in_s0[33]}), .c ({new_AGEMA_signal_967, stateFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({data_out_s1[10], data_out_s0[10]}), .a ({data_in_s1[34], data_in_s0[34]}), .c ({new_AGEMA_signal_970, stateFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({data_out_s1[14], data_out_s0[14]}), .a ({data_in_s1[35], data_in_s0[35]}), .c ({new_AGEMA_signal_973, stateFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({data_out_s1[18], data_out_s0[18]}), .a ({data_in_s1[36], data_in_s0[36]}), .c ({new_AGEMA_signal_976, stateFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({data_out_s1[22], data_out_s0[22]}), .a ({data_in_s1[37], data_in_s0[37]}), .c ({new_AGEMA_signal_979, stateFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({data_out_s1[26], data_out_s0[26]}), .a ({data_in_s1[38], data_in_s0[38]}), .c ({new_AGEMA_signal_982, stateFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({data_out_s1[30], data_out_s0[30]}), .a ({data_in_s1[39], data_in_s0[39]}), .c ({new_AGEMA_signal_985, stateFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({data_out_s1[34], data_out_s0[34]}), .a ({data_in_s1[40], data_in_s0[40]}), .c ({new_AGEMA_signal_988, stateFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({data_out_s1[38], data_out_s0[38]}), .a ({data_in_s1[41], data_in_s0[41]}), .c ({new_AGEMA_signal_991, stateFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({data_out_s1[42], data_out_s0[42]}), .a ({data_in_s1[42], data_in_s0[42]}), .c ({new_AGEMA_signal_994, stateFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({data_out_s1[46], data_out_s0[46]}), .a ({data_in_s1[43], data_in_s0[43]}), .c ({new_AGEMA_signal_997, stateFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({data_out_s1[50], data_out_s0[50]}), .a ({data_in_s1[44], data_in_s0[44]}), .c ({new_AGEMA_signal_1000, stateFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({data_out_s1[54], data_out_s0[54]}), .a ({data_in_s1[45], data_in_s0[45]}), .c ({new_AGEMA_signal_1003, stateFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({data_out_s1[58], data_out_s0[58]}), .a ({data_in_s1[46], data_in_s0[46]}), .c ({new_AGEMA_signal_1006, stateFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({data_out_s1[62], data_out_s0[62]}), .a ({data_in_s1[47], data_in_s0[47]}), .c ({new_AGEMA_signal_1008, stateFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({data_out_s1[3], data_out_s0[3]}), .a ({data_in_s1[48], data_in_s0[48]}), .c ({new_AGEMA_signal_1011, stateFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({data_out_s1[7], data_out_s0[7]}), .a ({data_in_s1[49], data_in_s0[49]}), .c ({new_AGEMA_signal_1014, stateFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({data_out_s1[11], data_out_s0[11]}), .a ({data_in_s1[50], data_in_s0[50]}), .c ({new_AGEMA_signal_1017, stateFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({data_out_s1[15], data_out_s0[15]}), .a ({data_in_s1[51], data_in_s0[51]}), .c ({new_AGEMA_signal_1020, stateFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({data_out_s1[19], data_out_s0[19]}), .a ({data_in_s1[52], data_in_s0[52]}), .c ({new_AGEMA_signal_1023, stateFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({data_out_s1[23], data_out_s0[23]}), .a ({data_in_s1[53], data_in_s0[53]}), .c ({new_AGEMA_signal_1026, stateFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({data_out_s1[27], data_out_s0[27]}), .a ({data_in_s1[54], data_in_s0[54]}), .c ({new_AGEMA_signal_1029, stateFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({data_out_s1[31], data_out_s0[31]}), .a ({data_in_s1[55], data_in_s0[55]}), .c ({new_AGEMA_signal_1032, stateFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({data_out_s1[35], data_out_s0[35]}), .a ({data_in_s1[56], data_in_s0[56]}), .c ({new_AGEMA_signal_1035, stateFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({data_out_s1[39], data_out_s0[39]}), .a ({data_in_s1[57], data_in_s0[57]}), .c ({new_AGEMA_signal_1038, stateFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({data_out_s1[43], data_out_s0[43]}), .a ({data_in_s1[58], data_in_s0[58]}), .c ({new_AGEMA_signal_1041, stateFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({data_out_s1[47], data_out_s0[47]}), .a ({data_in_s1[59], data_in_s0[59]}), .c ({new_AGEMA_signal_1044, stateFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({data_out_s1[51], data_out_s0[51]}), .a ({data_in_s1[60], data_in_s0[60]}), .c ({new_AGEMA_signal_1047, stateFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({data_out_s1[55], data_out_s0[55]}), .a ({data_in_s1[61], data_in_s0[61]}), .c ({new_AGEMA_signal_1050, stateFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({data_out_s1[59], data_out_s0[59]}), .a ({data_in_s1[62], data_in_s0[62]}), .c ({new_AGEMA_signal_1053, stateFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({data_out_s1[63], data_out_s0[63]}), .a ({data_in_s1[63], data_in_s0[63]}), .c ({new_AGEMA_signal_1055, stateFF_inputPar[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) keyFF_U5 ( .a ({1'b0, counter[4]}), .b ({new_AGEMA_signal_1056, keyFF_outputPar[22]}), .c ({new_AGEMA_signal_1057, keyFF_counterAdd[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) keyFF_U4 ( .a ({1'b0, counter[3]}), .b ({new_AGEMA_signal_1058, keyFF_outputPar[21]}), .c ({new_AGEMA_signal_1059, keyFF_counterAdd[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) keyFF_U3 ( .a ({1'b0, counter[2]}), .b ({new_AGEMA_signal_1060, keyFF_outputPar[20]}), .c ({new_AGEMA_signal_1061, keyFF_counterAdd[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) keyFF_U2 ( .a ({1'b0, counter[1]}), .b ({new_AGEMA_signal_1274, keyFF_outputPar[19]}), .c ({new_AGEMA_signal_1275, keyFF_counterAdd[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) keyFF_U1 ( .a ({1'b0, counter[0]}), .b ({new_AGEMA_signal_1062, keyFF_outputPar[18]}), .c ({new_AGEMA_signal_1063, keyFF_counterAdd[0]}) ) ;
    INV_X1 keyFF_keystate_U3 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n6) ) ;
    INV_X1 keyFF_keystate_U2 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n7) ) ;
    INV_X1 keyFF_keystate_U1 ( .A (ctrlData_0_), .ZN (keyFF_keystate_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_856, roundkey[0]}), .a ({new_AGEMA_signal_1066, keyFF_inputPar[0]}), .c ({new_AGEMA_signal_1374, keyFF_keystate_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_859, roundkey[1]}), .a ({new_AGEMA_signal_1069, keyFF_inputPar[1]}), .c ({new_AGEMA_signal_1375, keyFF_keystate_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_862, roundkey[2]}), .a ({new_AGEMA_signal_1072, keyFF_inputPar[2]}), .c ({new_AGEMA_signal_1376, keyFF_keystate_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_865, roundkey[3]}), .a ({new_AGEMA_signal_1075, keyFF_inputPar[3]}), .c ({new_AGEMA_signal_1377, keyFF_keystate_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1287, keyRegKS[1]}), .a ({new_AGEMA_signal_1078, keyFF_inputPar[4]}), .c ({new_AGEMA_signal_1378, keyFF_keystate_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1289, keyRegKS[2]}), .a ({new_AGEMA_signal_1081, keyFF_inputPar[5]}), .c ({new_AGEMA_signal_1379, keyFF_keystate_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1291, keyRegKS[3]}), .a ({new_AGEMA_signal_1084, keyFF_inputPar[6]}), .c ({new_AGEMA_signal_1380, keyFF_keystate_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1064, keyFF_outputPar[3]}), .a ({new_AGEMA_signal_1087, keyFF_inputPar[7]}), .c ({new_AGEMA_signal_1381, keyFF_keystate_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1067, keyFF_outputPar[4]}), .a ({new_AGEMA_signal_1090, keyFF_inputPar[8]}), .c ({new_AGEMA_signal_1382, keyFF_keystate_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1070, keyFF_outputPar[5]}), .a ({new_AGEMA_signal_1093, keyFF_inputPar[9]}), .c ({new_AGEMA_signal_1383, keyFF_keystate_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1073, keyFF_outputPar[6]}), .a ({new_AGEMA_signal_1096, keyFF_inputPar[10]}), .c ({new_AGEMA_signal_1384, keyFF_keystate_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1076, keyFF_outputPar[7]}), .a ({new_AGEMA_signal_1099, keyFF_inputPar[11]}), .c ({new_AGEMA_signal_1385, keyFF_keystate_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1079, keyFF_outputPar[8]}), .a ({new_AGEMA_signal_1102, keyFF_inputPar[12]}), .c ({new_AGEMA_signal_1386, keyFF_keystate_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1082, keyFF_outputPar[9]}), .a ({new_AGEMA_signal_1105, keyFF_inputPar[13]}), .c ({new_AGEMA_signal_1387, keyFF_keystate_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1085, keyFF_outputPar[10]}), .a ({new_AGEMA_signal_1108, keyFF_inputPar[14]}), .c ({new_AGEMA_signal_1388, keyFF_keystate_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1088, keyFF_outputPar[11]}), .a ({new_AGEMA_signal_1277, keyFF_inputPar[15]}), .c ({new_AGEMA_signal_1389, keyFF_keystate_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1091, keyFF_outputPar[12]}), .a ({new_AGEMA_signal_1285, keyFF_inputPar[16]}), .c ({new_AGEMA_signal_1303, keyFF_keystate_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1094, keyFF_outputPar[13]}), .a ({new_AGEMA_signal_1279, keyFF_inputPar[17]}), .c ({new_AGEMA_signal_1304, keyFF_keystate_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1097, keyFF_outputPar[14]}), .a ({new_AGEMA_signal_1281, keyFF_inputPar[18]}), .c ({new_AGEMA_signal_1305, keyFF_keystate_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1100, keyFF_outputPar[15]}), .a ({new_AGEMA_signal_1283, keyFF_inputPar[19]}), .c ({new_AGEMA_signal_1306, keyFF_keystate_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1103, keyFF_outputPar[16]}), .a ({new_AGEMA_signal_1111, keyFF_inputPar[20]}), .c ({new_AGEMA_signal_1307, keyFF_keystate_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1106, keyFF_outputPar[17]}), .a ({new_AGEMA_signal_1114, keyFF_inputPar[21]}), .c ({new_AGEMA_signal_1308, keyFF_keystate_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1062, keyFF_outputPar[18]}), .a ({new_AGEMA_signal_1117, keyFF_inputPar[22]}), .c ({new_AGEMA_signal_1309, keyFF_keystate_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1274, keyFF_outputPar[19]}), .a ({new_AGEMA_signal_1120, keyFF_inputPar[23]}), .c ({new_AGEMA_signal_1310, keyFF_keystate_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1060, keyFF_outputPar[20]}), .a ({new_AGEMA_signal_1123, keyFF_inputPar[24]}), .c ({new_AGEMA_signal_1390, keyFF_keystate_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1058, keyFF_outputPar[21]}), .a ({new_AGEMA_signal_1126, keyFF_inputPar[25]}), .c ({new_AGEMA_signal_1391, keyFF_keystate_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1056, keyFF_outputPar[22]}), .a ({new_AGEMA_signal_1129, keyFF_inputPar[26]}), .c ({new_AGEMA_signal_1392, keyFF_keystate_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1109, keyFF_outputPar[23]}), .a ({new_AGEMA_signal_1132, keyFF_inputPar[27]}), .c ({new_AGEMA_signal_1393, keyFF_keystate_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1112, keyFF_outputPar[24]}), .a ({new_AGEMA_signal_1135, keyFF_inputPar[28]}), .c ({new_AGEMA_signal_1394, keyFF_keystate_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1115, keyFF_outputPar[25]}), .a ({new_AGEMA_signal_1138, keyFF_inputPar[29]}), .c ({new_AGEMA_signal_1395, keyFF_keystate_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1118, keyFF_outputPar[26]}), .a ({new_AGEMA_signal_1141, keyFF_inputPar[30]}), .c ({new_AGEMA_signal_1396, keyFF_keystate_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1121, keyFF_outputPar[27]}), .a ({new_AGEMA_signal_1144, keyFF_inputPar[31]}), .c ({new_AGEMA_signal_1397, keyFF_keystate_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1124, keyFF_outputPar[28]}), .a ({new_AGEMA_signal_1147, keyFF_inputPar[32]}), .c ({new_AGEMA_signal_1398, keyFF_keystate_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1127, keyFF_outputPar[29]}), .a ({new_AGEMA_signal_1150, keyFF_inputPar[33]}), .c ({new_AGEMA_signal_1399, keyFF_keystate_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1130, keyFF_outputPar[30]}), .a ({new_AGEMA_signal_1153, keyFF_inputPar[34]}), .c ({new_AGEMA_signal_1400, keyFF_keystate_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1133, keyFF_outputPar[31]}), .a ({new_AGEMA_signal_1156, keyFF_inputPar[35]}), .c ({new_AGEMA_signal_1401, keyFF_keystate_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1136, keyFF_outputPar[32]}), .a ({new_AGEMA_signal_1159, keyFF_inputPar[36]}), .c ({new_AGEMA_signal_1402, keyFF_keystate_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1139, keyFF_outputPar[33]}), .a ({new_AGEMA_signal_1162, keyFF_inputPar[37]}), .c ({new_AGEMA_signal_1403, keyFF_keystate_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1142, keyFF_outputPar[34]}), .a ({new_AGEMA_signal_1165, keyFF_inputPar[38]}), .c ({new_AGEMA_signal_1404, keyFF_keystate_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1145, keyFF_outputPar[35]}), .a ({new_AGEMA_signal_1168, keyFF_inputPar[39]}), .c ({new_AGEMA_signal_1405, keyFF_keystate_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1148, keyFF_outputPar[36]}), .a ({new_AGEMA_signal_1171, keyFF_inputPar[40]}), .c ({new_AGEMA_signal_1406, keyFF_keystate_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1151, keyFF_outputPar[37]}), .a ({new_AGEMA_signal_1174, keyFF_inputPar[41]}), .c ({new_AGEMA_signal_1407, keyFF_keystate_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1154, keyFF_outputPar[38]}), .a ({new_AGEMA_signal_1177, keyFF_inputPar[42]}), .c ({new_AGEMA_signal_1408, keyFF_keystate_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1157, keyFF_outputPar[39]}), .a ({new_AGEMA_signal_1180, keyFF_inputPar[43]}), .c ({new_AGEMA_signal_1409, keyFF_keystate_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1160, keyFF_outputPar[40]}), .a ({new_AGEMA_signal_1183, keyFF_inputPar[44]}), .c ({new_AGEMA_signal_1410, keyFF_keystate_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1163, keyFF_outputPar[41]}), .a ({new_AGEMA_signal_1186, keyFF_inputPar[45]}), .c ({new_AGEMA_signal_1411, keyFF_keystate_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1166, keyFF_outputPar[42]}), .a ({new_AGEMA_signal_1189, keyFF_inputPar[46]}), .c ({new_AGEMA_signal_1412, keyFF_keystate_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1169, keyFF_outputPar[43]}), .a ({new_AGEMA_signal_1192, keyFF_inputPar[47]}), .c ({new_AGEMA_signal_1413, keyFF_keystate_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1172, keyFF_outputPar[44]}), .a ({new_AGEMA_signal_1195, keyFF_inputPar[48]}), .c ({new_AGEMA_signal_1414, keyFF_keystate_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1175, keyFF_outputPar[45]}), .a ({new_AGEMA_signal_1198, keyFF_inputPar[49]}), .c ({new_AGEMA_signal_1415, keyFF_keystate_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1178, keyFF_outputPar[46]}), .a ({new_AGEMA_signal_1201, keyFF_inputPar[50]}), .c ({new_AGEMA_signal_1416, keyFF_keystate_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1181, keyFF_outputPar[47]}), .a ({new_AGEMA_signal_1204, keyFF_inputPar[51]}), .c ({new_AGEMA_signal_1417, keyFF_keystate_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1184, keyFF_outputPar[48]}), .a ({new_AGEMA_signal_1207, keyFF_inputPar[52]}), .c ({new_AGEMA_signal_1418, keyFF_keystate_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1187, keyFF_outputPar[49]}), .a ({new_AGEMA_signal_1210, keyFF_inputPar[53]}), .c ({new_AGEMA_signal_1419, keyFF_keystate_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1190, keyFF_outputPar[50]}), .a ({new_AGEMA_signal_1213, keyFF_inputPar[54]}), .c ({new_AGEMA_signal_1420, keyFF_keystate_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1193, keyFF_outputPar[51]}), .a ({new_AGEMA_signal_1216, keyFF_inputPar[55]}), .c ({new_AGEMA_signal_1421, keyFF_keystate_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1196, keyFF_outputPar[52]}), .a ({new_AGEMA_signal_1219, keyFF_inputPar[56]}), .c ({new_AGEMA_signal_1422, keyFF_keystate_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1199, keyFF_outputPar[53]}), .a ({new_AGEMA_signal_1222, keyFF_inputPar[57]}), .c ({new_AGEMA_signal_1423, keyFF_keystate_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1202, keyFF_outputPar[54]}), .a ({new_AGEMA_signal_1225, keyFF_inputPar[58]}), .c ({new_AGEMA_signal_1424, keyFF_keystate_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1205, keyFF_outputPar[55]}), .a ({new_AGEMA_signal_1228, keyFF_inputPar[59]}), .c ({new_AGEMA_signal_1425, keyFF_keystate_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1208, keyFF_outputPar[56]}), .a ({new_AGEMA_signal_1231, keyFF_inputPar[60]}), .c ({new_AGEMA_signal_1426, keyFF_keystate_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1211, keyFF_outputPar[57]}), .a ({new_AGEMA_signal_1234, keyFF_inputPar[61]}), .c ({new_AGEMA_signal_1427, keyFF_keystate_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1214, keyFF_outputPar[58]}), .a ({new_AGEMA_signal_1237, keyFF_inputPar[62]}), .c ({new_AGEMA_signal_1428, keyFF_keystate_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1217, keyFF_outputPar[59]}), .a ({new_AGEMA_signal_1240, keyFF_inputPar[63]}), .c ({new_AGEMA_signal_1429, keyFF_keystate_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1220, keyFF_outputPar[60]}), .a ({new_AGEMA_signal_1243, keyFF_inputPar[64]}), .c ({new_AGEMA_signal_1430, keyFF_keystate_gff_17_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1223, keyFF_outputPar[61]}), .a ({new_AGEMA_signal_1246, keyFF_inputPar[65]}), .c ({new_AGEMA_signal_1431, keyFF_keystate_gff_17_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1226, keyFF_outputPar[62]}), .a ({new_AGEMA_signal_1249, keyFF_inputPar[66]}), .c ({new_AGEMA_signal_1432, keyFF_keystate_gff_17_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1229, keyFF_outputPar[63]}), .a ({new_AGEMA_signal_1252, keyFF_inputPar[67]}), .c ({new_AGEMA_signal_1433, keyFF_keystate_gff_17_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1232, keyFF_outputPar[64]}), .a ({new_AGEMA_signal_1255, keyFF_inputPar[68]}), .c ({new_AGEMA_signal_1434, keyFF_keystate_gff_18_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1235, keyFF_outputPar[65]}), .a ({new_AGEMA_signal_1258, keyFF_inputPar[69]}), .c ({new_AGEMA_signal_1435, keyFF_keystate_gff_18_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1238, keyFF_outputPar[66]}), .a ({new_AGEMA_signal_1261, keyFF_inputPar[70]}), .c ({new_AGEMA_signal_1436, keyFF_keystate_gff_18_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1241, keyFF_outputPar[67]}), .a ({new_AGEMA_signal_1264, keyFF_inputPar[71]}), .c ({new_AGEMA_signal_1437, keyFF_keystate_gff_18_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1244, keyFF_outputPar[68]}), .a ({new_AGEMA_signal_1267, keyFF_inputPar[72]}), .c ({new_AGEMA_signal_1438, keyFF_keystate_gff_19_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1247, keyFF_outputPar[69]}), .a ({new_AGEMA_signal_1269, keyFF_inputPar[73]}), .c ({new_AGEMA_signal_1439, keyFF_keystate_gff_19_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1250, keyFF_outputPar[70]}), .a ({new_AGEMA_signal_1271, keyFF_inputPar[74]}), .c ({new_AGEMA_signal_1440, keyFF_keystate_gff_19_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1253, keyFF_outputPar[71]}), .a ({new_AGEMA_signal_1273, keyFF_inputPar[75]}), .c ({new_AGEMA_signal_1441, keyFF_keystate_gff_19_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({new_AGEMA_signal_1064, keyFF_outputPar[3]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1066, keyFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({new_AGEMA_signal_1067, keyFF_outputPar[4]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1069, keyFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({new_AGEMA_signal_1070, keyFF_outputPar[5]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1072, keyFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({new_AGEMA_signal_1073, keyFF_outputPar[6]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1075, keyFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({new_AGEMA_signal_1076, keyFF_outputPar[7]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1078, keyFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({new_AGEMA_signal_1079, keyFF_outputPar[8]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1081, keyFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({new_AGEMA_signal_1082, keyFF_outputPar[9]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1084, keyFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({new_AGEMA_signal_1085, keyFF_outputPar[10]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1087, keyFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({new_AGEMA_signal_1088, keyFF_outputPar[11]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1090, keyFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({new_AGEMA_signal_1091, keyFF_outputPar[12]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1093, keyFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({new_AGEMA_signal_1094, keyFF_outputPar[13]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1096, keyFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({new_AGEMA_signal_1097, keyFF_outputPar[14]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1099, keyFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({new_AGEMA_signal_1100, keyFF_outputPar[15]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1102, keyFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({new_AGEMA_signal_1103, keyFF_outputPar[16]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1105, keyFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({new_AGEMA_signal_1106, keyFF_outputPar[17]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1108, keyFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({new_AGEMA_signal_1063, keyFF_counterAdd[0]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1277, keyFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({new_AGEMA_signal_1275, keyFF_counterAdd[1]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1285, keyFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({new_AGEMA_signal_1061, keyFF_counterAdd[2]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1279, keyFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({new_AGEMA_signal_1059, keyFF_counterAdd[3]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1281, keyFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({new_AGEMA_signal_1057, keyFF_counterAdd[4]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1283, keyFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({new_AGEMA_signal_1109, keyFF_outputPar[23]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1111, keyFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({new_AGEMA_signal_1112, keyFF_outputPar[24]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1114, keyFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({new_AGEMA_signal_1115, keyFF_outputPar[25]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1117, keyFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({new_AGEMA_signal_1118, keyFF_outputPar[26]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1120, keyFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({new_AGEMA_signal_1121, keyFF_outputPar[27]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1123, keyFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({new_AGEMA_signal_1124, keyFF_outputPar[28]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1126, keyFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({new_AGEMA_signal_1127, keyFF_outputPar[29]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1129, keyFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({new_AGEMA_signal_1130, keyFF_outputPar[30]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1132, keyFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({new_AGEMA_signal_1133, keyFF_outputPar[31]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1135, keyFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({new_AGEMA_signal_1136, keyFF_outputPar[32]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1138, keyFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({new_AGEMA_signal_1139, keyFF_outputPar[33]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1141, keyFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({new_AGEMA_signal_1142, keyFF_outputPar[34]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1144, keyFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({new_AGEMA_signal_1145, keyFF_outputPar[35]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_1147, keyFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({new_AGEMA_signal_1148, keyFF_outputPar[36]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1150, keyFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({new_AGEMA_signal_1151, keyFF_outputPar[37]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_1153, keyFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({new_AGEMA_signal_1154, keyFF_outputPar[38]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_1156, keyFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({new_AGEMA_signal_1157, keyFF_outputPar[39]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1159, keyFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({new_AGEMA_signal_1160, keyFF_outputPar[40]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1162, keyFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({new_AGEMA_signal_1163, keyFF_outputPar[41]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1165, keyFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({new_AGEMA_signal_1166, keyFF_outputPar[42]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1168, keyFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({new_AGEMA_signal_1169, keyFF_outputPar[43]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1171, keyFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({new_AGEMA_signal_1172, keyFF_outputPar[44]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1174, keyFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({new_AGEMA_signal_1175, keyFF_outputPar[45]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1177, keyFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({new_AGEMA_signal_1178, keyFF_outputPar[46]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1180, keyFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({new_AGEMA_signal_1181, keyFF_outputPar[47]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1183, keyFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({new_AGEMA_signal_1184, keyFF_outputPar[48]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1186, keyFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({new_AGEMA_signal_1187, keyFF_outputPar[49]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1189, keyFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({new_AGEMA_signal_1190, keyFF_outputPar[50]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1192, keyFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({new_AGEMA_signal_1193, keyFF_outputPar[51]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1195, keyFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({new_AGEMA_signal_1196, keyFF_outputPar[52]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1198, keyFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({new_AGEMA_signal_1199, keyFF_outputPar[53]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1201, keyFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({new_AGEMA_signal_1202, keyFF_outputPar[54]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1204, keyFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({new_AGEMA_signal_1205, keyFF_outputPar[55]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1207, keyFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({new_AGEMA_signal_1208, keyFF_outputPar[56]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1210, keyFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({new_AGEMA_signal_1211, keyFF_outputPar[57]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1213, keyFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({new_AGEMA_signal_1214, keyFF_outputPar[58]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1216, keyFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({new_AGEMA_signal_1217, keyFF_outputPar[59]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1219, keyFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({new_AGEMA_signal_1220, keyFF_outputPar[60]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1222, keyFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({new_AGEMA_signal_1223, keyFF_outputPar[61]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1225, keyFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({new_AGEMA_signal_1226, keyFF_outputPar[62]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1228, keyFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({new_AGEMA_signal_1229, keyFF_outputPar[63]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1231, keyFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({new_AGEMA_signal_1232, keyFF_outputPar[64]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1234, keyFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({new_AGEMA_signal_1235, keyFF_outputPar[65]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1237, keyFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({new_AGEMA_signal_1238, keyFF_outputPar[66]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1240, keyFF_inputPar[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_64_U1 ( .s (reset), .b ({new_AGEMA_signal_1241, keyFF_outputPar[67]}), .a ({key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1243, keyFF_inputPar[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_65_U1 ( .s (reset), .b ({new_AGEMA_signal_1244, keyFF_outputPar[68]}), .a ({key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1246, keyFF_inputPar[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_66_U1 ( .s (reset), .b ({new_AGEMA_signal_1247, keyFF_outputPar[69]}), .a ({key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1249, keyFF_inputPar[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_67_U1 ( .s (reset), .b ({new_AGEMA_signal_1250, keyFF_outputPar[70]}), .a ({key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1252, keyFF_inputPar[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_68_U1 ( .s (reset), .b ({new_AGEMA_signal_1253, keyFF_outputPar[71]}), .a ({key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1255, keyFF_inputPar[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_69_U1 ( .s (reset), .b ({new_AGEMA_signal_1256, keyFF_outputPar[72]}), .a ({key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1258, keyFF_inputPar[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_70_U1 ( .s (reset), .b ({new_AGEMA_signal_1259, keyFF_outputPar[73]}), .a ({key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1261, keyFF_inputPar[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_71_U1 ( .s (reset), .b ({new_AGEMA_signal_1262, keyFF_outputPar[74]}), .a ({key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_1264, keyFF_inputPar[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_72_U1 ( .s (reset), .b ({new_AGEMA_signal_1265, keyFF_outputPar[75]}), .a ({key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_1267, keyFF_inputPar[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_73_U1 ( .s (reset), .b ({new_AGEMA_signal_856, roundkey[0]}), .a ({key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_1269, keyFF_inputPar[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_74_U1 ( .s (reset), .b ({new_AGEMA_signal_859, roundkey[1]}), .a ({key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1271, keyFF_inputPar[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_75_U1 ( .s (reset), .b ({new_AGEMA_signal_862, roundkey[2]}), .a ({key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1273, keyFF_inputPar[75]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) sboxInst_U3 ( .a ({new_AGEMA_signal_1295, sboxInst_L0}), .b ({new_AGEMA_signal_1311, sboxInst_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) sboxInst_U2 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1293, sboxInst_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) sboxInst_U1 ( .a ({new_AGEMA_signal_1288, sboxIn[1]}), .b ({new_AGEMA_signal_1294, sboxInst_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR1_U1 ( .a ({new_AGEMA_signal_1290, sboxIn[2]}), .b ({new_AGEMA_signal_1288, sboxIn[1]}), .c ({new_AGEMA_signal_1295, sboxInst_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR2_U1 ( .a ({new_AGEMA_signal_1288, sboxIn[1]}), .b ({new_AGEMA_signal_1286, sboxIn[0]}), .c ({new_AGEMA_signal_1296, sboxInst_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR3_U1 ( .a ({new_AGEMA_signal_1296, sboxInst_L1}), .b ({new_AGEMA_signal_1292, sboxIn[3]}), .c ({new_AGEMA_signal_1312, sboxInst_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR4_U1 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1286, sboxIn[0]}), .c ({new_AGEMA_signal_1297, sboxInst_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR5_U1 ( .a ({new_AGEMA_signal_1297, sboxInst_L3}), .b ({new_AGEMA_signal_1295, sboxInst_L0}), .c ({new_AGEMA_signal_1313, sboxInst_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR6_U1 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1288, sboxIn[1]}), .c ({new_AGEMA_signal_1298, sboxInst_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR9_U1 ( .a ({new_AGEMA_signal_1296, sboxInst_L1}), .b ({new_AGEMA_signal_1290, sboxIn[2]}), .c ({new_AGEMA_signal_1314, sboxInst_Q7}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_sboxin_mux_inst_0_U1 ( .s (selSbox), .b ({new_AGEMA_signal_858, stateXORroundkey[0]}), .a ({new_AGEMA_signal_865, roundkey[3]}), .c ({new_AGEMA_signal_1286, sboxIn[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_sboxin_mux_inst_1_U1 ( .s (selSbox), .b ({new_AGEMA_signal_861, stateXORroundkey[1]}), .a ({new_AGEMA_signal_1287, keyRegKS[1]}), .c ({new_AGEMA_signal_1288, sboxIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_sboxin_mux_inst_2_U1 ( .s (selSbox), .b ({new_AGEMA_signal_864, stateXORroundkey[2]}), .a ({new_AGEMA_signal_1289, keyRegKS[2]}), .c ({new_AGEMA_signal_1290, sboxIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_sboxin_mux_inst_3_U1 ( .s (selSbox), .b ({new_AGEMA_signal_867, stateXORroundkey[3]}), .a ({new_AGEMA_signal_1291, keyRegKS[3]}), .c ({new_AGEMA_signal_1292, sboxIn[3]}) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1446, serialIn[0]}), .a ({new_AGEMA_signal_870, stateFF_inputPar[0]}), .c ({new_AGEMA_signal_1447, stateFF_state_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1256, keyFF_outputPar[72]}), .a ({new_AGEMA_signal_1443, keyFF_inputPar[76]}), .c ({new_AGEMA_signal_1448, keyFF_keystate_gff_20_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_76_U1 ( .s (reset), .b ({new_AGEMA_signal_1317, sboxOut[0]}), .a ({key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_1443, keyFF_inputPar[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR16_U1 ( .a ({new_AGEMA_signal_1316, sboxInst_T0}), .b ({new_AGEMA_signal_1312, sboxInst_L2}), .c ({new_AGEMA_signal_1444, sboxInst_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR7_U1 ( .a ({new_AGEMA_signal_1316, sboxInst_T0}), .b ({new_AGEMA_signal_1315, sboxInst_T2}), .c ({new_AGEMA_signal_1445, sboxInst_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR8_U1 ( .a ({new_AGEMA_signal_1298, sboxInst_L4}), .b ({new_AGEMA_signal_1445, sboxInst_L5}), .c ({new_AGEMA_signal_1449, sboxInst_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_AND1_U1 ( .a ({new_AGEMA_signal_1311, sboxInst_n1}), .b ({new_AGEMA_signal_1293, sboxInst_n2}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1316, sboxInst_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_AND3_U1 ( .a ({new_AGEMA_signal_1294, sboxInst_n3}), .b ({new_AGEMA_signal_1290, sboxIn[2]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1315, sboxInst_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR15_U1 ( .a ({new_AGEMA_signal_1297, sboxInst_L3}), .b ({new_AGEMA_signal_1315, sboxInst_T2}), .c ({new_AGEMA_signal_1317, sboxOut[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_serialIn_mux_inst_0_U1 ( .s (intDone), .b ({new_AGEMA_signal_1317, sboxOut[0]}), .a ({new_AGEMA_signal_858, stateXORroundkey[0]}), .c ({new_AGEMA_signal_1446, serialIn[0]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1461, serialIn[1]}), .a ({new_AGEMA_signal_873, stateFF_inputPar[1]}), .c ({new_AGEMA_signal_1463, stateFF_state_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1462, serialIn[2]}), .a ({new_AGEMA_signal_876, stateFF_inputPar[2]}), .c ({new_AGEMA_signal_1464, stateFF_state_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1469, serialIn[3]}), .a ({new_AGEMA_signal_879, stateFF_inputPar[3]}), .c ({new_AGEMA_signal_1470, stateFF_state_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1259, keyFF_outputPar[73]}), .a ({new_AGEMA_signal_1457, keyFF_inputPar[77]}), .c ({new_AGEMA_signal_1465, keyFF_keystate_gff_20_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1262, keyFF_outputPar[74]}), .a ({new_AGEMA_signal_1459, keyFF_inputPar[78]}), .c ({new_AGEMA_signal_1466, keyFF_keystate_gff_20_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1265, keyFF_outputPar[75]}), .a ({new_AGEMA_signal_1468, keyFF_inputPar[79]}), .c ({new_AGEMA_signal_1471, keyFF_keystate_gff_20_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_77_U1 ( .s (reset), .b ({new_AGEMA_signal_1455, sboxOut[1]}), .a ({key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1457, keyFF_inputPar[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_78_U1 ( .s (reset), .b ({new_AGEMA_signal_1454, sboxOut[2]}), .a ({key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1459, keyFF_inputPar[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) keyFF_MUX_inputPar_mux_inst_79_U1 ( .s (reset), .b ({new_AGEMA_signal_1460, sboxOut[3]}), .a ({key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1468, keyFF_inputPar[79]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_AND2_U1 ( .a ({new_AGEMA_signal_1444, sboxInst_Q2}), .b ({new_AGEMA_signal_1313, sboxInst_Q3}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1450, sboxInst_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_AND4_U1 ( .a ({new_AGEMA_signal_1449, sboxInst_Q6}), .b ({new_AGEMA_signal_1314, sboxInst_Q7}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1451, sboxInst_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR10_U1 ( .a ({new_AGEMA_signal_1445, sboxInst_L5}), .b ({new_AGEMA_signal_1451, sboxInst_T3}), .c ({new_AGEMA_signal_1453, sboxInst_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR11_U1 ( .a ({new_AGEMA_signal_1286, sboxIn[0]}), .b ({new_AGEMA_signal_1453, sboxInst_L7}), .c ({new_AGEMA_signal_1460, sboxOut[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR12_U1 ( .a ({new_AGEMA_signal_1445, sboxInst_L5}), .b ({new_AGEMA_signal_1450, sboxInst_T1}), .c ({new_AGEMA_signal_1452, sboxInst_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR13_U1 ( .a ({new_AGEMA_signal_1296, sboxInst_L1}), .b ({new_AGEMA_signal_1452, sboxInst_L8}), .c ({new_AGEMA_signal_1454, sboxOut[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sboxInst_XOR14_U1 ( .a ({new_AGEMA_signal_1298, sboxInst_L4}), .b ({new_AGEMA_signal_1451, sboxInst_T3}), .c ({new_AGEMA_signal_1455, sboxOut[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_serialIn_mux_inst_1_U1 ( .s (intDone), .b ({new_AGEMA_signal_1455, sboxOut[1]}), .a ({new_AGEMA_signal_861, stateXORroundkey[1]}), .c ({new_AGEMA_signal_1461, serialIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_serialIn_mux_inst_2_U1 ( .s (intDone), .b ({new_AGEMA_signal_1454, sboxOut[2]}), .a ({new_AGEMA_signal_864, stateXORroundkey[2]}), .c ({new_AGEMA_signal_1462, serialIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_serialIn_mux_inst_3_U1 ( .s (intDone), .b ({new_AGEMA_signal_1460, sboxOut[3]}), .a ({new_AGEMA_signal_867, stateXORroundkey[3]}), .c ({new_AGEMA_signal_1469, serialIn[3]}) ) ;

    /* register cells */
    DFF_X1 fsm_cnt_rnd_count_reg_reg_4__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n14), .Q (counter[4]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_2__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n16), .Q (counter[2]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n18), .Q (counter[0]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_3__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n1), .Q (counter[3]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_cnt_rnd_n41), .Q (fsm_cnt_rnd_n24), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_2__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n1), .Q (fsm_countSerial[2]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n3), .Q (fsm_countSerial[0]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_3__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n26), .Q (fsm_countSerial[3]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_cnt_ser_n28), .Q (fsm_countSerial[1]), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_0__FF_FF ( .CK (clk_gated), .D (fsm_n21), .Q (fsm_ps_state_0_), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_1__FF_FF ( .CK (clk_gated), .D (fsm_n20), .Q (fsm_ps_state_1_), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1447, stateFF_state_gff_1_s_next_state[0]}), .Q ({data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1464, stateFF_state_gff_1_s_next_state[2]}), .Q ({data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1463, stateFF_state_gff_1_s_next_state[1]}), .Q ({data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1470, stateFF_state_gff_1_s_next_state[3]}), .Q ({data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1302, stateFF_state_gff_2_s_next_state[3]}), .Q ({data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1301, stateFF_state_gff_2_s_next_state[2]}), .Q ({data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1300, stateFF_state_gff_2_s_next_state[1]}), .Q ({data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1299, stateFF_state_gff_2_s_next_state[0]}), .Q ({data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1321, stateFF_state_gff_3_s_next_state[3]}), .Q ({data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1320, stateFF_state_gff_3_s_next_state[2]}), .Q ({data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1319, stateFF_state_gff_3_s_next_state[1]}), .Q ({data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1318, stateFF_state_gff_3_s_next_state[0]}), .Q ({data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1325, stateFF_state_gff_4_s_next_state[3]}), .Q ({data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1324, stateFF_state_gff_4_s_next_state[2]}), .Q ({data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1323, stateFF_state_gff_4_s_next_state[1]}), .Q ({data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1322, stateFF_state_gff_4_s_next_state[0]}), .Q ({data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1329, stateFF_state_gff_5_s_next_state[3]}), .Q ({data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1328, stateFF_state_gff_5_s_next_state[2]}), .Q ({data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1327, stateFF_state_gff_5_s_next_state[1]}), .Q ({data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1326, stateFF_state_gff_5_s_next_state[0]}), .Q ({data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1333, stateFF_state_gff_6_s_next_state[3]}), .Q ({data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1332, stateFF_state_gff_6_s_next_state[2]}), .Q ({data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1331, stateFF_state_gff_6_s_next_state[1]}), .Q ({data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1330, stateFF_state_gff_6_s_next_state[0]}), .Q ({data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1337, stateFF_state_gff_7_s_next_state[3]}), .Q ({data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1336, stateFF_state_gff_7_s_next_state[2]}), .Q ({data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1335, stateFF_state_gff_7_s_next_state[1]}), .Q ({data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1334, stateFF_state_gff_7_s_next_state[0]}), .Q ({data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1341, stateFF_state_gff_8_s_next_state[3]}), .Q ({data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1340, stateFF_state_gff_8_s_next_state[2]}), .Q ({data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1339, stateFF_state_gff_8_s_next_state[1]}), .Q ({data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1338, stateFF_state_gff_8_s_next_state[0]}), .Q ({data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1345, stateFF_state_gff_9_s_next_state[3]}), .Q ({data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1344, stateFF_state_gff_9_s_next_state[2]}), .Q ({data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1343, stateFF_state_gff_9_s_next_state[1]}), .Q ({data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1342, stateFF_state_gff_9_s_next_state[0]}), .Q ({data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1349, stateFF_state_gff_10_s_next_state[3]}), .Q ({data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1348, stateFF_state_gff_10_s_next_state[2]}), .Q ({data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1347, stateFF_state_gff_10_s_next_state[1]}), .Q ({data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1346, stateFF_state_gff_10_s_next_state[0]}), .Q ({data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1353, stateFF_state_gff_11_s_next_state[3]}), .Q ({data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1352, stateFF_state_gff_11_s_next_state[2]}), .Q ({data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1351, stateFF_state_gff_11_s_next_state[1]}), .Q ({data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1350, stateFF_state_gff_11_s_next_state[0]}), .Q ({data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1357, stateFF_state_gff_12_s_next_state[3]}), .Q ({data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1356, stateFF_state_gff_12_s_next_state[2]}), .Q ({data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1355, stateFF_state_gff_12_s_next_state[1]}), .Q ({data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1354, stateFF_state_gff_12_s_next_state[0]}), .Q ({data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1361, stateFF_state_gff_13_s_next_state[3]}), .Q ({data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1360, stateFF_state_gff_13_s_next_state[2]}), .Q ({data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1359, stateFF_state_gff_13_s_next_state[1]}), .Q ({data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1358, stateFF_state_gff_13_s_next_state[0]}), .Q ({data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1365, stateFF_state_gff_14_s_next_state[3]}), .Q ({data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1364, stateFF_state_gff_14_s_next_state[2]}), .Q ({data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1363, stateFF_state_gff_14_s_next_state[1]}), .Q ({data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1362, stateFF_state_gff_14_s_next_state[0]}), .Q ({data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1369, stateFF_state_gff_15_s_next_state[3]}), .Q ({data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1368, stateFF_state_gff_15_s_next_state[2]}), .Q ({data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1367, stateFF_state_gff_15_s_next_state[1]}), .Q ({data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1366, stateFF_state_gff_15_s_next_state[0]}), .Q ({data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1373, stateFF_state_gff_16_s_next_state[3]}), .Q ({data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1372, stateFF_state_gff_16_s_next_state[2]}), .Q ({data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1371, stateFF_state_gff_16_s_next_state[1]}), .Q ({data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateFF_state_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1370, stateFF_state_gff_16_s_next_state[0]}), .Q ({data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1377, keyFF_keystate_gff_1_s_next_state[3]}), .Q ({new_AGEMA_signal_1064, keyFF_outputPar[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1376, keyFF_keystate_gff_1_s_next_state[2]}), .Q ({new_AGEMA_signal_1291, keyRegKS[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1375, keyFF_keystate_gff_1_s_next_state[1]}), .Q ({new_AGEMA_signal_1289, keyRegKS[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1374, keyFF_keystate_gff_1_s_next_state[0]}), .Q ({new_AGEMA_signal_1287, keyRegKS[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1381, keyFF_keystate_gff_2_s_next_state[3]}), .Q ({new_AGEMA_signal_1076, keyFF_outputPar[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1380, keyFF_keystate_gff_2_s_next_state[2]}), .Q ({new_AGEMA_signal_1073, keyFF_outputPar[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1379, keyFF_keystate_gff_2_s_next_state[1]}), .Q ({new_AGEMA_signal_1070, keyFF_outputPar[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1378, keyFF_keystate_gff_2_s_next_state[0]}), .Q ({new_AGEMA_signal_1067, keyFF_outputPar[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1385, keyFF_keystate_gff_3_s_next_state[3]}), .Q ({new_AGEMA_signal_1088, keyFF_outputPar[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1384, keyFF_keystate_gff_3_s_next_state[2]}), .Q ({new_AGEMA_signal_1085, keyFF_outputPar[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1383, keyFF_keystate_gff_3_s_next_state[1]}), .Q ({new_AGEMA_signal_1082, keyFF_outputPar[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1382, keyFF_keystate_gff_3_s_next_state[0]}), .Q ({new_AGEMA_signal_1079, keyFF_outputPar[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1389, keyFF_keystate_gff_4_s_next_state[3]}), .Q ({new_AGEMA_signal_1100, keyFF_outputPar[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1388, keyFF_keystate_gff_4_s_next_state[2]}), .Q ({new_AGEMA_signal_1097, keyFF_outputPar[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1387, keyFF_keystate_gff_4_s_next_state[1]}), .Q ({new_AGEMA_signal_1094, keyFF_outputPar[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1386, keyFF_keystate_gff_4_s_next_state[0]}), .Q ({new_AGEMA_signal_1091, keyFF_outputPar[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1306, keyFF_keystate_gff_5_s_next_state[3]}), .Q ({new_AGEMA_signal_1274, keyFF_outputPar[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1305, keyFF_keystate_gff_5_s_next_state[2]}), .Q ({new_AGEMA_signal_1062, keyFF_outputPar[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1304, keyFF_keystate_gff_5_s_next_state[1]}), .Q ({new_AGEMA_signal_1106, keyFF_outputPar[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1303, keyFF_keystate_gff_5_s_next_state[0]}), .Q ({new_AGEMA_signal_1103, keyFF_outputPar[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1310, keyFF_keystate_gff_6_s_next_state[3]}), .Q ({new_AGEMA_signal_1109, keyFF_outputPar[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1309, keyFF_keystate_gff_6_s_next_state[2]}), .Q ({new_AGEMA_signal_1056, keyFF_outputPar[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1308, keyFF_keystate_gff_6_s_next_state[1]}), .Q ({new_AGEMA_signal_1058, keyFF_outputPar[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1307, keyFF_keystate_gff_6_s_next_state[0]}), .Q ({new_AGEMA_signal_1060, keyFF_outputPar[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1393, keyFF_keystate_gff_7_s_next_state[3]}), .Q ({new_AGEMA_signal_1121, keyFF_outputPar[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1392, keyFF_keystate_gff_7_s_next_state[2]}), .Q ({new_AGEMA_signal_1118, keyFF_outputPar[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1391, keyFF_keystate_gff_7_s_next_state[1]}), .Q ({new_AGEMA_signal_1115, keyFF_outputPar[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1390, keyFF_keystate_gff_7_s_next_state[0]}), .Q ({new_AGEMA_signal_1112, keyFF_outputPar[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1397, keyFF_keystate_gff_8_s_next_state[3]}), .Q ({new_AGEMA_signal_1133, keyFF_outputPar[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1396, keyFF_keystate_gff_8_s_next_state[2]}), .Q ({new_AGEMA_signal_1130, keyFF_outputPar[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1395, keyFF_keystate_gff_8_s_next_state[1]}), .Q ({new_AGEMA_signal_1127, keyFF_outputPar[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1394, keyFF_keystate_gff_8_s_next_state[0]}), .Q ({new_AGEMA_signal_1124, keyFF_outputPar[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1401, keyFF_keystate_gff_9_s_next_state[3]}), .Q ({new_AGEMA_signal_1145, keyFF_outputPar[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1400, keyFF_keystate_gff_9_s_next_state[2]}), .Q ({new_AGEMA_signal_1142, keyFF_outputPar[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1399, keyFF_keystate_gff_9_s_next_state[1]}), .Q ({new_AGEMA_signal_1139, keyFF_outputPar[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1398, keyFF_keystate_gff_9_s_next_state[0]}), .Q ({new_AGEMA_signal_1136, keyFF_outputPar[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1405, keyFF_keystate_gff_10_s_next_state[3]}), .Q ({new_AGEMA_signal_1157, keyFF_outputPar[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1404, keyFF_keystate_gff_10_s_next_state[2]}), .Q ({new_AGEMA_signal_1154, keyFF_outputPar[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1403, keyFF_keystate_gff_10_s_next_state[1]}), .Q ({new_AGEMA_signal_1151, keyFF_outputPar[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1402, keyFF_keystate_gff_10_s_next_state[0]}), .Q ({new_AGEMA_signal_1148, keyFF_outputPar[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1409, keyFF_keystate_gff_11_s_next_state[3]}), .Q ({new_AGEMA_signal_1169, keyFF_outputPar[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1408, keyFF_keystate_gff_11_s_next_state[2]}), .Q ({new_AGEMA_signal_1166, keyFF_outputPar[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1407, keyFF_keystate_gff_11_s_next_state[1]}), .Q ({new_AGEMA_signal_1163, keyFF_outputPar[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1406, keyFF_keystate_gff_11_s_next_state[0]}), .Q ({new_AGEMA_signal_1160, keyFF_outputPar[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1413, keyFF_keystate_gff_12_s_next_state[3]}), .Q ({new_AGEMA_signal_1181, keyFF_outputPar[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1412, keyFF_keystate_gff_12_s_next_state[2]}), .Q ({new_AGEMA_signal_1178, keyFF_outputPar[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1411, keyFF_keystate_gff_12_s_next_state[1]}), .Q ({new_AGEMA_signal_1175, keyFF_outputPar[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1410, keyFF_keystate_gff_12_s_next_state[0]}), .Q ({new_AGEMA_signal_1172, keyFF_outputPar[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1417, keyFF_keystate_gff_13_s_next_state[3]}), .Q ({new_AGEMA_signal_1193, keyFF_outputPar[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1416, keyFF_keystate_gff_13_s_next_state[2]}), .Q ({new_AGEMA_signal_1190, keyFF_outputPar[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1415, keyFF_keystate_gff_13_s_next_state[1]}), .Q ({new_AGEMA_signal_1187, keyFF_outputPar[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1414, keyFF_keystate_gff_13_s_next_state[0]}), .Q ({new_AGEMA_signal_1184, keyFF_outputPar[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1421, keyFF_keystate_gff_14_s_next_state[3]}), .Q ({new_AGEMA_signal_1205, keyFF_outputPar[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1420, keyFF_keystate_gff_14_s_next_state[2]}), .Q ({new_AGEMA_signal_1202, keyFF_outputPar[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1419, keyFF_keystate_gff_14_s_next_state[1]}), .Q ({new_AGEMA_signal_1199, keyFF_outputPar[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1418, keyFF_keystate_gff_14_s_next_state[0]}), .Q ({new_AGEMA_signal_1196, keyFF_outputPar[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1425, keyFF_keystate_gff_15_s_next_state[3]}), .Q ({new_AGEMA_signal_1217, keyFF_outputPar[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1424, keyFF_keystate_gff_15_s_next_state[2]}), .Q ({new_AGEMA_signal_1214, keyFF_outputPar[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1423, keyFF_keystate_gff_15_s_next_state[1]}), .Q ({new_AGEMA_signal_1211, keyFF_outputPar[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1422, keyFF_keystate_gff_15_s_next_state[0]}), .Q ({new_AGEMA_signal_1208, keyFF_outputPar[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1429, keyFF_keystate_gff_16_s_next_state[3]}), .Q ({new_AGEMA_signal_1229, keyFF_outputPar[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1428, keyFF_keystate_gff_16_s_next_state[2]}), .Q ({new_AGEMA_signal_1226, keyFF_outputPar[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1427, keyFF_keystate_gff_16_s_next_state[1]}), .Q ({new_AGEMA_signal_1223, keyFF_outputPar[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1426, keyFF_keystate_gff_16_s_next_state[0]}), .Q ({new_AGEMA_signal_1220, keyFF_outputPar[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1433, keyFF_keystate_gff_17_s_next_state[3]}), .Q ({new_AGEMA_signal_1241, keyFF_outputPar[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1432, keyFF_keystate_gff_17_s_next_state[2]}), .Q ({new_AGEMA_signal_1238, keyFF_outputPar[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1431, keyFF_keystate_gff_17_s_next_state[1]}), .Q ({new_AGEMA_signal_1235, keyFF_outputPar[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_17_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1430, keyFF_keystate_gff_17_s_next_state[0]}), .Q ({new_AGEMA_signal_1232, keyFF_outputPar[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1437, keyFF_keystate_gff_18_s_next_state[3]}), .Q ({new_AGEMA_signal_1253, keyFF_outputPar[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1436, keyFF_keystate_gff_18_s_next_state[2]}), .Q ({new_AGEMA_signal_1250, keyFF_outputPar[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1435, keyFF_keystate_gff_18_s_next_state[1]}), .Q ({new_AGEMA_signal_1247, keyFF_outputPar[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_18_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1434, keyFF_keystate_gff_18_s_next_state[0]}), .Q ({new_AGEMA_signal_1244, keyFF_outputPar[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1441, keyFF_keystate_gff_19_s_next_state[3]}), .Q ({new_AGEMA_signal_1265, keyFF_outputPar[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1440, keyFF_keystate_gff_19_s_next_state[2]}), .Q ({new_AGEMA_signal_1262, keyFF_outputPar[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1439, keyFF_keystate_gff_19_s_next_state[1]}), .Q ({new_AGEMA_signal_1259, keyFF_outputPar[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_19_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1438, keyFF_keystate_gff_19_s_next_state[0]}), .Q ({new_AGEMA_signal_1256, keyFF_outputPar[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1471, keyFF_keystate_gff_20_s_next_state[3]}), .Q ({new_AGEMA_signal_865, roundkey[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1466, keyFF_keystate_gff_20_s_next_state[2]}), .Q ({new_AGEMA_signal_862, roundkey[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1465, keyFF_keystate_gff_20_s_next_state[1]}), .Q ({new_AGEMA_signal_859, roundkey[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) keyFF_keystate_gff_20_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1448, keyFF_keystate_gff_20_s_next_state[0]}), .Q ({new_AGEMA_signal_856, roundkey[0]}) ) ;
endmodule
