/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_BDDcudd_ClockGating_d1 (SI_s0, clk, SI_s1, Fresh, rst, SO_s0, SO_s1, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input rst ;
    input [405:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output Synch ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_2169 ;

    /* cells in depth 0 */
    ClockGatingController #(17) cell_1333 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_2169 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_927 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_1341, signal_942}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_928 ( .s ({SI_s1[5], SI_s0[5]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_1343, signal_943}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_929 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_1345, signal_944}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_930 ( .s ({SI_s1[5], SI_s0[5]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_1346, signal_945}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_931 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_1347, signal_946}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_932 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1343, signal_943}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_1348, signal_947}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_933 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_1349, signal_948}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_934 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_1350, signal_949}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_935 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_1351, signal_950}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_936 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_1352, signal_951}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_937 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_1353, signal_952}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_938 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_1354, signal_953}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_939 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1343, signal_943}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_1355, signal_954}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_940 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_1356, signal_955}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_941 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_1357, signal_956}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_942 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_1358, signal_957}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_943 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_1359, signal_958}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_944 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_1360, signal_959}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_945 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_1361, signal_960}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_946 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1346, signal_945}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_1362, signal_961}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1346, signal_945}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_1363, signal_962}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_1364, signal_963}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_1365, signal_964}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_1366, signal_965}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_951 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_1367, signal_966}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_952 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_1368, signal_967}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_953 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1346, signal_945}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_1369, signal_968}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_954 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_1370, signal_969}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_955 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_1371, signal_970}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_956 ( .s ({SI_s1[2], SI_s0[2]}), .b ({signal_1343, signal_943}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_1372, signal_971}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_957 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_1373, signal_972}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_958 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_1374, signal_973}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_959 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_1375, signal_974}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_960 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_1376, signal_975}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_961 ( .s ({SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_1377, signal_976}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_962 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_1378, signal_977}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_963 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_1379, signal_978}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_1380, signal_979}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_965 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_1381, signal_980}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_1382, signal_981}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1341, signal_942}), .a ({signal_1353, signal_952}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_1384, signal_982}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_1385, signal_983}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_1386, signal_984}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_970 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_1387, signal_985}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_1388, signal_986}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_1389, signal_987}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_1390, signal_988}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_974 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_1391, signal_989}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_1392, signal_990}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_1393, signal_991}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_1394, signal_992}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_978 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_1395, signal_993}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_979 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_1396, signal_994}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_980 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_1397, signal_995}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_981 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_1398, signal_996}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_982 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_1399, signal_997}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_983 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_1400, signal_998}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_984 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_1401, signal_999}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_985 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_1402, signal_1000}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_986 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_1403, signal_1001}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_987 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_1404, signal_1002}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_988 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_1405, signal_1003}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_989 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_1406, signal_1004}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_990 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_1407, signal_1005}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_991 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_1408, signal_1006}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_992 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_1409, signal_1007}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_993 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_1410, signal_1008}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_994 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_1411, signal_1009}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_995 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_1412, signal_1010}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_996 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_1413, signal_1011}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_997 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_1414, signal_1012}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_998 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_1415, signal_1013}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_999 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1375, signal_974}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_1416, signal_1014}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1000 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1359, signal_958}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_1417, signal_1015}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1001 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_1418, signal_1016}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1002 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_1419, signal_1017}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1003 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_1420, signal_1018}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1004 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_1421, signal_1019}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1005 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_1422, signal_1020}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1006 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_1423, signal_1021}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1007 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_1424, signal_1022}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1008 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_1425, signal_1023}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1009 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_1426, signal_1024}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1010 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_1427, signal_1025}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1011 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_1428, signal_1026}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1012 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_1429, signal_1027}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1013 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_1430, signal_1028}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1014 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_1431, signal_1029}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1015 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[88] ), .c ({signal_1432, signal_1030}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1016 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[89] ), .c ({signal_1433, signal_1031}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1017 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[90] ), .c ({signal_1434, signal_1032}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1018 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[91] ), .c ({signal_1435, signal_1033}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1019 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[92] ), .c ({signal_1436, signal_1034}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1020 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1376, signal_975}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[93] ), .c ({signal_1437, signal_1035}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1021 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[94] ), .c ({signal_1438, signal_1036}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1022 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1350, signal_949}), .a ({signal_1373, signal_972}), .clk ( clk ), .r ( Fresh[95] ), .c ({signal_1439, signal_1037}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1023 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[96] ), .c ({signal_1440, signal_1038}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1024 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[97] ), .c ({signal_1441, signal_1039}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1025 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[98] ), .c ({signal_1442, signal_1040}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1026 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[99] ), .c ({signal_1443, signal_1041}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1027 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1361, signal_960}), .a ({signal_1354, signal_953}), .clk ( clk ), .r ( Fresh[100] ), .c ({signal_1444, signal_1042}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1028 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[101] ), .c ({signal_1445, signal_1043}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1029 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[102] ), .c ({signal_1446, signal_1044}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1030 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1355, signal_954}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[103] ), .c ({signal_1447, signal_1045}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1031 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[104] ), .c ({signal_1448, signal_1046}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1032 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[105] ), .c ({signal_1449, signal_1047}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1033 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[106] ), .c ({signal_1450, signal_1048}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1034 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[107] ), .c ({signal_1451, signal_1049}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1035 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[108] ), .c ({signal_1452, signal_1050}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1036 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[109] ), .c ({signal_1453, signal_1051}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1037 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[110] ), .c ({signal_1454, signal_1052}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1038 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[111] ), .c ({signal_1455, signal_1053}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1039 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[112] ), .c ({signal_1456, signal_1054}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1040 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[113] ), .c ({signal_1457, signal_1055}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1041 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[114] ), .c ({signal_1458, signal_1056}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1042 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[115] ), .c ({signal_1459, signal_1057}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1043 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[116] ), .c ({signal_1460, signal_1058}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1044 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[117] ), .c ({signal_1461, signal_1059}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1045 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[118] ), .c ({signal_1462, signal_1060}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1046 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[119] ), .c ({signal_1463, signal_1061}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1047 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[120] ), .c ({signal_1464, signal_1062}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1048 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[121] ), .c ({signal_1465, signal_1063}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1049 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[122] ), .c ({signal_1466, signal_1064}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1050 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[123] ), .c ({signal_1467, signal_1065}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1051 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[124] ), .c ({signal_1468, signal_1066}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1052 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[125] ), .c ({signal_1469, signal_1067}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1053 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[126] ), .c ({signal_1470, signal_1068}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1054 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[127] ), .c ({signal_1471, signal_1069}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1055 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1346, signal_945}), .clk ( clk ), .r ( Fresh[128] ), .c ({signal_1472, signal_1070}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1056 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[129] ), .c ({signal_1473, signal_1071}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1057 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[130] ), .c ({signal_1474, signal_1072}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1058 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b0}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[131] ), .c ({signal_1475, signal_1073}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1059 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[132] ), .c ({signal_1476, signal_1074}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1060 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[133] ), .c ({signal_1477, signal_1075}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1061 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[134] ), .c ({signal_1478, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1062 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[135] ), .c ({signal_1479, signal_1077}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1063 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1362, signal_961}), .clk ( clk ), .r ( Fresh[136] ), .c ({signal_1480, signal_1078}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1064 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[137] ), .c ({signal_1481, signal_1079}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1065 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1345, signal_944}), .clk ( clk ), .r ( Fresh[138] ), .c ({signal_1482, signal_1080}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1066 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[139] ), .c ({signal_1483, signal_1081}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1067 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[140] ), .c ({signal_1484, signal_1082}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1068 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1348, signal_947}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[141] ), .c ({signal_1485, signal_1083}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1069 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[142] ), .c ({signal_1486, signal_1084}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1070 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1375, signal_974}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[143] ), .c ({signal_1487, signal_1085}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1071 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[144] ), .c ({signal_1488, signal_1086}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1072 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1371, signal_970}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[145] ), .c ({signal_1489, signal_1087}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1073 ( .s ({SI_s1[4], SI_s0[4]}), .b ({1'b0, 1'b1}), .a ({signal_1377, signal_976}), .clk ( clk ), .r ( Fresh[146] ), .c ({signal_1490, signal_1088}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1074 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1372, signal_971}), .clk ( clk ), .r ( Fresh[147] ), .c ({signal_1491, signal_1089}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1369, signal_968}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[148] ), .c ({signal_1492, signal_1090}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[149] ), .c ({signal_1493, signal_1091}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[150] ), .c ({signal_1494, signal_1092}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[151] ), .c ({signal_1495, signal_1093}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1363, signal_962}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[152] ), .c ({signal_1496, signal_1094}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[153] ), .c ({signal_1497, signal_1095}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1345, signal_944}), .a ({signal_1371, signal_970}), .clk ( clk ), .r ( Fresh[154] ), .c ({signal_1498, signal_1096}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[155] ), .c ({signal_1499, signal_1097}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[156] ), .c ({signal_1500, signal_1098}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1346, signal_945}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[157] ), .c ({signal_1501, signal_1099}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1361, signal_960}), .a ({signal_1375, signal_974}), .clk ( clk ), .r ( Fresh[158] ), .c ({signal_1502, signal_1100}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1377, signal_976}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[159] ), .c ({signal_1503, signal_1101}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1347, signal_946}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[160] ), .c ({signal_1504, signal_1102}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1362, signal_961}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[161] ), .c ({signal_1505, signal_1103}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1343, signal_943}), .a ({signal_1363, signal_962}), .clk ( clk ), .r ( Fresh[162] ), .c ({signal_1506, signal_1104}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .s ({SI_s1[4], SI_s0[4]}), .b ({signal_1372, signal_971}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[163] ), .c ({signal_1507, signal_1105}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1091 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1440, signal_1038}), .a ({signal_1420, signal_1018}), .clk ( clk ), .r ( Fresh[164] ), .c ({signal_1508, signal_1106}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1092 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1395, signal_993}), .a ({signal_1404, signal_1002}), .clk ( clk ), .r ( Fresh[165] ), .c ({signal_1509, signal_1107}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1093 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1438, signal_1036}), .a ({signal_1394, signal_992}), .clk ( clk ), .r ( Fresh[166] ), .c ({signal_1510, signal_1108}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1094 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1462, signal_1060}), .a ({signal_1366, signal_965}), .clk ( clk ), .r ( Fresh[167] ), .c ({signal_1511, signal_1109}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1468, signal_1066}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[168] ), .c ({signal_1512, signal_1110}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1365, signal_964}), .a ({signal_1428, signal_1026}), .clk ( clk ), .r ( Fresh[169] ), .c ({signal_1513, signal_1111}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1369, signal_968}), .a ({signal_1507, signal_1105}), .clk ( clk ), .r ( Fresh[170] ), .c ({signal_1514, signal_1112}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1457, signal_1055}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[171] ), .c ({signal_1515, signal_1113}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1491, signal_1089}), .a ({signal_1483, signal_1081}), .clk ( clk ), .r ( Fresh[172] ), .c ({signal_1516, signal_1114}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1357, signal_956}), .a ({signal_1441, signal_1039}), .clk ( clk ), .r ( Fresh[173] ), .c ({signal_1517, signal_1115}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1396, signal_994}), .a ({signal_1394, signal_992}), .clk ( clk ), .r ( Fresh[174] ), .c ({signal_1518, signal_1116}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1364, signal_963}), .a ({signal_1470, signal_1068}), .clk ( clk ), .r ( Fresh[175] ), .c ({signal_1519, signal_1117}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1403, signal_1001}), .a ({signal_1461, signal_1059}), .clk ( clk ), .r ( Fresh[176] ), .c ({signal_1520, signal_1118}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1460, signal_1058}), .a ({signal_1465, signal_1063}), .clk ( clk ), .r ( Fresh[177] ), .c ({signal_1521, signal_1119}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1445, signal_1043}), .a ({signal_1351, signal_950}), .clk ( clk ), .r ( Fresh[178] ), .c ({signal_1522, signal_1120}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1341, signal_942}), .a ({signal_1435, signal_1033}), .clk ( clk ), .r ( Fresh[179] ), .c ({signal_1523, signal_1121}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1107 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1459, signal_1057}), .a ({signal_1480, signal_1078}), .clk ( clk ), .r ( Fresh[180] ), .c ({signal_1524, signal_1122}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1108 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1445, signal_1043}), .a ({signal_1400, signal_998}), .clk ( clk ), .r ( Fresh[181] ), .c ({signal_1525, signal_1123}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1109 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1413, signal_1011}), .a ({signal_1359, signal_958}), .clk ( clk ), .r ( Fresh[182] ), .c ({signal_1526, signal_1124}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1110 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1397, signal_995}), .a ({signal_1471, signal_1069}), .clk ( clk ), .r ( Fresh[183] ), .c ({signal_1527, signal_1125}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1111 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1483, signal_1081}), .a ({signal_1505, signal_1103}), .clk ( clk ), .r ( Fresh[184] ), .c ({signal_1528, signal_1126}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1112 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1404, signal_1002}), .a ({signal_1458, signal_1056}), .clk ( clk ), .r ( Fresh[185] ), .c ({signal_1529, signal_1127}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1113 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1497, signal_1095}), .a ({signal_1478, signal_1076}), .clk ( clk ), .r ( Fresh[186] ), .c ({signal_1530, signal_1128}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1114 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1482, signal_1080}), .a ({signal_1449, signal_1047}), .clk ( clk ), .r ( Fresh[187] ), .c ({signal_1531, signal_1129}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1115 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1410, signal_1008}), .a ({signal_1424, signal_1022}), .clk ( clk ), .r ( Fresh[188] ), .c ({signal_1532, signal_1130}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1116 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1485, signal_1083}), .a ({signal_1477, signal_1075}), .clk ( clk ), .r ( Fresh[189] ), .c ({signal_1533, signal_1131}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1117 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1419, signal_1017}), .a ({signal_1431, signal_1029}), .clk ( clk ), .r ( Fresh[190] ), .c ({signal_1534, signal_1132}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1118 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1488, signal_1086}), .a ({signal_1467, signal_1065}), .clk ( clk ), .r ( Fresh[191] ), .c ({signal_1535, signal_1133}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1119 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1385, signal_983}), .a ({signal_1488, signal_1086}), .clk ( clk ), .r ( Fresh[192] ), .c ({signal_1536, signal_1134}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1120 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1504, signal_1102}), .a ({signal_1357, signal_956}), .clk ( clk ), .r ( Fresh[193] ), .c ({signal_1537, signal_1135}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1121 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1451, signal_1049}), .a ({signal_1386, signal_984}), .clk ( clk ), .r ( Fresh[194] ), .c ({signal_1538, signal_1136}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1122 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1473, signal_1071}), .a ({signal_1442, signal_1040}), .clk ( clk ), .r ( Fresh[195] ), .c ({signal_1539, signal_1137}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1123 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1429, signal_1027}), .a ({signal_1443, signal_1041}), .clk ( clk ), .r ( Fresh[196] ), .c ({signal_1540, signal_1138}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1124 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1418, signal_1016}), .a ({signal_1466, signal_1064}), .clk ( clk ), .r ( Fresh[197] ), .c ({signal_1541, signal_1139}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1125 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1374, signal_973}), .a ({signal_1427, signal_1025}), .clk ( clk ), .r ( Fresh[198] ), .c ({signal_1542, signal_1140}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1126 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1401, signal_999}), .a ({signal_1498, signal_1096}), .clk ( clk ), .r ( Fresh[199] ), .c ({signal_1543, signal_1141}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1127 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1489, signal_1087}), .a ({signal_1498, signal_1096}), .clk ( clk ), .r ( Fresh[200] ), .c ({signal_1544, signal_1142}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1128 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1391, signal_989}), .a ({signal_1390, signal_988}), .clk ( clk ), .r ( Fresh[201] ), .c ({signal_1545, signal_1143}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1129 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1499, signal_1097}), .a ({signal_1468, signal_1066}), .clk ( clk ), .r ( Fresh[202] ), .c ({signal_1546, signal_1144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1130 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1407, signal_1005}), .a ({signal_1440, signal_1038}), .clk ( clk ), .r ( Fresh[203] ), .c ({signal_1547, signal_1145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1131 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1458, signal_1056}), .a ({signal_1447, signal_1045}), .clk ( clk ), .r ( Fresh[204] ), .c ({signal_1548, signal_1146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1132 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1449, signal_1047}), .a ({signal_1393, signal_991}), .clk ( clk ), .r ( Fresh[205] ), .c ({signal_1549, signal_1147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1133 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1389, signal_987}), .a ({signal_1387, signal_985}), .clk ( clk ), .r ( Fresh[206] ), .c ({signal_1550, signal_1148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1134 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1491, signal_1089}), .a ({signal_1395, signal_993}), .clk ( clk ), .r ( Fresh[207] ), .c ({signal_1551, signal_1149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1135 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1421, signal_1019}), .a ({signal_1471, signal_1069}), .clk ( clk ), .r ( Fresh[208] ), .c ({signal_1552, signal_1150}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1136 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1490, signal_1088}), .a ({signal_1378, signal_977}), .clk ( clk ), .r ( Fresh[209] ), .c ({signal_1553, signal_1151}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1137 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1341, signal_942}), .a ({signal_1430, signal_1028}), .clk ( clk ), .r ( Fresh[210] ), .c ({signal_1554, signal_1152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1138 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1421, signal_1019}), .a ({signal_1385, signal_983}), .clk ( clk ), .r ( Fresh[211] ), .c ({signal_1555, signal_1153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1407, signal_1005}), .a ({signal_1412, signal_1010}), .clk ( clk ), .r ( Fresh[212] ), .c ({signal_1556, signal_1154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1438, signal_1036}), .a ({signal_1450, signal_1048}), .clk ( clk ), .r ( Fresh[213] ), .c ({signal_1557, signal_1155}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1463, signal_1061}), .a ({signal_1464, signal_1062}), .clk ( clk ), .r ( Fresh[214] ), .c ({signal_1558, signal_1156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1492, signal_1090}), .a ({signal_1435, signal_1033}), .clk ( clk ), .r ( Fresh[215] ), .c ({signal_1559, signal_1157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1486, signal_1084}), .a ({signal_1412, signal_1010}), .clk ( clk ), .r ( Fresh[216] ), .c ({signal_1560, signal_1158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1490, signal_1088}), .a ({signal_1355, signal_954}), .clk ( clk ), .r ( Fresh[217] ), .c ({signal_1561, signal_1159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1506, signal_1104}), .a ({signal_1414, signal_1012}), .clk ( clk ), .r ( Fresh[218] ), .c ({signal_1562, signal_1160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1474, signal_1072}), .a ({signal_1500, signal_1098}), .clk ( clk ), .r ( Fresh[219] ), .c ({signal_1563, signal_1161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1445, signal_1043}), .a ({signal_1361, signal_960}), .clk ( clk ), .r ( Fresh[220] ), .c ({signal_1564, signal_1162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1458, signal_1056}), .a ({signal_1481, signal_1079}), .clk ( clk ), .r ( Fresh[221] ), .c ({signal_1565, signal_1163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1418, signal_1016}), .a ({signal_1452, signal_1050}), .clk ( clk ), .r ( Fresh[222] ), .c ({signal_1566, signal_1164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1490, signal_1088}), .a ({signal_1477, signal_1075}), .clk ( clk ), .r ( Fresh[223] ), .c ({signal_1567, signal_1165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1415, signal_1013}), .a ({signal_1442, signal_1040}), .clk ( clk ), .r ( Fresh[224] ), .c ({signal_1568, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1449, signal_1047}), .a ({signal_1445, signal_1043}), .clk ( clk ), .r ( Fresh[225] ), .c ({signal_1569, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1396, signal_994}), .a ({signal_1503, signal_1101}), .clk ( clk ), .r ( Fresh[226] ), .c ({signal_1570, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1393, signal_991}), .a ({signal_1470, signal_1068}), .clk ( clk ), .r ( Fresh[227] ), .c ({signal_1571, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1411, signal_1009}), .a ({signal_1484, signal_1082}), .clk ( clk ), .r ( Fresh[228] ), .c ({signal_1572, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1405, signal_1003}), .a ({signal_1479, signal_1077}), .clk ( clk ), .r ( Fresh[229] ), .c ({signal_1573, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1456, signal_1054}), .a ({signal_1476, signal_1074}), .clk ( clk ), .r ( Fresh[230] ), .c ({signal_1574, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1480, signal_1078}), .a ({signal_1484, signal_1082}), .clk ( clk ), .r ( Fresh[231] ), .c ({signal_1575, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1424, signal_1022}), .a ({signal_1351, signal_950}), .clk ( clk ), .r ( Fresh[232] ), .c ({signal_1576, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1349, signal_948}), .a ({signal_1434, signal_1032}), .clk ( clk ), .r ( Fresh[233] ), .c ({signal_1577, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1432, signal_1030}), .a ({signal_1393, signal_991}), .clk ( clk ), .r ( Fresh[234] ), .c ({signal_1578, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1414, signal_1012}), .a ({signal_1469, signal_1067}), .clk ( clk ), .r ( Fresh[235] ), .c ({signal_1579, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1352, signal_951}), .a ({signal_1504, signal_1102}), .clk ( clk ), .r ( Fresh[236] ), .c ({signal_1580, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1463, signal_1061}), .a ({signal_1494, signal_1092}), .clk ( clk ), .r ( Fresh[237] ), .c ({signal_1581, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1472, signal_1070}), .a ({signal_1370, signal_969}), .clk ( clk ), .r ( Fresh[238] ), .c ({signal_1582, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1362, signal_961}), .a ({signal_1400, signal_998}), .clk ( clk ), .r ( Fresh[239] ), .c ({signal_1583, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1389, signal_987}), .a ({signal_1366, signal_965}), .clk ( clk ), .r ( Fresh[240] ), .c ({signal_1584, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1406, signal_1004}), .a ({signal_1368, signal_967}), .clk ( clk ), .r ( Fresh[241] ), .c ({signal_1585, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1396, signal_994}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[242] ), .c ({signal_1586, signal_1184}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1407, signal_1005}), .a ({signal_1368, signal_967}), .clk ( clk ), .r ( Fresh[243] ), .c ({signal_1587, signal_1185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1464, signal_1062}), .a ({signal_1341, signal_942}), .clk ( clk ), .r ( Fresh[244] ), .c ({signal_1588, signal_1186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1363, signal_962}), .a ({signal_1496, signal_1094}), .clk ( clk ), .r ( Fresh[245] ), .c ({signal_1589, signal_1187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1499, signal_1097}), .a ({signal_1399, signal_997}), .clk ( clk ), .r ( Fresh[246] ), .c ({signal_1590, signal_1188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1468, signal_1066}), .a ({signal_1401, signal_999}), .clk ( clk ), .r ( Fresh[247] ), .c ({signal_1591, signal_1189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1433, signal_1031}), .a ({signal_1453, signal_1051}), .clk ( clk ), .r ( Fresh[248] ), .c ({signal_1592, signal_1190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1448, signal_1046}), .a ({signal_1409, signal_1007}), .clk ( clk ), .r ( Fresh[249] ), .c ({signal_1593, signal_1191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1479, signal_1077}), .a ({signal_1343, signal_943}), .clk ( clk ), .r ( Fresh[250] ), .c ({signal_1594, signal_1192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1382, signal_981}), .a ({signal_1408, signal_1006}), .clk ( clk ), .r ( Fresh[251] ), .c ({signal_1595, signal_1193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1357, signal_956}), .a ({signal_1392, signal_990}), .clk ( clk ), .r ( Fresh[252] ), .c ({signal_1596, signal_1194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1367, signal_966}), .a ({signal_1449, signal_1047}), .clk ( clk ), .r ( Fresh[253] ), .c ({signal_1597, signal_1195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1475, signal_1073}), .a ({signal_1426, signal_1024}), .clk ( clk ), .r ( Fresh[254] ), .c ({signal_1598, signal_1196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1392, signal_990}), .a ({signal_1421, signal_1019}), .clk ( clk ), .r ( Fresh[255] ), .c ({signal_1599, signal_1197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1414, signal_1012}), .a ({signal_1411, signal_1009}), .clk ( clk ), .r ( Fresh[256] ), .c ({signal_1600, signal_1198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1446, signal_1044}), .a ({signal_1436, signal_1034}), .clk ( clk ), .r ( Fresh[257] ), .c ({signal_1601, signal_1199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1493, signal_1091}), .a ({signal_1455, signal_1053}), .clk ( clk ), .r ( Fresh[258] ), .c ({signal_1602, signal_1200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1493, signal_1091}), .a ({signal_1347, signal_946}), .clk ( clk ), .r ( Fresh[259] ), .c ({signal_1603, signal_1201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1433, signal_1031}), .a ({signal_1496, signal_1094}), .clk ( clk ), .r ( Fresh[260] ), .c ({signal_1604, signal_1202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1397, signal_995}), .a ({signal_1419, signal_1017}), .clk ( clk ), .r ( Fresh[261] ), .c ({signal_1605, signal_1203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1453, signal_1051}), .a ({signal_1456, signal_1054}), .clk ( clk ), .r ( Fresh[262] ), .c ({signal_1606, signal_1204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1396, signal_994}), .a ({signal_1493, signal_1091}), .clk ( clk ), .r ( Fresh[263] ), .c ({signal_1607, signal_1205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1487, signal_1085}), .a ({signal_1369, signal_968}), .clk ( clk ), .r ( Fresh[264] ), .c ({signal_1608, signal_1206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1376, signal_975}), .a ({signal_1425, signal_1023}), .clk ( clk ), .r ( Fresh[265] ), .c ({signal_1609, signal_1207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1360, signal_959}), .a ({signal_1495, signal_1093}), .clk ( clk ), .r ( Fresh[266] ), .c ({signal_1610, signal_1208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1454, signal_1052}), .a ({signal_1410, signal_1008}), .clk ( clk ), .r ( Fresh[267] ), .c ({signal_1611, signal_1209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1356, signal_955}), .a ({signal_1418, signal_1016}), .clk ( clk ), .r ( Fresh[268] ), .c ({signal_1612, signal_1210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1393, signal_991}), .a ({signal_1348, signal_947}), .clk ( clk ), .r ( Fresh[269] ), .c ({signal_1613, signal_1211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1503, signal_1101}), .a ({signal_1461, signal_1059}), .clk ( clk ), .r ( Fresh[270] ), .c ({signal_1614, signal_1212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1423, signal_1021}), .a ({signal_1471, signal_1069}), .clk ( clk ), .r ( Fresh[271] ), .c ({signal_1615, signal_1213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1387, signal_985}), .a ({signal_1379, signal_978}), .clk ( clk ), .r ( Fresh[272] ), .c ({signal_1616, signal_1214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1502, signal_1100}), .a ({signal_1449, signal_1047}), .clk ( clk ), .r ( Fresh[273] ), .c ({signal_1617, signal_1215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1358, signal_957}), .a ({signal_1405, signal_1003}), .clk ( clk ), .r ( Fresh[274] ), .c ({signal_1618, signal_1216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1445, signal_1043}), .a ({signal_1402, signal_1000}), .clk ( clk ), .r ( Fresh[275] ), .c ({signal_1619, signal_1217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1388, signal_986}), .a ({signal_1350, signal_949}), .clk ( clk ), .r ( Fresh[276] ), .c ({signal_1620, signal_1218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1390, signal_988}), .a ({signal_1501, signal_1099}), .clk ( clk ), .r ( Fresh[277] ), .c ({signal_1621, signal_1219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1403, signal_1001}), .a ({signal_1380, signal_979}), .clk ( clk ), .r ( Fresh[278] ), .c ({signal_1622, signal_1220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1447, signal_1045}), .a ({signal_1422, signal_1020}), .clk ( clk ), .r ( Fresh[279] ), .c ({signal_1623, signal_1221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1436, signal_1034}), .a ({signal_1398, signal_996}), .clk ( clk ), .r ( Fresh[280] ), .c ({signal_1624, signal_1222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .s ({SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0}), .a ({signal_1381, signal_980}), .clk ( clk ), .r ( Fresh[281] ), .c ({signal_1625, signal_1223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1463, signal_1061}), .a ({signal_1498, signal_1096}), .clk ( clk ), .r ( Fresh[282] ), .c ({signal_1626, signal_1224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1484, signal_1082}), .a ({signal_1455, signal_1053}), .clk ( clk ), .r ( Fresh[283] ), .c ({signal_1627, signal_1225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1401, signal_999}), .a ({signal_1351, signal_950}), .clk ( clk ), .r ( Fresh[284] ), .c ({signal_1628, signal_1226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .s ({SI_s1[1], SI_s0[1]}), .b ({signal_1343, signal_943}), .a ({signal_1400, signal_998}), .clk ( clk ), .r ( Fresh[285] ), .c ({signal_1629, signal_1227}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1587, signal_1185}), .a ({signal_1624, signal_1222}), .clk ( clk ), .r ( Fresh[286] ), .c ({signal_1631, signal_1228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1618, signal_1216}), .a ({signal_1595, signal_1193}), .clk ( clk ), .r ( Fresh[287] ), .c ({signal_1632, signal_1229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1215 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1563, signal_1161}), .a ({signal_1518, signal_1116}), .clk ( clk ), .r ( Fresh[288] ), .c ({signal_1633, signal_1230}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1216 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1617, signal_1215}), .a ({signal_1585, signal_1183}), .clk ( clk ), .r ( Fresh[289] ), .c ({signal_1634, signal_1231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1217 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1444, signal_1042}), .a ({signal_1544, signal_1142}), .clk ( clk ), .r ( Fresh[290] ), .c ({signal_1635, signal_1232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1218 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1580, signal_1178}), .a ({signal_1612, signal_1210}), .clk ( clk ), .r ( Fresh[291] ), .c ({signal_1636, signal_1233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1219 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1553, signal_1151}), .a ({signal_1557, signal_1155}), .clk ( clk ), .r ( Fresh[292] ), .c ({signal_1637, signal_1234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1220 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1546, signal_1144}), .a ({signal_1613, signal_1211}), .clk ( clk ), .r ( Fresh[293] ), .c ({signal_1638, signal_1235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1221 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1559, signal_1157}), .a ({signal_1600, signal_1198}), .clk ( clk ), .r ( Fresh[294] ), .c ({signal_1639, signal_1236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1222 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1525, signal_1123}), .a ({signal_1543, signal_1141}), .clk ( clk ), .r ( Fresh[295] ), .c ({signal_1640, signal_1237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1223 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1586, signal_1184}), .a ({signal_1524, signal_1122}), .clk ( clk ), .r ( Fresh[296] ), .c ({signal_1641, signal_1238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1224 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1561, signal_1159}), .a ({signal_1515, signal_1113}), .clk ( clk ), .r ( Fresh[297] ), .c ({signal_1642, signal_1239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1225 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1537, signal_1135}), .a ({signal_1522, signal_1120}), .clk ( clk ), .r ( Fresh[298] ), .c ({signal_1643, signal_1240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1226 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1545, signal_1143}), .a ({signal_1527, signal_1125}), .clk ( clk ), .r ( Fresh[299] ), .c ({signal_1644, signal_1241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1227 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1599, signal_1197}), .a ({signal_1531, signal_1129}), .clk ( clk ), .r ( Fresh[300] ), .c ({signal_1645, signal_1242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1228 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1581, signal_1179}), .a ({signal_1567, signal_1165}), .clk ( clk ), .r ( Fresh[301] ), .c ({signal_1646, signal_1243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1229 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1614, signal_1212}), .a ({signal_1628, signal_1226}), .clk ( clk ), .r ( Fresh[302] ), .c ({signal_1647, signal_1244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1230 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1517, signal_1115}), .a ({signal_1555, signal_1153}), .clk ( clk ), .r ( Fresh[303] ), .c ({signal_1648, signal_1245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1231 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1568, signal_1166}), .a ({signal_1416, signal_1014}), .clk ( clk ), .r ( Fresh[304] ), .c ({signal_1649, signal_1246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1232 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1542, signal_1140}), .a ({signal_1619, signal_1217}), .clk ( clk ), .r ( Fresh[305] ), .c ({signal_1650, signal_1247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1233 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1592, signal_1190}), .a ({signal_1437, signal_1035}), .clk ( clk ), .r ( Fresh[306] ), .c ({signal_1651, signal_1248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1234 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1558, signal_1156}), .a ({signal_1593, signal_1191}), .clk ( clk ), .r ( Fresh[307] ), .c ({signal_1652, signal_1249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1235 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1520, signal_1118}), .a ({signal_1511, signal_1109}), .clk ( clk ), .r ( Fresh[308] ), .c ({signal_1653, signal_1250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1236 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1594, signal_1192}), .a ({signal_1548, signal_1146}), .clk ( clk ), .r ( Fresh[309] ), .c ({signal_1654, signal_1251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1237 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1596, signal_1194}), .a ({signal_1540, signal_1138}), .clk ( clk ), .r ( Fresh[310] ), .c ({signal_1655, signal_1252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1238 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1590, signal_1188}), .a ({signal_1508, signal_1106}), .clk ( clk ), .r ( Fresh[311] ), .c ({signal_1656, signal_1253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1239 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1582, signal_1180}), .a ({signal_1562, signal_1160}), .clk ( clk ), .r ( Fresh[312] ), .c ({signal_1657, signal_1254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1240 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1529, signal_1127}), .a ({signal_1616, signal_1214}), .clk ( clk ), .r ( Fresh[313] ), .c ({signal_1658, signal_1255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1241 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1584, signal_1182}), .a ({signal_1541, signal_1139}), .clk ( clk ), .r ( Fresh[314] ), .c ({signal_1659, signal_1256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1242 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1579, signal_1177}), .a ({signal_1551, signal_1149}), .clk ( clk ), .r ( Fresh[315] ), .c ({signal_1660, signal_1257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1243 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1575, signal_1173}), .a ({signal_1523, signal_1121}), .clk ( clk ), .r ( Fresh[316] ), .c ({signal_1661, signal_1258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1244 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1589, signal_1187}), .a ({signal_1519, signal_1117}), .clk ( clk ), .r ( Fresh[317] ), .c ({signal_1662, signal_1259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1245 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1513, signal_1111}), .a ({signal_1560, signal_1158}), .clk ( clk ), .r ( Fresh[318] ), .c ({signal_1663, signal_1260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1246 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1384, signal_982}), .a ({signal_1509, signal_1107}), .clk ( clk ), .r ( Fresh[319] ), .c ({signal_1664, signal_1261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1247 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1556, signal_1154}), .a ({signal_1622, signal_1220}), .clk ( clk ), .r ( Fresh[320] ), .c ({signal_1665, signal_1262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1248 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1530, signal_1128}), .a ({signal_1521, signal_1119}), .clk ( clk ), .r ( Fresh[321] ), .c ({signal_1666, signal_1263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1249 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1533, signal_1131}), .a ({signal_1604, signal_1202}), .clk ( clk ), .r ( Fresh[322] ), .c ({signal_1667, signal_1264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1250 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1569, signal_1167}), .a ({signal_1554, signal_1152}), .clk ( clk ), .r ( Fresh[323] ), .c ({signal_1668, signal_1265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1251 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1591, signal_1189}), .a ({signal_1606, signal_1204}), .clk ( clk ), .r ( Fresh[324] ), .c ({signal_1669, signal_1266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1252 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1552, signal_1150}), .a ({signal_1610, signal_1208}), .clk ( clk ), .r ( Fresh[325] ), .c ({signal_1670, signal_1267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1253 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1578, signal_1176}), .a ({signal_1535, signal_1133}), .clk ( clk ), .r ( Fresh[326] ), .c ({signal_1671, signal_1268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1254 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1621, signal_1219}), .a ({signal_1607, signal_1205}), .clk ( clk ), .r ( Fresh[327] ), .c ({signal_1672, signal_1269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1255 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1577, signal_1175}), .a ({signal_1532, signal_1130}), .clk ( clk ), .r ( Fresh[328] ), .c ({signal_1673, signal_1270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1256 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1550, signal_1148}), .a ({signal_1570, signal_1168}), .clk ( clk ), .r ( Fresh[329] ), .c ({signal_1674, signal_1271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1257 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1597, signal_1195}), .a ({signal_1538, signal_1136}), .clk ( clk ), .r ( Fresh[330] ), .c ({signal_1675, signal_1272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1258 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1605, signal_1203}), .a ({signal_1598, signal_1196}), .clk ( clk ), .r ( Fresh[331] ), .c ({signal_1676, signal_1273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1259 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1528, signal_1126}), .a ({signal_1601, signal_1199}), .clk ( clk ), .r ( Fresh[332] ), .c ({signal_1677, signal_1274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1260 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1539, signal_1137}), .a ({signal_1611, signal_1209}), .clk ( clk ), .r ( Fresh[333] ), .c ({signal_1678, signal_1275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1261 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1608, signal_1206}), .a ({signal_1571, signal_1169}), .clk ( clk ), .r ( Fresh[334] ), .c ({signal_1679, signal_1276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1262 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1603, signal_1201}), .a ({signal_1623, signal_1221}), .clk ( clk ), .r ( Fresh[335] ), .c ({signal_1680, signal_1277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1263 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1625, signal_1223}), .a ({signal_1514, signal_1112}), .clk ( clk ), .r ( Fresh[336] ), .c ({signal_1681, signal_1278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1264 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1572, signal_1170}), .a ({signal_1564, signal_1162}), .clk ( clk ), .r ( Fresh[337] ), .c ({signal_1682, signal_1279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1265 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1439, signal_1037}), .a ({signal_1512, signal_1110}), .clk ( clk ), .r ( Fresh[338] ), .c ({signal_1683, signal_1280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1266 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1626, signal_1224}), .a ({signal_1620, signal_1218}), .clk ( clk ), .r ( Fresh[339] ), .c ({signal_1684, signal_1281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1267 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1549, signal_1147}), .a ({signal_1510, signal_1108}), .clk ( clk ), .r ( Fresh[340] ), .c ({signal_1685, signal_1282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1268 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1534, signal_1132}), .a ({signal_1565, signal_1163}), .clk ( clk ), .r ( Fresh[341] ), .c ({signal_1686, signal_1283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1269 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1627, signal_1225}), .a ({signal_1526, signal_1124}), .clk ( clk ), .r ( Fresh[342] ), .c ({signal_1687, signal_1284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1270 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1417, signal_1015}), .a ({signal_1588, signal_1186}), .clk ( clk ), .r ( Fresh[343] ), .c ({signal_1688, signal_1285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1271 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1609, signal_1207}), .a ({signal_1602, signal_1200}), .clk ( clk ), .r ( Fresh[344] ), .c ({signal_1689, signal_1286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1272 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1629, signal_1227}), .a ({signal_1574, signal_1172}), .clk ( clk ), .r ( Fresh[345] ), .c ({signal_1690, signal_1287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1273 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1576, signal_1174}), .a ({signal_1573, signal_1171}), .clk ( clk ), .r ( Fresh[346] ), .c ({signal_1691, signal_1288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1274 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1536, signal_1134}), .a ({signal_1583, signal_1181}), .clk ( clk ), .r ( Fresh[347] ), .c ({signal_1692, signal_1289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1275 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1615, signal_1213}), .a ({signal_1547, signal_1145}), .clk ( clk ), .r ( Fresh[348] ), .c ({signal_1693, signal_1290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1276 ( .s ({SI_s1[3], SI_s0[3]}), .b ({signal_1566, signal_1164}), .a ({signal_1516, signal_1114}), .clk ( clk ), .r ( Fresh[349] ), .c ({signal_1694, signal_1291}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1277 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1637, signal_1234}), .a ({signal_1664, signal_1261}), .clk ( clk ), .r ( Fresh[350] ), .c ({signal_1696, signal_1292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1278 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1636, signal_1233}), .a ({signal_1638, signal_1235}), .clk ( clk ), .r ( Fresh[351] ), .c ({signal_1697, signal_1293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1279 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1645, signal_1242}), .a ({signal_1662, signal_1259}), .clk ( clk ), .r ( Fresh[352] ), .c ({signal_1698, signal_1294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1280 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1681, signal_1278}), .a ({signal_1652, signal_1249}), .clk ( clk ), .r ( Fresh[353] ), .c ({signal_1699, signal_1295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1281 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1676, signal_1273}), .a ({signal_1689, signal_1286}), .clk ( clk ), .r ( Fresh[354] ), .c ({signal_1700, signal_1296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1282 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1632, signal_1229}), .a ({signal_1684, signal_1281}), .clk ( clk ), .r ( Fresh[355] ), .c ({signal_1701, signal_1297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1283 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1675, signal_1272}), .a ({signal_1673, signal_1270}), .clk ( clk ), .r ( Fresh[356] ), .c ({signal_1702, signal_1298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1284 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1672, signal_1269}), .a ({signal_1639, signal_1236}), .clk ( clk ), .r ( Fresh[357] ), .c ({signal_1703, signal_1299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1285 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1690, signal_1287}), .a ({signal_1671, signal_1268}), .clk ( clk ), .r ( Fresh[358] ), .c ({signal_1704, signal_1300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1286 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1649, signal_1246}), .a ({signal_1668, signal_1265}), .clk ( clk ), .r ( Fresh[359] ), .c ({signal_1705, signal_1301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1287 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1647, signal_1244}), .a ({signal_1692, signal_1289}), .clk ( clk ), .r ( Fresh[360] ), .c ({signal_1706, signal_1302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1288 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1674, signal_1271}), .a ({signal_1642, signal_1239}), .clk ( clk ), .r ( Fresh[361] ), .c ({signal_1707, signal_1303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1289 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1667, signal_1264}), .a ({signal_1641, signal_1238}), .clk ( clk ), .r ( Fresh[362] ), .c ({signal_1708, signal_1304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1290 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1669, signal_1266}), .a ({signal_1635, signal_1232}), .clk ( clk ), .r ( Fresh[363] ), .c ({signal_1709, signal_1305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1291 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1666, signal_1263}), .a ({signal_1651, signal_1248}), .clk ( clk ), .r ( Fresh[364] ), .c ({signal_1710, signal_1306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1292 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1663, signal_1260}), .a ({signal_1660, signal_1257}), .clk ( clk ), .r ( Fresh[365] ), .c ({signal_1711, signal_1307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1293 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1655, signal_1252}), .a ({signal_1693, signal_1290}), .clk ( clk ), .r ( Fresh[366] ), .c ({signal_1712, signal_1308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1294 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1683, signal_1280}), .a ({signal_1634, signal_1231}), .clk ( clk ), .r ( Fresh[367] ), .c ({signal_1713, signal_1309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1295 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1682, signal_1279}), .a ({signal_1686, signal_1283}), .clk ( clk ), .r ( Fresh[368] ), .c ({signal_1714, signal_1310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1296 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1640, signal_1237}), .a ({signal_1685, signal_1282}), .clk ( clk ), .r ( Fresh[369] ), .c ({signal_1715, signal_1311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1297 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1680, signal_1277}), .a ({signal_1659, signal_1256}), .clk ( clk ), .r ( Fresh[370] ), .c ({signal_1716, signal_1312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1298 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1661, signal_1258}), .a ({signal_1665, signal_1262}), .clk ( clk ), .r ( Fresh[371] ), .c ({signal_1717, signal_1313}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1299 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1654, signal_1251}), .a ({signal_1658, signal_1255}), .clk ( clk ), .r ( Fresh[372] ), .c ({signal_1718, signal_1314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1300 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1646, signal_1243}), .a ({signal_1670, signal_1267}), .clk ( clk ), .r ( Fresh[373] ), .c ({signal_1719, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1301 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1648, signal_1245}), .a ({signal_1657, signal_1254}), .clk ( clk ), .r ( Fresh[374] ), .c ({signal_1720, signal_1316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1302 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1677, signal_1274}), .a ({signal_1653, signal_1250}), .clk ( clk ), .r ( Fresh[375] ), .c ({signal_1721, signal_1317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1303 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1687, signal_1284}), .a ({signal_1694, signal_1291}), .clk ( clk ), .r ( Fresh[376] ), .c ({signal_1722, signal_1318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1304 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1650, signal_1247}), .a ({signal_1643, signal_1240}), .clk ( clk ), .r ( Fresh[377] ), .c ({signal_1723, signal_1319}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1305 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1644, signal_1241}), .a ({signal_1631, signal_1228}), .clk ( clk ), .r ( Fresh[378] ), .c ({signal_1724, signal_1320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1306 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1656, signal_1253}), .a ({signal_1633, signal_1230}), .clk ( clk ), .r ( Fresh[379] ), .c ({signal_1725, signal_1321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1307 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1678, signal_1275}), .a ({signal_1679, signal_1276}), .clk ( clk ), .r ( Fresh[380] ), .c ({signal_1726, signal_1322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1308 ( .s ({SI_s1[0], SI_s0[0]}), .b ({signal_1688, signal_1285}), .a ({signal_1691, signal_1288}), .clk ( clk ), .r ( Fresh[381] ), .c ({signal_1727, signal_1323}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1309 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1698, signal_1294}), .a ({signal_1718, signal_1314}), .clk ( clk ), .r ( Fresh[382] ), .c ({signal_1729, signal_1324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1310 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1727, signal_1323}), .a ({signal_1705, signal_1301}), .clk ( clk ), .r ( Fresh[383] ), .c ({signal_1730, signal_1325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1311 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1722, signal_1318}), .a ({signal_1697, signal_1293}), .clk ( clk ), .r ( Fresh[384] ), .c ({signal_1731, signal_1326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1312 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1703, signal_1299}), .a ({signal_1712, signal_1308}), .clk ( clk ), .r ( Fresh[385] ), .c ({signal_1732, signal_1327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1313 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1700, signal_1296}), .a ({signal_1720, signal_1316}), .clk ( clk ), .r ( Fresh[386] ), .c ({signal_1733, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1314 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1696, signal_1292}), .a ({signal_1714, signal_1310}), .clk ( clk ), .r ( Fresh[387] ), .c ({signal_1734, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1315 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1701, signal_1297}), .a ({signal_1717, signal_1313}), .clk ( clk ), .r ( Fresh[388] ), .c ({signal_1735, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1316 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1721, signal_1317}), .a ({signal_1708, signal_1304}), .clk ( clk ), .r ( Fresh[389] ), .c ({signal_1736, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1317 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1711, signal_1307}), .a ({signal_1713, signal_1309}), .clk ( clk ), .r ( Fresh[390] ), .c ({signal_1737, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1318 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1716, signal_1312}), .a ({signal_1724, signal_1320}), .clk ( clk ), .r ( Fresh[391] ), .c ({signal_1738, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1319 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1704, signal_1300}), .a ({signal_1702, signal_1298}), .clk ( clk ), .r ( Fresh[392] ), .c ({signal_1739, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1320 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1719, signal_1315}), .a ({signal_1706, signal_1302}), .clk ( clk ), .r ( Fresh[393] ), .c ({signal_1740, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1321 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1709, signal_1305}), .a ({signal_1726, signal_1322}), .clk ( clk ), .r ( Fresh[394] ), .c ({signal_1741, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1322 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1707, signal_1303}), .a ({signal_1725, signal_1321}), .clk ( clk ), .r ( Fresh[395] ), .c ({signal_1742, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1323 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1723, signal_1319}), .a ({signal_1710, signal_1306}), .clk ( clk ), .r ( Fresh[396] ), .c ({signal_1743, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1324 ( .s ({SI_s1[7], SI_s0[7]}), .b ({signal_1699, signal_1295}), .a ({signal_1715, signal_1311}), .clk ( clk ), .r ( Fresh[397] ), .c ({signal_1744, signal_1339}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1325 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1730, signal_1325}), .a ({signal_1741, signal_1336}), .clk ( clk ), .r ( Fresh[398] ), .c ({signal_1746, signal_30}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1326 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1732, signal_1327}), .a ({signal_1733, signal_1328}), .clk ( clk ), .r ( Fresh[399] ), .c ({signal_1747, signal_23}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1327 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1743, signal_1338}), .a ({signal_1736, signal_1331}), .clk ( clk ), .r ( Fresh[400] ), .c ({signal_1748, signal_29}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1328 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1731, signal_1326}), .a ({signal_1744, signal_1339}), .clk ( clk ), .r ( Fresh[401] ), .c ({signal_1749, signal_28}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1329 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1740, signal_1335}), .a ({signal_1738, signal_1333}), .clk ( clk ), .r ( Fresh[402] ), .c ({signal_1750, signal_26}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1330 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1742, signal_1337}), .a ({signal_1735, signal_1330}), .clk ( clk ), .r ( Fresh[403] ), .c ({signal_1751, signal_27}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1331 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1739, signal_1334}), .a ({signal_1737, signal_1332}), .clk ( clk ), .r ( Fresh[404] ), .c ({signal_1752, signal_24}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_1332 ( .s ({SI_s1[6], SI_s0[6]}), .b ({signal_1734, signal_1329}), .a ({signal_1729, signal_1324}), .clk ( clk ), .r ( Fresh[405] ), .c ({signal_1753, signal_25}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_0 ( .clk ( signal_2169 ), .D ({signal_1747, signal_23}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1 ( .clk ( signal_2169 ), .D ({signal_1752, signal_24}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_2 ( .clk ( signal_2169 ), .D ({signal_1753, signal_25}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3 ( .clk ( signal_2169 ), .D ({signal_1750, signal_26}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_4 ( .clk ( signal_2169 ), .D ({signal_1751, signal_27}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_5 ( .clk ( signal_2169 ), .D ({signal_1749, signal_28}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_6 ( .clk ( signal_2169 ), .D ({signal_1748, signal_29}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_7 ( .clk ( signal_2169 ), .D ({signal_1746, signal_30}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
