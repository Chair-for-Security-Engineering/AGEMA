/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module LED_HPC2_ClockGating_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1, Synch);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    output Synch ;
    wire n15 ;
    wire n14 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n34 ;
    wire LED_128_Instance_n33 ;
    wire LED_128_Instance_n32 ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n21 ;
    wire LED_128_Instance_n20 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n15 ;
    wire LED_128_Instance_n14 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n10 ;
    wire LED_128_Instance_n2 ;
    wire LED_128_Instance_n1 ;
    wire LED_128_Instance_n27 ;
    wire LED_128_Instance_N9 ;
    wire LED_128_Instance_n28 ;
    wire LED_128_Instance_N8 ;
    wire LED_128_Instance_n30 ;
    wire LED_128_Instance_N7 ;
    wire LED_128_Instance_n5 ;
    wire LED_128_Instance_N6 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_N5 ;
    wire LED_128_Instance_n6 ;
    wire LED_128_Instance_N4 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_N13 ;
    wire LED_128_Instance_n25 ;
    wire LED_128_Instance_N12 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n26 ;
    wire LED_128_Instance_N11 ;
    wire LED_128_Instance_n4 ;
    wire LED_128_Instance_N10 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_addroundkey_out_0_ ;
    wire LED_128_Instance_addroundkey_out_1_ ;
    wire LED_128_Instance_addroundkey_out_2_ ;
    wire LED_128_Instance_addroundkey_out_3_ ;
    wire LED_128_Instance_addroundkey_out_4_ ;
    wire LED_128_Instance_addroundkey_out_5_ ;
    wire LED_128_Instance_addroundkey_out_6_ ;
    wire LED_128_Instance_addroundkey_out_16_ ;
    wire LED_128_Instance_addroundkey_out_17_ ;
    wire LED_128_Instance_addroundkey_out_18_ ;
    wire LED_128_Instance_addroundkey_out_19_ ;
    wire LED_128_Instance_addroundkey_out_20_ ;
    wire LED_128_Instance_addroundkey_out_21_ ;
    wire LED_128_Instance_addroundkey_out_22_ ;
    wire LED_128_Instance_addroundkey_out_32_ ;
    wire LED_128_Instance_addroundkey_out_33_ ;
    wire LED_128_Instance_addroundkey_out_34_ ;
    wire LED_128_Instance_addroundkey_out_35_ ;
    wire LED_128_Instance_addroundkey_out_36_ ;
    wire LED_128_Instance_addroundkey_out_37_ ;
    wire LED_128_Instance_addroundkey_out_38_ ;
    wire LED_128_Instance_addroundkey_out_48_ ;
    wire LED_128_Instance_addroundkey_out_49_ ;
    wire LED_128_Instance_addroundkey_out_50_ ;
    wire LED_128_Instance_addroundkey_out_51_ ;
    wire LED_128_Instance_addroundkey_out_52_ ;
    wire LED_128_Instance_addroundkey_out_53_ ;
    wire LED_128_Instance_addroundkey_out_54_ ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_n11 ;
    wire LED_128_Instance_MUX_state0_n10 ;
    wire LED_128_Instance_MUX_state0_n9 ;
    wire LED_128_Instance_MUX_state0_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n10 ;
    wire LED_128_Instance_MUX_current_roundkey_n9 ;
    wire LED_128_Instance_MUX_current_roundkey_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n7 ;
    wire LED_128_Instance_MUX_addroundkey_out_n9 ;
    wire LED_128_Instance_MUX_addroundkey_out_n8 ;
    wire LED_128_Instance_MUX_addroundkey_out_n7 ;
    wire LED_128_Instance_SBox_Instance_0_n3 ;
    wire LED_128_Instance_SBox_Instance_0_n2 ;
    wire LED_128_Instance_SBox_Instance_0_n1 ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_n3 ;
    wire LED_128_Instance_SBox_Instance_1_n2 ;
    wire LED_128_Instance_SBox_Instance_1_n1 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_n3 ;
    wire LED_128_Instance_SBox_Instance_2_n2 ;
    wire LED_128_Instance_SBox_Instance_2_n1 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_n3 ;
    wire LED_128_Instance_SBox_Instance_3_n2 ;
    wire LED_128_Instance_SBox_Instance_3_n1 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_n3 ;
    wire LED_128_Instance_SBox_Instance_4_n2 ;
    wire LED_128_Instance_SBox_Instance_4_n1 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_n3 ;
    wire LED_128_Instance_SBox_Instance_5_n2 ;
    wire LED_128_Instance_SBox_Instance_5_n1 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_n3 ;
    wire LED_128_Instance_SBox_Instance_6_n2 ;
    wire LED_128_Instance_SBox_Instance_6_n1 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_n3 ;
    wire LED_128_Instance_SBox_Instance_7_n2 ;
    wire LED_128_Instance_SBox_Instance_7_n1 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_n3 ;
    wire LED_128_Instance_SBox_Instance_8_n2 ;
    wire LED_128_Instance_SBox_Instance_8_n1 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_n3 ;
    wire LED_128_Instance_SBox_Instance_9_n2 ;
    wire LED_128_Instance_SBox_Instance_9_n1 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_n3 ;
    wire LED_128_Instance_SBox_Instance_10_n2 ;
    wire LED_128_Instance_SBox_Instance_10_n1 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_n3 ;
    wire LED_128_Instance_SBox_Instance_11_n2 ;
    wire LED_128_Instance_SBox_Instance_11_n1 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_n3 ;
    wire LED_128_Instance_SBox_Instance_12_n2 ;
    wire LED_128_Instance_SBox_Instance_12_n1 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_n3 ;
    wire LED_128_Instance_SBox_Instance_13_n2 ;
    wire LED_128_Instance_SBox_Instance_13_n1 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_n3 ;
    wire LED_128_Instance_SBox_Instance_14_n2 ;
    wire LED_128_Instance_SBox_Instance_14_n1 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_n3 ;
    wire LED_128_Instance_SBox_Instance_15_n2 ;
    wire LED_128_Instance_SBox_Instance_15_n1 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_0__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state1 ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2515 ;
    wire clk_gated ;

    /* cells in depth 0 */
    NOR2_X1 U16 ( .A1 (roundconstant[4]), .A2 (roundconstant[1]), .ZN (n14) ) ;
    NAND2_X1 U17 ( .A1 (roundconstant[0]), .A2 (n14), .ZN (n16) ) ;
    NOR2_X1 U18 ( .A1 (roundconstant[5]), .A2 (n16), .ZN (n17) ) ;
    NAND2_X1 U19 ( .A1 (roundconstant[3]), .A2 (n17), .ZN (n18) ) ;
    NOR2_X1 U20 ( .A1 (roundconstant[2]), .A2 (n18), .ZN (n19) ) ;
    NOR2_X1 U21 ( .A1 (OUT_done), .A2 (n19), .ZN (n20) ) ;
    NOR2_X1 U22 ( .A1 (IN_reset), .A2 (n20), .ZN (n15) ) ;
    NAND2_X1 LED_128_Instance_U30 ( .A1 (LED_128_Instance_n33), .A2 (LED_128_Instance_n32), .ZN (LED_128_Instance_n34) ) ;
    XNOR2_X1 LED_128_Instance_U29 ( .A (LED_128_Instance_n25), .B (LED_128_Instance_n23), .ZN (LED_128_Instance_n32) ) ;
    XOR2_X1 LED_128_Instance_U28 ( .A (LED_128_Instance_n4), .B (LED_128_Instance_n26), .Z (LED_128_Instance_n23) ) ;
    NAND2_X1 LED_128_Instance_U27 ( .A1 (LED_128_Instance_n21), .A2 (LED_128_Instance_n20), .ZN (LED_128_Instance_n33) ) ;
    NAND2_X1 LED_128_Instance_U26 ( .A1 (LED_128_Instance_n19), .A2 (LED_128_Instance_n18), .ZN (LED_128_Instance_n20) ) ;
    NOR2_X1 LED_128_Instance_U25 ( .A1 (LED_128_Instance_n24), .A2 (LED_128_Instance_n1), .ZN (LED_128_Instance_n18) ) ;
    NOR2_X1 LED_128_Instance_U24 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n19) ) ;
    NAND2_X1 LED_128_Instance_U23 ( .A1 (LED_128_Instance_n1), .A2 (LED_128_Instance_n17), .ZN (LED_128_Instance_n21) ) ;
    AND2_X1 LED_128_Instance_U22 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n17) ) ;
    NAND2_X1 LED_128_Instance_U21 ( .A1 (LED_128_Instance_n29), .A2 (LED_128_Instance_n14), .ZN (LED_128_Instance_n15) ) ;
    NOR2_X1 LED_128_Instance_U20 ( .A1 (LED_128_Instance_n6), .A2 (LED_128_Instance_n13), .ZN (LED_128_Instance_n14) ) ;
    NAND2_X1 LED_128_Instance_U19 ( .A1 (LED_128_Instance_n5), .A2 (roundconstant[3]), .ZN (LED_128_Instance_n13) ) ;
    NAND2_X1 LED_128_Instance_U18 ( .A1 (LED_128_Instance_n28), .A2 (LED_128_Instance_n27), .ZN (LED_128_Instance_n16) ) ;
    NOR2_X1 LED_128_Instance_U17 ( .A1 (LED_128_Instance_n28), .A2 (IN_reset), .ZN (LED_128_Instance_N9) ) ;
    NOR2_X1 LED_128_Instance_U16 ( .A1 (IN_reset), .A2 (LED_128_Instance_n30), .ZN (LED_128_Instance_N8) ) ;
    NOR2_X1 LED_128_Instance_U15 ( .A1 (IN_reset), .A2 (LED_128_Instance_n5), .ZN (LED_128_Instance_N7) ) ;
    NOR2_X1 LED_128_Instance_U14 ( .A1 (IN_reset), .A2 (LED_128_Instance_n29), .ZN (LED_128_Instance_N6) ) ;
    NOR2_X1 LED_128_Instance_U13 ( .A1 (IN_reset), .A2 (LED_128_Instance_n6), .ZN (LED_128_Instance_N5) ) ;
    NOR2_X1 LED_128_Instance_U12 ( .A1 (LED_128_Instance_n1), .A2 (IN_reset), .ZN (LED_128_Instance_N13) ) ;
    NOR2_X1 LED_128_Instance_U11 ( .A1 (LED_128_Instance_n8), .A2 (IN_reset), .ZN (LED_128_Instance_N12) ) ;
    NOR2_X1 LED_128_Instance_U10 ( .A1 (LED_128_Instance_n4), .A2 (IN_reset), .ZN (LED_128_Instance_N11) ) ;
    NOR2_X1 LED_128_Instance_U9 ( .A1 (LED_128_Instance_n2), .A2 (IN_reset), .ZN (LED_128_Instance_N10) ) ;
    OR2_X1 LED_128_Instance_U8 ( .A1 (LED_128_Instance_n2), .A2 (LED_128_Instance_n21), .ZN (LED_128_Instance_n11) ) ;
    NAND2_X1 LED_128_Instance_U7 ( .A1 (LED_128_Instance_n34), .A2 (LED_128_Instance_n11), .ZN (LED_128_Instance_n31) ) ;
    NOR2_X1 LED_128_Instance_U6 ( .A1 (LED_128_Instance_n16), .A2 (LED_128_Instance_n15), .ZN (LED_128_Instance_n22) ) ;
    INV_X1 LED_128_Instance_U5 ( .A (LED_128_Instance_n11), .ZN (LED_128_Instance_n12) ) ;
    OR2_X1 LED_128_Instance_U4 ( .A1 (IN_reset), .A2 (LED_128_Instance_n10), .ZN (LED_128_Instance_N4) ) ;
    XNOR2_X1 LED_128_Instance_U3 ( .A (LED_128_Instance_n28), .B (LED_128_Instance_n27), .ZN (LED_128_Instance_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U4 ( .A (LED_128_Instance_n22), .ZN (LED_128_Instance_MUX_state0_n11) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U3 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n8) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U2 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U1 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U4 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U3 ( .A (LED_128_Instance_n12), .ZN (LED_128_Instance_MUX_current_roundkey_n10) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U2 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n7) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U1 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({new_AGEMA_signal_1330, LED_128_Instance_current_roundkey[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({new_AGEMA_signal_1395, LED_128_Instance_current_roundkey[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({new_AGEMA_signal_1333, LED_128_Instance_current_roundkey[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({new_AGEMA_signal_1401, LED_128_Instance_current_roundkey[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({new_AGEMA_signal_1407, LED_128_Instance_current_roundkey[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({new_AGEMA_signal_1413, LED_128_Instance_current_roundkey[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({new_AGEMA_signal_1416, LED_128_Instance_current_roundkey[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({new_AGEMA_signal_1419, LED_128_Instance_current_roundkey[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({new_AGEMA_signal_1422, LED_128_Instance_current_roundkey[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({new_AGEMA_signal_1425, LED_128_Instance_current_roundkey[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({new_AGEMA_signal_1428, LED_128_Instance_current_roundkey[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({new_AGEMA_signal_1431, LED_128_Instance_current_roundkey[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({new_AGEMA_signal_1434, LED_128_Instance_current_roundkey[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({new_AGEMA_signal_1336, LED_128_Instance_current_roundkey[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({new_AGEMA_signal_1437, LED_128_Instance_current_roundkey[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({new_AGEMA_signal_1440, LED_128_Instance_current_roundkey[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({new_AGEMA_signal_1339, LED_128_Instance_current_roundkey[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({new_AGEMA_signal_1443, LED_128_Instance_current_roundkey[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({new_AGEMA_signal_1446, LED_128_Instance_current_roundkey[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({new_AGEMA_signal_1342, LED_128_Instance_current_roundkey[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({new_AGEMA_signal_1449, LED_128_Instance_current_roundkey[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({new_AGEMA_signal_1345, LED_128_Instance_current_roundkey[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({new_AGEMA_signal_1452, LED_128_Instance_current_roundkey[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({new_AGEMA_signal_1348, LED_128_Instance_current_roundkey[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({new_AGEMA_signal_1455, LED_128_Instance_current_roundkey[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({new_AGEMA_signal_1351, LED_128_Instance_current_roundkey[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({new_AGEMA_signal_1458, LED_128_Instance_current_roundkey[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({new_AGEMA_signal_1461, LED_128_Instance_current_roundkey[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({new_AGEMA_signal_1464, LED_128_Instance_current_roundkey[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({new_AGEMA_signal_1354, LED_128_Instance_current_roundkey[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({new_AGEMA_signal_1467, LED_128_Instance_current_roundkey[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({new_AGEMA_signal_1357, LED_128_Instance_current_roundkey[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({new_AGEMA_signal_1360, LED_128_Instance_current_roundkey[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({new_AGEMA_signal_1363, LED_128_Instance_current_roundkey[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({new_AGEMA_signal_1473, LED_128_Instance_current_roundkey[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({new_AGEMA_signal_1366, LED_128_Instance_current_roundkey[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({new_AGEMA_signal_1479, LED_128_Instance_current_roundkey[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({new_AGEMA_signal_1485, LED_128_Instance_current_roundkey[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({new_AGEMA_signal_1491, LED_128_Instance_current_roundkey[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({new_AGEMA_signal_1497, LED_128_Instance_current_roundkey[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({new_AGEMA_signal_1503, LED_128_Instance_current_roundkey[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({new_AGEMA_signal_1509, LED_128_Instance_current_roundkey[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({new_AGEMA_signal_1515, LED_128_Instance_current_roundkey[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({new_AGEMA_signal_1521, LED_128_Instance_current_roundkey[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({new_AGEMA_signal_1527, LED_128_Instance_current_roundkey[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({new_AGEMA_signal_1533, LED_128_Instance_current_roundkey[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({new_AGEMA_signal_1539, LED_128_Instance_current_roundkey[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({new_AGEMA_signal_1545, LED_128_Instance_current_roundkey[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U64 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({new_AGEMA_signal_1416, LED_128_Instance_current_roundkey[9]}), .c ({new_AGEMA_signal_1554, LED_128_Instance_addroundkey_tmp[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U63 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({new_AGEMA_signal_1413, LED_128_Instance_current_roundkey[8]}), .c ({new_AGEMA_signal_1556, LED_128_Instance_addroundkey_tmp[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U62 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[7]}), .c ({new_AGEMA_signal_1558, LED_128_Instance_addroundkey_tmp[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U61 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({new_AGEMA_signal_1407, LED_128_Instance_current_roundkey[6]}), .c ({new_AGEMA_signal_1560, LED_128_Instance_addroundkey_tmp[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U60 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({new_AGEMA_signal_1545, LED_128_Instance_current_roundkey[63]}), .c ({new_AGEMA_signal_1562, LED_128_Instance_addroundkey_tmp[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U59 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[62]}), .c ({new_AGEMA_signal_1564, LED_128_Instance_addroundkey_tmp[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U58 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({new_AGEMA_signal_1539, LED_128_Instance_current_roundkey[61]}), .c ({new_AGEMA_signal_1566, LED_128_Instance_addroundkey_tmp[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U57 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[60]}), .c ({new_AGEMA_signal_1568, LED_128_Instance_addroundkey_tmp[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U56 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[5]}), .c ({new_AGEMA_signal_1570, LED_128_Instance_addroundkey_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U55 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({new_AGEMA_signal_1533, LED_128_Instance_current_roundkey[59]}), .c ({new_AGEMA_signal_1572, LED_128_Instance_addroundkey_tmp[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U54 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[58]}), .c ({new_AGEMA_signal_1574, LED_128_Instance_addroundkey_tmp[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U53 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({new_AGEMA_signal_1527, LED_128_Instance_current_roundkey[57]}), .c ({new_AGEMA_signal_1576, LED_128_Instance_addroundkey_tmp[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U52 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[56]}), .c ({new_AGEMA_signal_1578, LED_128_Instance_addroundkey_tmp[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U51 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({new_AGEMA_signal_1521, LED_128_Instance_current_roundkey[55]}), .c ({new_AGEMA_signal_1580, LED_128_Instance_addroundkey_tmp[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U50 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[54]}), .c ({new_AGEMA_signal_1582, LED_128_Instance_addroundkey_tmp[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U49 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({new_AGEMA_signal_1515, LED_128_Instance_current_roundkey[53]}), .c ({new_AGEMA_signal_1584, LED_128_Instance_addroundkey_tmp[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U48 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[52]}), .c ({new_AGEMA_signal_1586, LED_128_Instance_addroundkey_tmp[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U47 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({new_AGEMA_signal_1509, LED_128_Instance_current_roundkey[51]}), .c ({new_AGEMA_signal_1588, LED_128_Instance_addroundkey_tmp[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U46 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[50]}), .c ({new_AGEMA_signal_1590, LED_128_Instance_addroundkey_tmp[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U45 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({new_AGEMA_signal_1401, LED_128_Instance_current_roundkey[4]}), .c ({new_AGEMA_signal_1592, LED_128_Instance_addroundkey_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U44 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({new_AGEMA_signal_1503, LED_128_Instance_current_roundkey[49]}), .c ({new_AGEMA_signal_1594, LED_128_Instance_addroundkey_tmp[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U43 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[48]}), .c ({new_AGEMA_signal_1596, LED_128_Instance_addroundkey_tmp[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U42 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({new_AGEMA_signal_1497, LED_128_Instance_current_roundkey[47]}), .c ({new_AGEMA_signal_1598, LED_128_Instance_addroundkey_tmp[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U41 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[46]}), .c ({new_AGEMA_signal_1600, LED_128_Instance_addroundkey_tmp[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U40 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({new_AGEMA_signal_1491, LED_128_Instance_current_roundkey[45]}), .c ({new_AGEMA_signal_1602, LED_128_Instance_addroundkey_tmp[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U39 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[44]}), .c ({new_AGEMA_signal_1604, LED_128_Instance_addroundkey_tmp[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U38 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({new_AGEMA_signal_1485, LED_128_Instance_current_roundkey[43]}), .c ({new_AGEMA_signal_1606, LED_128_Instance_addroundkey_tmp[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U37 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[42]}), .c ({new_AGEMA_signal_1608, LED_128_Instance_addroundkey_tmp[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U36 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({new_AGEMA_signal_1479, LED_128_Instance_current_roundkey[41]}), .c ({new_AGEMA_signal_1610, LED_128_Instance_addroundkey_tmp[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U35 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[40]}), .c ({new_AGEMA_signal_1612, LED_128_Instance_addroundkey_tmp[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U34 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({new_AGEMA_signal_1333, LED_128_Instance_current_roundkey[3]}), .c ({new_AGEMA_signal_1368, LED_128_Instance_addroundkey_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U33 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({new_AGEMA_signal_1366, LED_128_Instance_current_roundkey[39]}), .c ({new_AGEMA_signal_1370, LED_128_Instance_addroundkey_tmp[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U32 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({new_AGEMA_signal_1473, LED_128_Instance_current_roundkey[38]}), .c ({new_AGEMA_signal_1614, LED_128_Instance_addroundkey_tmp[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U31 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[37]}), .c ({new_AGEMA_signal_1616, LED_128_Instance_addroundkey_tmp[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U30 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({new_AGEMA_signal_1363, LED_128_Instance_current_roundkey[36]}), .c ({new_AGEMA_signal_1372, LED_128_Instance_addroundkey_tmp[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U29 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({new_AGEMA_signal_1360, LED_128_Instance_current_roundkey[35]}), .c ({new_AGEMA_signal_1374, LED_128_Instance_addroundkey_tmp[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U28 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({new_AGEMA_signal_1357, LED_128_Instance_current_roundkey[34]}), .c ({new_AGEMA_signal_1376, LED_128_Instance_addroundkey_tmp[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U27 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({new_AGEMA_signal_1467, LED_128_Instance_current_roundkey[33]}), .c ({new_AGEMA_signal_1618, LED_128_Instance_addroundkey_tmp[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U26 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({new_AGEMA_signal_1354, LED_128_Instance_current_roundkey[32]}), .c ({new_AGEMA_signal_1378, LED_128_Instance_addroundkey_tmp[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U25 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({new_AGEMA_signal_1464, LED_128_Instance_current_roundkey[31]}), .c ({new_AGEMA_signal_1620, LED_128_Instance_addroundkey_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U24 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({new_AGEMA_signal_1461, LED_128_Instance_current_roundkey[30]}), .c ({new_AGEMA_signal_1622, LED_128_Instance_addroundkey_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U23 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[2]}), .c ({new_AGEMA_signal_1624, LED_128_Instance_addroundkey_tmp[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U22 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({new_AGEMA_signal_1458, LED_128_Instance_current_roundkey[29]}), .c ({new_AGEMA_signal_1626, LED_128_Instance_addroundkey_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U21 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({new_AGEMA_signal_1351, LED_128_Instance_current_roundkey[28]}), .c ({new_AGEMA_signal_1380, LED_128_Instance_addroundkey_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U20 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({new_AGEMA_signal_1455, LED_128_Instance_current_roundkey[27]}), .c ({new_AGEMA_signal_1628, LED_128_Instance_addroundkey_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U19 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({new_AGEMA_signal_1348, LED_128_Instance_current_roundkey[26]}), .c ({new_AGEMA_signal_1382, LED_128_Instance_addroundkey_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U18 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({new_AGEMA_signal_1452, LED_128_Instance_current_roundkey[25]}), .c ({new_AGEMA_signal_1630, LED_128_Instance_addroundkey_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U17 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({new_AGEMA_signal_1345, LED_128_Instance_current_roundkey[24]}), .c ({new_AGEMA_signal_1384, LED_128_Instance_addroundkey_tmp[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U16 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({new_AGEMA_signal_1449, LED_128_Instance_current_roundkey[23]}), .c ({new_AGEMA_signal_1632, LED_128_Instance_addroundkey_tmp[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U15 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({new_AGEMA_signal_1342, LED_128_Instance_current_roundkey[22]}), .c ({new_AGEMA_signal_1386, LED_128_Instance_addroundkey_tmp[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U14 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({new_AGEMA_signal_1446, LED_128_Instance_current_roundkey[21]}), .c ({new_AGEMA_signal_1634, LED_128_Instance_addroundkey_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U13 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({new_AGEMA_signal_1443, LED_128_Instance_current_roundkey[20]}), .c ({new_AGEMA_signal_1636, LED_128_Instance_addroundkey_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U12 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({new_AGEMA_signal_1395, LED_128_Instance_current_roundkey[1]}), .c ({new_AGEMA_signal_1638, LED_128_Instance_addroundkey_tmp[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U11 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({new_AGEMA_signal_1339, LED_128_Instance_current_roundkey[19]}), .c ({new_AGEMA_signal_1388, LED_128_Instance_addroundkey_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U10 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({new_AGEMA_signal_1440, LED_128_Instance_current_roundkey[18]}), .c ({new_AGEMA_signal_1640, LED_128_Instance_addroundkey_tmp[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U9 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({new_AGEMA_signal_1437, LED_128_Instance_current_roundkey[17]}), .c ({new_AGEMA_signal_1642, LED_128_Instance_addroundkey_tmp[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U8 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({new_AGEMA_signal_1336, LED_128_Instance_current_roundkey[16]}), .c ({new_AGEMA_signal_1390, LED_128_Instance_addroundkey_tmp[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U7 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({new_AGEMA_signal_1434, LED_128_Instance_current_roundkey[15]}), .c ({new_AGEMA_signal_1644, LED_128_Instance_addroundkey_tmp[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U6 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({new_AGEMA_signal_1431, LED_128_Instance_current_roundkey[14]}), .c ({new_AGEMA_signal_1646, LED_128_Instance_addroundkey_tmp[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U5 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({new_AGEMA_signal_1428, LED_128_Instance_current_roundkey[13]}), .c ({new_AGEMA_signal_1648, LED_128_Instance_addroundkey_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U4 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({new_AGEMA_signal_1425, LED_128_Instance_current_roundkey[12]}), .c ({new_AGEMA_signal_1650, LED_128_Instance_addroundkey_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U3 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({new_AGEMA_signal_1422, LED_128_Instance_current_roundkey[11]}), .c ({new_AGEMA_signal_1652, LED_128_Instance_addroundkey_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U2 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({new_AGEMA_signal_1419, LED_128_Instance_current_roundkey[10]}), .c ({new_AGEMA_signal_1654, LED_128_Instance_addroundkey_tmp[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_addRoundKey_instance_U1 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({new_AGEMA_signal_1330, LED_128_Instance_current_roundkey[0]}), .c ({new_AGEMA_signal_1392, LED_128_Instance_addroundkey_tmp[0]}) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U3 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n7) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U2 ( .A (LED_128_Instance_n31), .ZN (LED_128_Instance_MUX_addroundkey_out_n9) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U1 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({new_AGEMA_signal_1392, LED_128_Instance_addroundkey_tmp[0]}), .c ({new_AGEMA_signal_1546, LED_128_Instance_addroundkey_out_0_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({new_AGEMA_signal_1638, LED_128_Instance_addroundkey_tmp[1]}), .c ({new_AGEMA_signal_1666, LED_128_Instance_addroundkey_out_1_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({new_AGEMA_signal_1624, LED_128_Instance_addroundkey_tmp[2]}), .c ({new_AGEMA_signal_1667, LED_128_Instance_addroundkey_out_2_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({new_AGEMA_signal_1368, LED_128_Instance_addroundkey_tmp[3]}), .c ({new_AGEMA_signal_1547, LED_128_Instance_addroundkey_out_3_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({new_AGEMA_signal_1592, LED_128_Instance_addroundkey_tmp[4]}), .c ({new_AGEMA_signal_1668, LED_128_Instance_addroundkey_out_4_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({new_AGEMA_signal_1570, LED_128_Instance_addroundkey_tmp[5]}), .c ({new_AGEMA_signal_1669, LED_128_Instance_addroundkey_out_5_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({new_AGEMA_signal_1560, LED_128_Instance_addroundkey_tmp[6]}), .c ({new_AGEMA_signal_1670, LED_128_Instance_addroundkey_out_6_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({new_AGEMA_signal_1558, LED_128_Instance_addroundkey_tmp[7]}), .c ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({new_AGEMA_signal_1556, LED_128_Instance_addroundkey_tmp[8]}), .c ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({new_AGEMA_signal_1554, LED_128_Instance_addroundkey_tmp[9]}), .c ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({new_AGEMA_signal_1654, LED_128_Instance_addroundkey_tmp[10]}), .c ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({new_AGEMA_signal_1652, LED_128_Instance_addroundkey_tmp[11]}), .c ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({new_AGEMA_signal_1650, LED_128_Instance_addroundkey_tmp[12]}), .c ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({new_AGEMA_signal_1648, LED_128_Instance_addroundkey_tmp[13]}), .c ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({new_AGEMA_signal_1646, LED_128_Instance_addroundkey_tmp[14]}), .c ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({new_AGEMA_signal_1644, LED_128_Instance_addroundkey_tmp[15]}), .c ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({new_AGEMA_signal_1390, LED_128_Instance_addroundkey_tmp[16]}), .c ({new_AGEMA_signal_1548, LED_128_Instance_addroundkey_out_16_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({new_AGEMA_signal_1642, LED_128_Instance_addroundkey_tmp[17]}), .c ({new_AGEMA_signal_1680, LED_128_Instance_addroundkey_out_17_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({new_AGEMA_signal_1640, LED_128_Instance_addroundkey_tmp[18]}), .c ({new_AGEMA_signal_1681, LED_128_Instance_addroundkey_out_18_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({new_AGEMA_signal_1388, LED_128_Instance_addroundkey_tmp[19]}), .c ({new_AGEMA_signal_1549, LED_128_Instance_addroundkey_out_19_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({new_AGEMA_signal_1636, LED_128_Instance_addroundkey_tmp[20]}), .c ({new_AGEMA_signal_1682, LED_128_Instance_addroundkey_out_20_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({new_AGEMA_signal_1634, LED_128_Instance_addroundkey_tmp[21]}), .c ({new_AGEMA_signal_1683, LED_128_Instance_addroundkey_out_21_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({new_AGEMA_signal_1386, LED_128_Instance_addroundkey_tmp[22]}), .c ({new_AGEMA_signal_1550, LED_128_Instance_addroundkey_out_22_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({new_AGEMA_signal_1632, LED_128_Instance_addroundkey_tmp[23]}), .c ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({new_AGEMA_signal_1384, LED_128_Instance_addroundkey_tmp[24]}), .c ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({new_AGEMA_signal_1630, LED_128_Instance_addroundkey_tmp[25]}), .c ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({new_AGEMA_signal_1382, LED_128_Instance_addroundkey_tmp[26]}), .c ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({new_AGEMA_signal_1628, LED_128_Instance_addroundkey_tmp[27]}), .c ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({new_AGEMA_signal_1380, LED_128_Instance_addroundkey_tmp[28]}), .c ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({new_AGEMA_signal_1626, LED_128_Instance_addroundkey_tmp[29]}), .c ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({new_AGEMA_signal_1622, LED_128_Instance_addroundkey_tmp[30]}), .c ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({new_AGEMA_signal_1620, LED_128_Instance_addroundkey_tmp[31]}), .c ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({new_AGEMA_signal_1378, LED_128_Instance_addroundkey_tmp[32]}), .c ({new_AGEMA_signal_1656, LED_128_Instance_addroundkey_out_32_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({new_AGEMA_signal_1618, LED_128_Instance_addroundkey_tmp[33]}), .c ({new_AGEMA_signal_1690, LED_128_Instance_addroundkey_out_33_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({new_AGEMA_signal_1376, LED_128_Instance_addroundkey_tmp[34]}), .c ({new_AGEMA_signal_1657, LED_128_Instance_addroundkey_out_34_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({new_AGEMA_signal_1374, LED_128_Instance_addroundkey_tmp[35]}), .c ({new_AGEMA_signal_1658, LED_128_Instance_addroundkey_out_35_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({new_AGEMA_signal_1372, LED_128_Instance_addroundkey_tmp[36]}), .c ({new_AGEMA_signal_1659, LED_128_Instance_addroundkey_out_36_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({new_AGEMA_signal_1616, LED_128_Instance_addroundkey_tmp[37]}), .c ({new_AGEMA_signal_1691, LED_128_Instance_addroundkey_out_37_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({new_AGEMA_signal_1614, LED_128_Instance_addroundkey_tmp[38]}), .c ({new_AGEMA_signal_1692, LED_128_Instance_addroundkey_out_38_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({new_AGEMA_signal_1370, LED_128_Instance_addroundkey_tmp[39]}), .c ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({new_AGEMA_signal_1612, LED_128_Instance_addroundkey_tmp[40]}), .c ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({new_AGEMA_signal_1610, LED_128_Instance_addroundkey_tmp[41]}), .c ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({new_AGEMA_signal_1608, LED_128_Instance_addroundkey_tmp[42]}), .c ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({new_AGEMA_signal_1606, LED_128_Instance_addroundkey_tmp[43]}), .c ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({new_AGEMA_signal_1604, LED_128_Instance_addroundkey_tmp[44]}), .c ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({new_AGEMA_signal_1602, LED_128_Instance_addroundkey_tmp[45]}), .c ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({new_AGEMA_signal_1600, LED_128_Instance_addroundkey_tmp[46]}), .c ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({new_AGEMA_signal_1598, LED_128_Instance_addroundkey_tmp[47]}), .c ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({new_AGEMA_signal_1596, LED_128_Instance_addroundkey_tmp[48]}), .c ({new_AGEMA_signal_1701, LED_128_Instance_addroundkey_out_48_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({new_AGEMA_signal_1594, LED_128_Instance_addroundkey_tmp[49]}), .c ({new_AGEMA_signal_1702, LED_128_Instance_addroundkey_out_49_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({new_AGEMA_signal_1590, LED_128_Instance_addroundkey_tmp[50]}), .c ({new_AGEMA_signal_1703, LED_128_Instance_addroundkey_out_50_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({new_AGEMA_signal_1588, LED_128_Instance_addroundkey_tmp[51]}), .c ({new_AGEMA_signal_1704, LED_128_Instance_addroundkey_out_51_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({new_AGEMA_signal_1586, LED_128_Instance_addroundkey_tmp[52]}), .c ({new_AGEMA_signal_1705, LED_128_Instance_addroundkey_out_52_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({new_AGEMA_signal_1584, LED_128_Instance_addroundkey_tmp[53]}), .c ({new_AGEMA_signal_1706, LED_128_Instance_addroundkey_out_53_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({new_AGEMA_signal_1582, LED_128_Instance_addroundkey_tmp[54]}), .c ({new_AGEMA_signal_1707, LED_128_Instance_addroundkey_out_54_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({new_AGEMA_signal_1580, LED_128_Instance_addroundkey_tmp[55]}), .c ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({new_AGEMA_signal_1578, LED_128_Instance_addroundkey_tmp[56]}), .c ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({new_AGEMA_signal_1576, LED_128_Instance_addroundkey_tmp[57]}), .c ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({new_AGEMA_signal_1574, LED_128_Instance_addroundkey_tmp[58]}), .c ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({new_AGEMA_signal_1572, LED_128_Instance_addroundkey_tmp[59]}), .c ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({new_AGEMA_signal_1568, LED_128_Instance_addroundkey_tmp[60]}), .c ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({new_AGEMA_signal_1566, LED_128_Instance_addroundkey_tmp[61]}), .c ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({new_AGEMA_signal_1564, LED_128_Instance_addroundkey_tmp[62]}), .c ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({new_AGEMA_signal_1562, LED_128_Instance_addroundkey_tmp[63]}), .c ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U28 ( .a ({1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_1670, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U27 ( .a ({1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_1669, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U26 ( .a ({1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1707, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U25 ( .a ({1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_1706, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U24 ( .a ({1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_1705, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U23 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1704, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U22 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1703, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U21 ( .a ({1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_1668, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U20 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1702, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U19 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1701, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U18 ( .a ({1'b0, 1'b1}), .b ({new_AGEMA_signal_1547, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U17 ( .a ({1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_1692, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U16 ( .a ({1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_1691, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U15 ( .a ({1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_1659, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U14 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1658, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U13 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1657, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U12 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1690, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U11 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1656, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U10 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1667, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U9 ( .a ({1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1550, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U8 ( .a ({1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_1683, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U7 ( .a ({1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_1682, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U6 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1666, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U5 ( .a ({1'b0, 1'b1}), .b ({new_AGEMA_signal_1549, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U4 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1681, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U3 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1680, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U2 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1548, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_AddConstants_instance_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1546, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_U3 ( .a ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}), .b ({new_AGEMA_signal_1876, LED_128_Instance_SBox_Instance_0_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_U2 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1721, LED_128_Instance_SBox_Instance_0_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_U1 ( .a ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_1799, LED_128_Instance_SBox_Instance_0_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .a ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .b ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .a ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .a ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .c ({new_AGEMA_signal_1877, LED_128_Instance_SBox_Instance_0_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_1722, LED_128_Instance_SBox_Instance_0_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .a ({new_AGEMA_signal_1722, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}), .c ({new_AGEMA_signal_1878, LED_128_Instance_SBox_Instance_0_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_1802, LED_128_Instance_SBox_Instance_0_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .a ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .c ({new_AGEMA_signal_1879, LED_128_Instance_SBox_Instance_0_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_U3 ( .a ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}), .b ({new_AGEMA_signal_1881, LED_128_Instance_SBox_Instance_1_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_U2 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1745, LED_128_Instance_SBox_Instance_1_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_U1 ( .a ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_1803, LED_128_Instance_SBox_Instance_1_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .a ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .b ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .a ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .a ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_1882, LED_128_Instance_SBox_Instance_1_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_1806, LED_128_Instance_SBox_Instance_1_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .a ({new_AGEMA_signal_1806, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}), .c ({new_AGEMA_signal_1883, LED_128_Instance_SBox_Instance_1_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_1807, LED_128_Instance_SBox_Instance_1_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .a ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .c ({new_AGEMA_signal_1884, LED_128_Instance_SBox_Instance_1_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_U3 ( .a ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}), .b ({new_AGEMA_signal_1808, LED_128_Instance_SBox_Instance_2_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_U2 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1746, LED_128_Instance_SBox_Instance_2_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_U1 ( .a ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_1747, LED_128_Instance_SBox_Instance_2_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .a ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .b ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .a ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .a ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_1809, LED_128_Instance_SBox_Instance_2_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_1750, LED_128_Instance_SBox_Instance_2_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .a ({new_AGEMA_signal_1750, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}), .c ({new_AGEMA_signal_1810, LED_128_Instance_SBox_Instance_2_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_1751, LED_128_Instance_SBox_Instance_2_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .a ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_1811, LED_128_Instance_SBox_Instance_2_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_U3 ( .a ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}), .b ({new_AGEMA_signal_1813, LED_128_Instance_SBox_Instance_3_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_U2 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1752, LED_128_Instance_SBox_Instance_3_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_U1 ( .a ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_1753, LED_128_Instance_SBox_Instance_3_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .a ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .b ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .a ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .a ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_1814, LED_128_Instance_SBox_Instance_3_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_1756, LED_128_Instance_SBox_Instance_3_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .a ({new_AGEMA_signal_1756, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}), .c ({new_AGEMA_signal_1815, LED_128_Instance_SBox_Instance_3_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_1757, LED_128_Instance_SBox_Instance_3_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .a ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_1816, LED_128_Instance_SBox_Instance_3_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_U3 ( .a ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}), .b ({new_AGEMA_signal_1890, LED_128_Instance_SBox_Instance_4_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_U2 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1723, LED_128_Instance_SBox_Instance_4_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_U1 ( .a ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_1818, LED_128_Instance_SBox_Instance_4_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .a ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .b ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .a ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .a ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .c ({new_AGEMA_signal_1891, LED_128_Instance_SBox_Instance_4_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_1724, LED_128_Instance_SBox_Instance_4_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .a ({new_AGEMA_signal_1724, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}), .c ({new_AGEMA_signal_1892, LED_128_Instance_SBox_Instance_4_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_1821, LED_128_Instance_SBox_Instance_4_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .a ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .c ({new_AGEMA_signal_1893, LED_128_Instance_SBox_Instance_4_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_U3 ( .a ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}), .b ({new_AGEMA_signal_1895, LED_128_Instance_SBox_Instance_5_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_U2 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1758, LED_128_Instance_SBox_Instance_5_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_U1 ( .a ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_1822, LED_128_Instance_SBox_Instance_5_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .a ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .b ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .a ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .a ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_1896, LED_128_Instance_SBox_Instance_5_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_1825, LED_128_Instance_SBox_Instance_5_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .a ({new_AGEMA_signal_1825, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}), .c ({new_AGEMA_signal_1897, LED_128_Instance_SBox_Instance_5_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_1826, LED_128_Instance_SBox_Instance_5_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .a ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .c ({new_AGEMA_signal_1898, LED_128_Instance_SBox_Instance_5_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_U3 ( .a ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}), .b ({new_AGEMA_signal_1827, LED_128_Instance_SBox_Instance_6_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_U2 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1759, LED_128_Instance_SBox_Instance_6_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_U1 ( .a ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1760, LED_128_Instance_SBox_Instance_6_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .a ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .b ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .a ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .a ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_1828, LED_128_Instance_SBox_Instance_6_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_1763, LED_128_Instance_SBox_Instance_6_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .a ({new_AGEMA_signal_1763, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}), .c ({new_AGEMA_signal_1829, LED_128_Instance_SBox_Instance_6_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_1764, LED_128_Instance_SBox_Instance_6_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .a ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_1830, LED_128_Instance_SBox_Instance_6_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_U3 ( .a ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}), .b ({new_AGEMA_signal_1832, LED_128_Instance_SBox_Instance_7_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_U2 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1765, LED_128_Instance_SBox_Instance_7_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_U1 ( .a ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1766, LED_128_Instance_SBox_Instance_7_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .a ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .b ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .a ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .a ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_1833, LED_128_Instance_SBox_Instance_7_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_1769, LED_128_Instance_SBox_Instance_7_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .a ({new_AGEMA_signal_1769, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}), .c ({new_AGEMA_signal_1834, LED_128_Instance_SBox_Instance_7_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_1770, LED_128_Instance_SBox_Instance_7_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .a ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_1835, LED_128_Instance_SBox_Instance_7_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_U3 ( .a ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}), .b ({new_AGEMA_signal_1904, LED_128_Instance_SBox_Instance_8_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_U2 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1771, LED_128_Instance_SBox_Instance_8_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_U1 ( .a ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_1837, LED_128_Instance_SBox_Instance_8_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .a ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .b ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .a ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .a ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .c ({new_AGEMA_signal_1905, LED_128_Instance_SBox_Instance_8_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_1772, LED_128_Instance_SBox_Instance_8_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .a ({new_AGEMA_signal_1772, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}), .c ({new_AGEMA_signal_1906, LED_128_Instance_SBox_Instance_8_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_1840, LED_128_Instance_SBox_Instance_8_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .a ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .c ({new_AGEMA_signal_1907, LED_128_Instance_SBox_Instance_8_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_U3 ( .a ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}), .b ({new_AGEMA_signal_1909, LED_128_Instance_SBox_Instance_9_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_U2 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1725, LED_128_Instance_SBox_Instance_9_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_U1 ( .a ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_1841, LED_128_Instance_SBox_Instance_9_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .a ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .b ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .a ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .a ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_1910, LED_128_Instance_SBox_Instance_9_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_1773, LED_128_Instance_SBox_Instance_9_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .a ({new_AGEMA_signal_1773, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}), .c ({new_AGEMA_signal_1911, LED_128_Instance_SBox_Instance_9_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_1844, LED_128_Instance_SBox_Instance_9_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .a ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .c ({new_AGEMA_signal_1912, LED_128_Instance_SBox_Instance_9_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_U3 ( .a ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}), .b ({new_AGEMA_signal_1845, LED_128_Instance_SBox_Instance_10_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_U2 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1774, LED_128_Instance_SBox_Instance_10_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_U1 ( .a ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_1775, LED_128_Instance_SBox_Instance_10_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .a ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .b ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .a ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .a ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_1846, LED_128_Instance_SBox_Instance_10_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_1778, LED_128_Instance_SBox_Instance_10_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .a ({new_AGEMA_signal_1778, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}), .c ({new_AGEMA_signal_1847, LED_128_Instance_SBox_Instance_10_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_1779, LED_128_Instance_SBox_Instance_10_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .a ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_1848, LED_128_Instance_SBox_Instance_10_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_U3 ( .a ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}), .b ({new_AGEMA_signal_1850, LED_128_Instance_SBox_Instance_11_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_U2 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1780, LED_128_Instance_SBox_Instance_11_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_U1 ( .a ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_1781, LED_128_Instance_SBox_Instance_11_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .a ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .b ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .a ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .a ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_1851, LED_128_Instance_SBox_Instance_11_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_1784, LED_128_Instance_SBox_Instance_11_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .a ({new_AGEMA_signal_1784, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}), .c ({new_AGEMA_signal_1852, LED_128_Instance_SBox_Instance_11_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_1785, LED_128_Instance_SBox_Instance_11_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .a ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_1853, LED_128_Instance_SBox_Instance_11_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_U3 ( .a ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}), .b ({new_AGEMA_signal_1918, LED_128_Instance_SBox_Instance_12_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_U2 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1855, LED_128_Instance_SBox_Instance_12_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_U1 ( .a ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_1856, LED_128_Instance_SBox_Instance_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .a ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .b ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .a ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .a ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .c ({new_AGEMA_signal_1919, LED_128_Instance_SBox_Instance_12_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_1859, LED_128_Instance_SBox_Instance_12_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .a ({new_AGEMA_signal_1859, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}), .c ({new_AGEMA_signal_1920, LED_128_Instance_SBox_Instance_12_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_1860, LED_128_Instance_SBox_Instance_12_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .a ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .c ({new_AGEMA_signal_1921, LED_128_Instance_SBox_Instance_12_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_U3 ( .a ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}), .b ({new_AGEMA_signal_1923, LED_128_Instance_SBox_Instance_13_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_U2 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1786, LED_128_Instance_SBox_Instance_13_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_U1 ( .a ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_1861, LED_128_Instance_SBox_Instance_13_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .a ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .b ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .a ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .a ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_1924, LED_128_Instance_SBox_Instance_13_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_1864, LED_128_Instance_SBox_Instance_13_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .a ({new_AGEMA_signal_1864, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}), .c ({new_AGEMA_signal_1925, LED_128_Instance_SBox_Instance_13_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_1865, LED_128_Instance_SBox_Instance_13_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .a ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .c ({new_AGEMA_signal_1926, LED_128_Instance_SBox_Instance_13_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_U3 ( .a ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}), .b ({new_AGEMA_signal_1866, LED_128_Instance_SBox_Instance_14_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_U2 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1787, LED_128_Instance_SBox_Instance_14_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_U1 ( .a ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_1788, LED_128_Instance_SBox_Instance_14_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .a ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .b ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .a ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .a ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_1867, LED_128_Instance_SBox_Instance_14_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_1791, LED_128_Instance_SBox_Instance_14_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .a ({new_AGEMA_signal_1791, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}), .c ({new_AGEMA_signal_1868, LED_128_Instance_SBox_Instance_14_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_1792, LED_128_Instance_SBox_Instance_14_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .a ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_1869, LED_128_Instance_SBox_Instance_14_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_U3 ( .a ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}), .b ({new_AGEMA_signal_1871, LED_128_Instance_SBox_Instance_15_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_U2 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1793, LED_128_Instance_SBox_Instance_15_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_U1 ( .a ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_1794, LED_128_Instance_SBox_Instance_15_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .a ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .b ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .a ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .a ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_1872, LED_128_Instance_SBox_Instance_15_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_1797, LED_128_Instance_SBox_Instance_15_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .a ({new_AGEMA_signal_1797, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}), .c ({new_AGEMA_signal_1873, LED_128_Instance_SBox_Instance_15_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_1798, LED_128_Instance_SBox_Instance_15_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .a ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_1874, LED_128_Instance_SBox_Instance_15_Q7}) ) ;
    INV_X1 LED_128_Instance_ks_reg_0__U1 ( .A (LED_128_Instance_ks_reg_0__Q), .ZN (LED_128_Instance_n4) ) ;
    INV_X1 LED_128_Instance_ks_reg_1__U1 ( .A (LED_128_Instance_n26), .ZN (LED_128_Instance_n8) ) ;
    INV_X1 LED_128_Instance_ks_reg_2__U1 ( .A (LED_128_Instance_n25), .ZN (LED_128_Instance_n1) ) ;
    INV_X1 LED_128_Instance_ks_reg_3__U1 ( .A (LED_128_Instance_n2), .ZN (LED_128_Instance_n24) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_0__U1 ( .A (roundconstant[0]), .ZN (LED_128_Instance_n6) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_1__U1 ( .A (roundconstant[1]), .ZN (LED_128_Instance_n29) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_2__U1 ( .A (roundconstant[2]), .ZN (LED_128_Instance_n5) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_3__U1 ( .A (roundconstant[3]), .ZN (LED_128_Instance_n30) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_4__U1 ( .A (roundconstant[4]), .ZN (LED_128_Instance_n28) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_5__U1 ( .A (roundconstant[5]), .ZN (LED_128_Instance_n27) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (CLK), .rst (IN_reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .a ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_1877, LED_128_Instance_SBox_Instance_0_L2}), .c ({new_AGEMA_signal_1964, LED_128_Instance_SBox_Instance_0_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .a ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .a ({new_AGEMA_signal_1802, LED_128_Instance_SBox_Instance_0_L4}), .b ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}), .c ({new_AGEMA_signal_1996, LED_128_Instance_SBox_Instance_0_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .a ({new_AGEMA_signal_1876, LED_128_Instance_SBox_Instance_0_n1}), .b ({new_AGEMA_signal_1721, LED_128_Instance_SBox_Instance_0_n2}), .clk (CLK), .r (Fresh[0]), .c ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .a ({new_AGEMA_signal_1799, LED_128_Instance_SBox_Instance_0_n3}), .b ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .clk (CLK), .r (Fresh[1]), .c ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .a ({new_AGEMA_signal_1722, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_1933, LED_128_Instance_subcells_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .a ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_1882, LED_128_Instance_SBox_Instance_1_L2}), .c ({new_AGEMA_signal_1966, LED_128_Instance_SBox_Instance_1_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .a ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .a ({new_AGEMA_signal_1807, LED_128_Instance_SBox_Instance_1_L4}), .b ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}), .c ({new_AGEMA_signal_1998, LED_128_Instance_SBox_Instance_1_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .a ({new_AGEMA_signal_1881, LED_128_Instance_SBox_Instance_1_n1}), .b ({new_AGEMA_signal_1745, LED_128_Instance_SBox_Instance_1_n2}), .clk (CLK), .r (Fresh[2]), .c ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .a ({new_AGEMA_signal_1803, LED_128_Instance_SBox_Instance_1_n3}), .b ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .clk (CLK), .r (Fresh[3]), .c ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .a ({new_AGEMA_signal_1806, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_1935, LED_128_Instance_subcells_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .a ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_1809, LED_128_Instance_SBox_Instance_2_L2}), .c ({new_AGEMA_signal_1936, LED_128_Instance_SBox_Instance_2_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .a ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .a ({new_AGEMA_signal_1751, LED_128_Instance_SBox_Instance_2_L4}), .b ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}), .c ({new_AGEMA_signal_1968, LED_128_Instance_SBox_Instance_2_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .a ({new_AGEMA_signal_1808, LED_128_Instance_SBox_Instance_2_n1}), .b ({new_AGEMA_signal_1746, LED_128_Instance_SBox_Instance_2_n2}), .clk (CLK), .r (Fresh[4]), .c ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .a ({new_AGEMA_signal_1747, LED_128_Instance_SBox_Instance_2_n3}), .b ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .clk (CLK), .r (Fresh[5]), .c ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .a ({new_AGEMA_signal_1750, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_1887, LED_128_Instance_subcells_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .a ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_1814, LED_128_Instance_SBox_Instance_3_L2}), .c ({new_AGEMA_signal_1938, LED_128_Instance_SBox_Instance_3_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .a ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .a ({new_AGEMA_signal_1757, LED_128_Instance_SBox_Instance_3_L4}), .b ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}), .c ({new_AGEMA_signal_1970, LED_128_Instance_SBox_Instance_3_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .a ({new_AGEMA_signal_1813, LED_128_Instance_SBox_Instance_3_n1}), .b ({new_AGEMA_signal_1752, LED_128_Instance_SBox_Instance_3_n2}), .clk (CLK), .r (Fresh[6]), .c ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .a ({new_AGEMA_signal_1753, LED_128_Instance_SBox_Instance_3_n3}), .b ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .clk (CLK), .r (Fresh[7]), .c ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .a ({new_AGEMA_signal_1756, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_1889, LED_128_Instance_subcells_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .a ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_1891, LED_128_Instance_SBox_Instance_4_L2}), .c ({new_AGEMA_signal_1972, LED_128_Instance_SBox_Instance_4_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .a ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .a ({new_AGEMA_signal_1821, LED_128_Instance_SBox_Instance_4_L4}), .b ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}), .c ({new_AGEMA_signal_2004, LED_128_Instance_SBox_Instance_4_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .a ({new_AGEMA_signal_1890, LED_128_Instance_SBox_Instance_4_n1}), .b ({new_AGEMA_signal_1723, LED_128_Instance_SBox_Instance_4_n2}), .clk (CLK), .r (Fresh[8]), .c ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .a ({new_AGEMA_signal_1818, LED_128_Instance_SBox_Instance_4_n3}), .b ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .clk (CLK), .r (Fresh[9]), .c ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .a ({new_AGEMA_signal_1724, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_1941, LED_128_Instance_subcells_out[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .a ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_1896, LED_128_Instance_SBox_Instance_5_L2}), .c ({new_AGEMA_signal_1974, LED_128_Instance_SBox_Instance_5_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .a ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .a ({new_AGEMA_signal_1826, LED_128_Instance_SBox_Instance_5_L4}), .b ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}), .c ({new_AGEMA_signal_2006, LED_128_Instance_SBox_Instance_5_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .a ({new_AGEMA_signal_1895, LED_128_Instance_SBox_Instance_5_n1}), .b ({new_AGEMA_signal_1758, LED_128_Instance_SBox_Instance_5_n2}), .clk (CLK), .r (Fresh[10]), .c ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .a ({new_AGEMA_signal_1822, LED_128_Instance_SBox_Instance_5_n3}), .b ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .clk (CLK), .r (Fresh[11]), .c ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .a ({new_AGEMA_signal_1825, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_1943, LED_128_Instance_subcells_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .a ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_1828, LED_128_Instance_SBox_Instance_6_L2}), .c ({new_AGEMA_signal_1944, LED_128_Instance_SBox_Instance_6_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .a ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .a ({new_AGEMA_signal_1764, LED_128_Instance_SBox_Instance_6_L4}), .b ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}), .c ({new_AGEMA_signal_1976, LED_128_Instance_SBox_Instance_6_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .a ({new_AGEMA_signal_1827, LED_128_Instance_SBox_Instance_6_n1}), .b ({new_AGEMA_signal_1759, LED_128_Instance_SBox_Instance_6_n2}), .clk (CLK), .r (Fresh[12]), .c ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .a ({new_AGEMA_signal_1760, LED_128_Instance_SBox_Instance_6_n3}), .b ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .clk (CLK), .r (Fresh[13]), .c ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .a ({new_AGEMA_signal_1763, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_1901, LED_128_Instance_subcells_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .a ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_1833, LED_128_Instance_SBox_Instance_7_L2}), .c ({new_AGEMA_signal_1946, LED_128_Instance_SBox_Instance_7_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .a ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .a ({new_AGEMA_signal_1770, LED_128_Instance_SBox_Instance_7_L4}), .b ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}), .c ({new_AGEMA_signal_1978, LED_128_Instance_SBox_Instance_7_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .a ({new_AGEMA_signal_1832, LED_128_Instance_SBox_Instance_7_n1}), .b ({new_AGEMA_signal_1765, LED_128_Instance_SBox_Instance_7_n2}), .clk (CLK), .r (Fresh[14]), .c ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .a ({new_AGEMA_signal_1766, LED_128_Instance_SBox_Instance_7_n3}), .b ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .clk (CLK), .r (Fresh[15]), .c ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .a ({new_AGEMA_signal_1769, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_1903, LED_128_Instance_subcells_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .a ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_1905, LED_128_Instance_SBox_Instance_8_L2}), .c ({new_AGEMA_signal_1980, LED_128_Instance_SBox_Instance_8_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .a ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .a ({new_AGEMA_signal_1840, LED_128_Instance_SBox_Instance_8_L4}), .b ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}), .c ({new_AGEMA_signal_2012, LED_128_Instance_SBox_Instance_8_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .a ({new_AGEMA_signal_1904, LED_128_Instance_SBox_Instance_8_n1}), .b ({new_AGEMA_signal_1771, LED_128_Instance_SBox_Instance_8_n2}), .clk (CLK), .r (Fresh[16]), .c ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .a ({new_AGEMA_signal_1837, LED_128_Instance_SBox_Instance_8_n3}), .b ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .clk (CLK), .r (Fresh[17]), .c ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .a ({new_AGEMA_signal_1772, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_1949, LED_128_Instance_subcells_out[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .a ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_1910, LED_128_Instance_SBox_Instance_9_L2}), .c ({new_AGEMA_signal_1982, LED_128_Instance_SBox_Instance_9_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .a ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .a ({new_AGEMA_signal_1844, LED_128_Instance_SBox_Instance_9_L4}), .b ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}), .c ({new_AGEMA_signal_2014, LED_128_Instance_SBox_Instance_9_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .a ({new_AGEMA_signal_1909, LED_128_Instance_SBox_Instance_9_n1}), .b ({new_AGEMA_signal_1725, LED_128_Instance_SBox_Instance_9_n2}), .clk (CLK), .r (Fresh[18]), .c ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .a ({new_AGEMA_signal_1841, LED_128_Instance_SBox_Instance_9_n3}), .b ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .clk (CLK), .r (Fresh[19]), .c ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .a ({new_AGEMA_signal_1773, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_1951, LED_128_Instance_subcells_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .a ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_1846, LED_128_Instance_SBox_Instance_10_L2}), .c ({new_AGEMA_signal_1952, LED_128_Instance_SBox_Instance_10_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .a ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .a ({new_AGEMA_signal_1779, LED_128_Instance_SBox_Instance_10_L4}), .b ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}), .c ({new_AGEMA_signal_1984, LED_128_Instance_SBox_Instance_10_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .a ({new_AGEMA_signal_1845, LED_128_Instance_SBox_Instance_10_n1}), .b ({new_AGEMA_signal_1774, LED_128_Instance_SBox_Instance_10_n2}), .clk (CLK), .r (Fresh[20]), .c ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .a ({new_AGEMA_signal_1775, LED_128_Instance_SBox_Instance_10_n3}), .b ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .clk (CLK), .r (Fresh[21]), .c ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .a ({new_AGEMA_signal_1778, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_1915, LED_128_Instance_subcells_out[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .a ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_1851, LED_128_Instance_SBox_Instance_11_L2}), .c ({new_AGEMA_signal_1954, LED_128_Instance_SBox_Instance_11_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .a ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .a ({new_AGEMA_signal_1785, LED_128_Instance_SBox_Instance_11_L4}), .b ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}), .c ({new_AGEMA_signal_1986, LED_128_Instance_SBox_Instance_11_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .a ({new_AGEMA_signal_1850, LED_128_Instance_SBox_Instance_11_n1}), .b ({new_AGEMA_signal_1780, LED_128_Instance_SBox_Instance_11_n2}), .clk (CLK), .r (Fresh[22]), .c ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .a ({new_AGEMA_signal_1781, LED_128_Instance_SBox_Instance_11_n3}), .b ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .clk (CLK), .r (Fresh[23]), .c ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .a ({new_AGEMA_signal_1784, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_1917, LED_128_Instance_subcells_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .a ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_1919, LED_128_Instance_SBox_Instance_12_L2}), .c ({new_AGEMA_signal_1988, LED_128_Instance_SBox_Instance_12_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .a ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .a ({new_AGEMA_signal_1860, LED_128_Instance_SBox_Instance_12_L4}), .b ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}), .c ({new_AGEMA_signal_2020, LED_128_Instance_SBox_Instance_12_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .a ({new_AGEMA_signal_1918, LED_128_Instance_SBox_Instance_12_n1}), .b ({new_AGEMA_signal_1855, LED_128_Instance_SBox_Instance_12_n2}), .clk (CLK), .r (Fresh[24]), .c ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .a ({new_AGEMA_signal_1856, LED_128_Instance_SBox_Instance_12_n3}), .b ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .clk (CLK), .r (Fresh[25]), .c ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .a ({new_AGEMA_signal_1859, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_1957, LED_128_Instance_subcells_out[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .a ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_1924, LED_128_Instance_SBox_Instance_13_L2}), .c ({new_AGEMA_signal_1990, LED_128_Instance_SBox_Instance_13_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .a ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .a ({new_AGEMA_signal_1865, LED_128_Instance_SBox_Instance_13_L4}), .b ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}), .c ({new_AGEMA_signal_2022, LED_128_Instance_SBox_Instance_13_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .a ({new_AGEMA_signal_1923, LED_128_Instance_SBox_Instance_13_n1}), .b ({new_AGEMA_signal_1786, LED_128_Instance_SBox_Instance_13_n2}), .clk (CLK), .r (Fresh[26]), .c ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .a ({new_AGEMA_signal_1861, LED_128_Instance_SBox_Instance_13_n3}), .b ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .clk (CLK), .r (Fresh[27]), .c ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .a ({new_AGEMA_signal_1864, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_1959, LED_128_Instance_subcells_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .a ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_1867, LED_128_Instance_SBox_Instance_14_L2}), .c ({new_AGEMA_signal_1960, LED_128_Instance_SBox_Instance_14_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .a ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .a ({new_AGEMA_signal_1792, LED_128_Instance_SBox_Instance_14_L4}), .b ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}), .c ({new_AGEMA_signal_1992, LED_128_Instance_SBox_Instance_14_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .a ({new_AGEMA_signal_1866, LED_128_Instance_SBox_Instance_14_n1}), .b ({new_AGEMA_signal_1787, LED_128_Instance_SBox_Instance_14_n2}), .clk (CLK), .r (Fresh[28]), .c ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .a ({new_AGEMA_signal_1788, LED_128_Instance_SBox_Instance_14_n3}), .b ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .clk (CLK), .r (Fresh[29]), .c ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .a ({new_AGEMA_signal_1791, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_1929, LED_128_Instance_subcells_out[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .a ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_1872, LED_128_Instance_SBox_Instance_15_L2}), .c ({new_AGEMA_signal_1962, LED_128_Instance_SBox_Instance_15_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .a ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .a ({new_AGEMA_signal_1798, LED_128_Instance_SBox_Instance_15_L4}), .b ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}), .c ({new_AGEMA_signal_1994, LED_128_Instance_SBox_Instance_15_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .a ({new_AGEMA_signal_1871, LED_128_Instance_SBox_Instance_15_n1}), .b ({new_AGEMA_signal_1793, LED_128_Instance_SBox_Instance_15_n2}), .clk (CLK), .r (Fresh[30]), .c ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .a ({new_AGEMA_signal_1794, LED_128_Instance_SBox_Instance_15_n3}), .b ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .clk (CLK), .r (Fresh[31]), .c ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .a ({new_AGEMA_signal_1797, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_1931, LED_128_Instance_subcells_out[60]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_0_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .a ({new_AGEMA_signal_1546, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_2171, LED_128_Instance_state0[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_1_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .a ({new_AGEMA_signal_1666, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_2268, LED_128_Instance_state0[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_2_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .a ({new_AGEMA_signal_1667, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_2191, LED_128_Instance_state0[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_3_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .a ({new_AGEMA_signal_1547, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_2222, LED_128_Instance_state0[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .a ({new_AGEMA_signal_1668, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_2192, LED_128_Instance_state0[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .a ({new_AGEMA_signal_1669, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_2269, LED_128_Instance_state0[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .a ({new_AGEMA_signal_1670, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_2193, LED_128_Instance_state0[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_2194, LED_128_Instance_state0[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .a ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_2195, LED_128_Instance_state0[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .a ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_2223, LED_128_Instance_state0[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .a ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_2196, LED_128_Instance_state0[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_2197, LED_128_Instance_state0[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .a ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_2198, LED_128_Instance_state0[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .a ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_2224, LED_128_Instance_state0[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .a ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_2199, LED_128_Instance_state0[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_2225, LED_128_Instance_state0[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_16_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}), .a ({new_AGEMA_signal_1548, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_2310, LED_128_Instance_state0[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_17_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2340, LED_128_Instance_mixcolumns_out[17]}), .a ({new_AGEMA_signal_1680, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_2355, LED_128_Instance_state0[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_18_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .a ({new_AGEMA_signal_1681, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_2356, LED_128_Instance_state0[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_19_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .a ({new_AGEMA_signal_1549, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_2270, LED_128_Instance_state0[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}), .a ({new_AGEMA_signal_1682, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_2271, LED_128_Instance_state0[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_21_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2297, LED_128_Instance_mixcolumns_out[21]}), .a ({new_AGEMA_signal_1683, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_2311, LED_128_Instance_state0[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_22_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .a ({new_AGEMA_signal_1550, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_2357, LED_128_Instance_state0[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_23_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_2272, LED_128_Instance_state0[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_24_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}), .a ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_2273, LED_128_Instance_state0[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_25_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2304, LED_128_Instance_mixcolumns_out[25]}), .a ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_2312, LED_128_Instance_state0[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_26_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .a ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_2313, LED_128_Instance_state0[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_27_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_2274, LED_128_Instance_state0[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_28_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}), .a ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_2314, LED_128_Instance_state0[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2354, LED_128_Instance_mixcolumns_out[29]}), .a ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_2358, LED_128_Instance_state0[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .a ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_2315, LED_128_Instance_state0[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_2275, LED_128_Instance_state0[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_32_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}), .a ({new_AGEMA_signal_1656, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_2359, LED_128_Instance_state0[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}), .a ({new_AGEMA_signal_1690, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_2395, LED_128_Instance_state0[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_34_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}), .a ({new_AGEMA_signal_1657, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_2360, LED_128_Instance_state0[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_35_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}), .a ({new_AGEMA_signal_1658, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_2435, LED_128_Instance_state0[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_36_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}), .a ({new_AGEMA_signal_1659, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_2361, LED_128_Instance_state0[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_37_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}), .a ({new_AGEMA_signal_1691, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_2362, LED_128_Instance_state0[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}), .a ({new_AGEMA_signal_1692, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_2316, LED_128_Instance_state0[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_39_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}), .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_2436, LED_128_Instance_state0[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}), .a ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_2363, LED_128_Instance_state0[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}), .a ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_2364, LED_128_Instance_state0[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}), .a ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_2317, LED_128_Instance_state0[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_43_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}), .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_2396, LED_128_Instance_state0[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}), .a ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_2365, LED_128_Instance_state0[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}), .a ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_2397, LED_128_Instance_state0[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}), .a ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_2366, LED_128_Instance_state0[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_47_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}), .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_2398, LED_128_Instance_state0[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_48_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2487, LED_128_Instance_mixcolumns_out[48]}), .a ({new_AGEMA_signal_1701, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_2492, LED_128_Instance_state0[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_49_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2500, LED_128_Instance_mixcolumns_out[49]}), .a ({new_AGEMA_signal_1702, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_2502, LED_128_Instance_state0[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_50_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2427, LED_128_Instance_mixcolumns_out[50]}), .a ({new_AGEMA_signal_1703, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_2437, LED_128_Instance_state0[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_51_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2426, LED_128_Instance_mixcolumns_out[51]}), .a ({new_AGEMA_signal_1704, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_2438, LED_128_Instance_state0[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_52_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2489, LED_128_Instance_mixcolumns_out[52]}), .a ({new_AGEMA_signal_1705, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_2493, LED_128_Instance_state0[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_53_U1 ( .s (LED_128_Instance_n22), .b ({new_AGEMA_signal_2501, LED_128_Instance_mixcolumns_out[53]}), .a ({new_AGEMA_signal_1706, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_2503, LED_128_Instance_state0[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2387, LED_128_Instance_mixcolumns_out[54]}), .a ({new_AGEMA_signal_1707, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_2399, LED_128_Instance_state0[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2429, LED_128_Instance_mixcolumns_out[55]}), .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_2439, LED_128_Instance_state0[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2481, LED_128_Instance_mixcolumns_out[56]}), .a ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_2484, LED_128_Instance_state0[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2490, LED_128_Instance_mixcolumns_out[57]}), .a ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_2494, LED_128_Instance_state0[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2390, LED_128_Instance_mixcolumns_out[58]}), .a ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_2400, LED_128_Instance_state0[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2389, LED_128_Instance_mixcolumns_out[59]}), .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_2401, LED_128_Instance_state0[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_state0_n9), .b ({new_AGEMA_signal_2483, LED_128_Instance_mixcolumns_out[60]}), .a ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_2485, LED_128_Instance_state0[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_state0_n10), .b ({new_AGEMA_signal_2491, LED_128_Instance_mixcolumns_out[61]}), .a ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_2495, LED_128_Instance_state0[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2433, LED_128_Instance_mixcolumns_out[62]}), .a ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_2440, LED_128_Instance_state0[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state0_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_state0_n8), .b ({new_AGEMA_signal_2432, LED_128_Instance_mixcolumns_out[63]}), .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_2441, LED_128_Instance_state0[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_0_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2171, LED_128_Instance_state0[0]}), .a ({IN_plaintext_s1[0], IN_plaintext_s0[0]}), .c ({new_AGEMA_signal_2201, LED_128_Instance_state1[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_1_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2268, LED_128_Instance_state0[1]}), .a ({IN_plaintext_s1[1], IN_plaintext_s0[1]}), .c ({new_AGEMA_signal_2319, LED_128_Instance_state1[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_2_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2191, LED_128_Instance_state0[2]}), .a ({IN_plaintext_s1[2], IN_plaintext_s0[2]}), .c ({new_AGEMA_signal_2227, LED_128_Instance_state1[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_3_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2222, LED_128_Instance_state0[3]}), .a ({IN_plaintext_s1[3], IN_plaintext_s0[3]}), .c ({new_AGEMA_signal_2277, LED_128_Instance_state1[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_4_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2192, LED_128_Instance_state0[4]}), .a ({IN_plaintext_s1[4], IN_plaintext_s0[4]}), .c ({new_AGEMA_signal_2229, LED_128_Instance_state1[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_5_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2269, LED_128_Instance_state0[5]}), .a ({IN_plaintext_s1[5], IN_plaintext_s0[5]}), .c ({new_AGEMA_signal_2321, LED_128_Instance_state1[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_6_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2193, LED_128_Instance_state0[6]}), .a ({IN_plaintext_s1[6], IN_plaintext_s0[6]}), .c ({new_AGEMA_signal_2231, LED_128_Instance_state1[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_7_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2194, LED_128_Instance_state0[7]}), .a ({IN_plaintext_s1[7], IN_plaintext_s0[7]}), .c ({new_AGEMA_signal_2233, LED_128_Instance_state1[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_8_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2195, LED_128_Instance_state0[8]}), .a ({IN_plaintext_s1[8], IN_plaintext_s0[8]}), .c ({new_AGEMA_signal_2235, LED_128_Instance_state1[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_9_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2223, LED_128_Instance_state0[9]}), .a ({IN_plaintext_s1[9], IN_plaintext_s0[9]}), .c ({new_AGEMA_signal_2279, LED_128_Instance_state1[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_10_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2196, LED_128_Instance_state0[10]}), .a ({IN_plaintext_s1[10], IN_plaintext_s0[10]}), .c ({new_AGEMA_signal_2237, LED_128_Instance_state1[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_11_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2197, LED_128_Instance_state0[11]}), .a ({IN_plaintext_s1[11], IN_plaintext_s0[11]}), .c ({new_AGEMA_signal_2239, LED_128_Instance_state1[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_12_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2198, LED_128_Instance_state0[12]}), .a ({IN_plaintext_s1[12], IN_plaintext_s0[12]}), .c ({new_AGEMA_signal_2241, LED_128_Instance_state1[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_13_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2224, LED_128_Instance_state0[13]}), .a ({IN_plaintext_s1[13], IN_plaintext_s0[13]}), .c ({new_AGEMA_signal_2281, LED_128_Instance_state1[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_14_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2199, LED_128_Instance_state0[14]}), .a ({IN_plaintext_s1[14], IN_plaintext_s0[14]}), .c ({new_AGEMA_signal_2243, LED_128_Instance_state1[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_15_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2225, LED_128_Instance_state0[15]}), .a ({IN_plaintext_s1[15], IN_plaintext_s0[15]}), .c ({new_AGEMA_signal_2283, LED_128_Instance_state1[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_16_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2310, LED_128_Instance_state0[16]}), .a ({IN_plaintext_s1[16], IN_plaintext_s0[16]}), .c ({new_AGEMA_signal_2368, LED_128_Instance_state1[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_17_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2355, LED_128_Instance_state0[17]}), .a ({IN_plaintext_s1[17], IN_plaintext_s0[17]}), .c ({new_AGEMA_signal_2403, LED_128_Instance_state1[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_18_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2356, LED_128_Instance_state0[18]}), .a ({IN_plaintext_s1[18], IN_plaintext_s0[18]}), .c ({new_AGEMA_signal_2405, LED_128_Instance_state1[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_19_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2270, LED_128_Instance_state0[19]}), .a ({IN_plaintext_s1[19], IN_plaintext_s0[19]}), .c ({new_AGEMA_signal_2323, LED_128_Instance_state1[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_20_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2271, LED_128_Instance_state0[20]}), .a ({IN_plaintext_s1[20], IN_plaintext_s0[20]}), .c ({new_AGEMA_signal_2325, LED_128_Instance_state1[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_21_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2311, LED_128_Instance_state0[21]}), .a ({IN_plaintext_s1[21], IN_plaintext_s0[21]}), .c ({new_AGEMA_signal_2370, LED_128_Instance_state1[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_22_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2357, LED_128_Instance_state0[22]}), .a ({IN_plaintext_s1[22], IN_plaintext_s0[22]}), .c ({new_AGEMA_signal_2407, LED_128_Instance_state1[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_23_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2272, LED_128_Instance_state0[23]}), .a ({IN_plaintext_s1[23], IN_plaintext_s0[23]}), .c ({new_AGEMA_signal_2327, LED_128_Instance_state1[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_24_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2273, LED_128_Instance_state0[24]}), .a ({IN_plaintext_s1[24], IN_plaintext_s0[24]}), .c ({new_AGEMA_signal_2329, LED_128_Instance_state1[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_25_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2312, LED_128_Instance_state0[25]}), .a ({IN_plaintext_s1[25], IN_plaintext_s0[25]}), .c ({new_AGEMA_signal_2372, LED_128_Instance_state1[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_26_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2313, LED_128_Instance_state0[26]}), .a ({IN_plaintext_s1[26], IN_plaintext_s0[26]}), .c ({new_AGEMA_signal_2374, LED_128_Instance_state1[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_27_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2274, LED_128_Instance_state0[27]}), .a ({IN_plaintext_s1[27], IN_plaintext_s0[27]}), .c ({new_AGEMA_signal_2331, LED_128_Instance_state1[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_28_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2314, LED_128_Instance_state0[28]}), .a ({IN_plaintext_s1[28], IN_plaintext_s0[28]}), .c ({new_AGEMA_signal_2376, LED_128_Instance_state1[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_29_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2358, LED_128_Instance_state0[29]}), .a ({IN_plaintext_s1[29], IN_plaintext_s0[29]}), .c ({new_AGEMA_signal_2409, LED_128_Instance_state1[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_30_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2315, LED_128_Instance_state0[30]}), .a ({IN_plaintext_s1[30], IN_plaintext_s0[30]}), .c ({new_AGEMA_signal_2378, LED_128_Instance_state1[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_31_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2275, LED_128_Instance_state0[31]}), .a ({IN_plaintext_s1[31], IN_plaintext_s0[31]}), .c ({new_AGEMA_signal_2333, LED_128_Instance_state1[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_32_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2359, LED_128_Instance_state0[32]}), .a ({IN_plaintext_s1[32], IN_plaintext_s0[32]}), .c ({new_AGEMA_signal_2411, LED_128_Instance_state1[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_33_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2395, LED_128_Instance_state0[33]}), .a ({IN_plaintext_s1[33], IN_plaintext_s0[33]}), .c ({new_AGEMA_signal_2443, LED_128_Instance_state1[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_34_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2360, LED_128_Instance_state0[34]}), .a ({IN_plaintext_s1[34], IN_plaintext_s0[34]}), .c ({new_AGEMA_signal_2413, LED_128_Instance_state1[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_35_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2435, LED_128_Instance_state0[35]}), .a ({IN_plaintext_s1[35], IN_plaintext_s0[35]}), .c ({new_AGEMA_signal_2463, LED_128_Instance_state1[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_36_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2361, LED_128_Instance_state0[36]}), .a ({IN_plaintext_s1[36], IN_plaintext_s0[36]}), .c ({new_AGEMA_signal_2415, LED_128_Instance_state1[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_37_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2362, LED_128_Instance_state0[37]}), .a ({IN_plaintext_s1[37], IN_plaintext_s0[37]}), .c ({new_AGEMA_signal_2417, LED_128_Instance_state1[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_38_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2316, LED_128_Instance_state0[38]}), .a ({IN_plaintext_s1[38], IN_plaintext_s0[38]}), .c ({new_AGEMA_signal_2380, LED_128_Instance_state1[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_39_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2436, LED_128_Instance_state0[39]}), .a ({IN_plaintext_s1[39], IN_plaintext_s0[39]}), .c ({new_AGEMA_signal_2465, LED_128_Instance_state1[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_40_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2363, LED_128_Instance_state0[40]}), .a ({IN_plaintext_s1[40], IN_plaintext_s0[40]}), .c ({new_AGEMA_signal_2419, LED_128_Instance_state1[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_41_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2364, LED_128_Instance_state0[41]}), .a ({IN_plaintext_s1[41], IN_plaintext_s0[41]}), .c ({new_AGEMA_signal_2421, LED_128_Instance_state1[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_42_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2317, LED_128_Instance_state0[42]}), .a ({IN_plaintext_s1[42], IN_plaintext_s0[42]}), .c ({new_AGEMA_signal_2382, LED_128_Instance_state1[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_43_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2396, LED_128_Instance_state0[43]}), .a ({IN_plaintext_s1[43], IN_plaintext_s0[43]}), .c ({new_AGEMA_signal_2445, LED_128_Instance_state1[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_44_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2365, LED_128_Instance_state0[44]}), .a ({IN_plaintext_s1[44], IN_plaintext_s0[44]}), .c ({new_AGEMA_signal_2423, LED_128_Instance_state1[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_45_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2397, LED_128_Instance_state0[45]}), .a ({IN_plaintext_s1[45], IN_plaintext_s0[45]}), .c ({new_AGEMA_signal_2447, LED_128_Instance_state1[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_46_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2366, LED_128_Instance_state0[46]}), .a ({IN_plaintext_s1[46], IN_plaintext_s0[46]}), .c ({new_AGEMA_signal_2425, LED_128_Instance_state1[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_47_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2398, LED_128_Instance_state0[47]}), .a ({IN_plaintext_s1[47], IN_plaintext_s0[47]}), .c ({new_AGEMA_signal_2449, LED_128_Instance_state1[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_48_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2492, LED_128_Instance_state0[48]}), .a ({IN_plaintext_s1[48], IN_plaintext_s0[48]}), .c ({new_AGEMA_signal_2505, LED_128_Instance_state1[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_49_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2502, LED_128_Instance_state0[49]}), .a ({IN_plaintext_s1[49], IN_plaintext_s0[49]}), .c ({new_AGEMA_signal_2513, LED_128_Instance_state1[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_50_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2437, LED_128_Instance_state0[50]}), .a ({IN_plaintext_s1[50], IN_plaintext_s0[50]}), .c ({new_AGEMA_signal_2467, LED_128_Instance_state1[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_51_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2438, LED_128_Instance_state0[51]}), .a ({IN_plaintext_s1[51], IN_plaintext_s0[51]}), .c ({new_AGEMA_signal_2469, LED_128_Instance_state1[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_52_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2493, LED_128_Instance_state0[52]}), .a ({IN_plaintext_s1[52], IN_plaintext_s0[52]}), .c ({new_AGEMA_signal_2507, LED_128_Instance_state1[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_53_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2503, LED_128_Instance_state0[53]}), .a ({IN_plaintext_s1[53], IN_plaintext_s0[53]}), .c ({new_AGEMA_signal_2515, LED_128_Instance_state1[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_54_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2399, LED_128_Instance_state0[54]}), .a ({IN_plaintext_s1[54], IN_plaintext_s0[54]}), .c ({new_AGEMA_signal_2451, LED_128_Instance_state1[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_55_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2439, LED_128_Instance_state0[55]}), .a ({IN_plaintext_s1[55], IN_plaintext_s0[55]}), .c ({new_AGEMA_signal_2471, LED_128_Instance_state1[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_56_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2484, LED_128_Instance_state0[56]}), .a ({IN_plaintext_s1[56], IN_plaintext_s0[56]}), .c ({new_AGEMA_signal_2497, LED_128_Instance_state1[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_57_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2494, LED_128_Instance_state0[57]}), .a ({IN_plaintext_s1[57], IN_plaintext_s0[57]}), .c ({new_AGEMA_signal_2509, LED_128_Instance_state1[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_58_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2400, LED_128_Instance_state0[58]}), .a ({IN_plaintext_s1[58], IN_plaintext_s0[58]}), .c ({new_AGEMA_signal_2453, LED_128_Instance_state1[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_59_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2401, LED_128_Instance_state0[59]}), .a ({IN_plaintext_s1[59], IN_plaintext_s0[59]}), .c ({new_AGEMA_signal_2455, LED_128_Instance_state1[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_60_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2485, LED_128_Instance_state0[60]}), .a ({IN_plaintext_s1[60], IN_plaintext_s0[60]}), .c ({new_AGEMA_signal_2499, LED_128_Instance_state1[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_61_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2495, LED_128_Instance_state0[61]}), .a ({IN_plaintext_s1[61], IN_plaintext_s0[61]}), .c ({new_AGEMA_signal_2511, LED_128_Instance_state1[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_62_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2440, LED_128_Instance_state0[62]}), .a ({IN_plaintext_s1[62], IN_plaintext_s0[62]}), .c ({new_AGEMA_signal_2473, LED_128_Instance_state1[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_MUX_state1_mux_inst_63_U1 ( .s (IN_reset), .b ({new_AGEMA_signal_2441, LED_128_Instance_state0[63]}), .a ({IN_plaintext_s1[63], IN_plaintext_s0[63]}), .c ({new_AGEMA_signal_2475, LED_128_Instance_state1[63]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .a ({new_AGEMA_signal_1964, LED_128_Instance_SBox_Instance_0_Q2}), .b ({new_AGEMA_signal_1878, LED_128_Instance_SBox_Instance_0_Q3}), .clk (CLK), .r (Fresh[32]), .c ({new_AGEMA_signal_1997, LED_128_Instance_SBox_Instance_0_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .a ({new_AGEMA_signal_1996, LED_128_Instance_SBox_Instance_0_Q6}), .b ({new_AGEMA_signal_1879, LED_128_Instance_SBox_Instance_0_Q7}), .clk (CLK), .r (Fresh[33]), .c ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .a ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}), .b ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2068, LED_128_Instance_SBox_Instance_0_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .a ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}), .b ({new_AGEMA_signal_2068, LED_128_Instance_SBox_Instance_0_L7}), .c ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .a ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}), .b ({new_AGEMA_signal_1997, LED_128_Instance_SBox_Instance_0_T1}), .c ({new_AGEMA_signal_2029, LED_128_Instance_SBox_Instance_0_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .a ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_2029, LED_128_Instance_SBox_Instance_0_L8}), .c ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .a ({new_AGEMA_signal_1802, LED_128_Instance_SBox_Instance_0_L4}), .b ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2070, LED_128_Instance_subcells_out[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .a ({new_AGEMA_signal_1966, LED_128_Instance_SBox_Instance_1_Q2}), .b ({new_AGEMA_signal_1883, LED_128_Instance_SBox_Instance_1_Q3}), .clk (CLK), .r (Fresh[34]), .c ({new_AGEMA_signal_1999, LED_128_Instance_SBox_Instance_1_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .a ({new_AGEMA_signal_1998, LED_128_Instance_SBox_Instance_1_Q6}), .b ({new_AGEMA_signal_1884, LED_128_Instance_SBox_Instance_1_Q7}), .clk (CLK), .r (Fresh[35]), .c ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .a ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}), .b ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2071, LED_128_Instance_SBox_Instance_1_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .a ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}), .b ({new_AGEMA_signal_2071, LED_128_Instance_SBox_Instance_1_L7}), .c ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .a ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}), .b ({new_AGEMA_signal_1999, LED_128_Instance_SBox_Instance_1_T1}), .c ({new_AGEMA_signal_2031, LED_128_Instance_SBox_Instance_1_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .a ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_2031, LED_128_Instance_SBox_Instance_1_L8}), .c ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .a ({new_AGEMA_signal_1807, LED_128_Instance_SBox_Instance_1_L4}), .b ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2073, LED_128_Instance_subcells_out[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .a ({new_AGEMA_signal_1936, LED_128_Instance_SBox_Instance_2_Q2}), .b ({new_AGEMA_signal_1810, LED_128_Instance_SBox_Instance_2_Q3}), .clk (CLK), .r (Fresh[36]), .c ({new_AGEMA_signal_1969, LED_128_Instance_SBox_Instance_2_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .a ({new_AGEMA_signal_1968, LED_128_Instance_SBox_Instance_2_Q6}), .b ({new_AGEMA_signal_1811, LED_128_Instance_SBox_Instance_2_Q7}), .clk (CLK), .r (Fresh[37]), .c ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .a ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}), .b ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2032, LED_128_Instance_SBox_Instance_2_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .a ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .b ({new_AGEMA_signal_2032, LED_128_Instance_SBox_Instance_2_L7}), .c ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .a ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}), .b ({new_AGEMA_signal_1969, LED_128_Instance_SBox_Instance_2_T1}), .c ({new_AGEMA_signal_2001, LED_128_Instance_SBox_Instance_2_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .a ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_2001, LED_128_Instance_SBox_Instance_2_L8}), .c ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .a ({new_AGEMA_signal_1751, LED_128_Instance_SBox_Instance_2_L4}), .b ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2034, LED_128_Instance_subcells_out[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .a ({new_AGEMA_signal_1938, LED_128_Instance_SBox_Instance_3_Q2}), .b ({new_AGEMA_signal_1815, LED_128_Instance_SBox_Instance_3_Q3}), .clk (CLK), .r (Fresh[38]), .c ({new_AGEMA_signal_1971, LED_128_Instance_SBox_Instance_3_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .a ({new_AGEMA_signal_1970, LED_128_Instance_SBox_Instance_3_Q6}), .b ({new_AGEMA_signal_1816, LED_128_Instance_SBox_Instance_3_Q7}), .clk (CLK), .r (Fresh[39]), .c ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .a ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}), .b ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2035, LED_128_Instance_SBox_Instance_3_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .a ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .b ({new_AGEMA_signal_2035, LED_128_Instance_SBox_Instance_3_L7}), .c ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .a ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}), .b ({new_AGEMA_signal_1971, LED_128_Instance_SBox_Instance_3_T1}), .c ({new_AGEMA_signal_2003, LED_128_Instance_SBox_Instance_3_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .a ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_2003, LED_128_Instance_SBox_Instance_3_L8}), .c ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .a ({new_AGEMA_signal_1757, LED_128_Instance_SBox_Instance_3_L4}), .b ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2037, LED_128_Instance_subcells_out[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .a ({new_AGEMA_signal_1972, LED_128_Instance_SBox_Instance_4_Q2}), .b ({new_AGEMA_signal_1892, LED_128_Instance_SBox_Instance_4_Q3}), .clk (CLK), .r (Fresh[40]), .c ({new_AGEMA_signal_2005, LED_128_Instance_SBox_Instance_4_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .a ({new_AGEMA_signal_2004, LED_128_Instance_SBox_Instance_4_Q6}), .b ({new_AGEMA_signal_1893, LED_128_Instance_SBox_Instance_4_Q7}), .clk (CLK), .r (Fresh[41]), .c ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .a ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}), .b ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2076, LED_128_Instance_SBox_Instance_4_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .a ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}), .b ({new_AGEMA_signal_2076, LED_128_Instance_SBox_Instance_4_L7}), .c ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .a ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}), .b ({new_AGEMA_signal_2005, LED_128_Instance_SBox_Instance_4_T1}), .c ({new_AGEMA_signal_2039, LED_128_Instance_SBox_Instance_4_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .a ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_2039, LED_128_Instance_SBox_Instance_4_L8}), .c ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .a ({new_AGEMA_signal_1821, LED_128_Instance_SBox_Instance_4_L4}), .b ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .a ({new_AGEMA_signal_1974, LED_128_Instance_SBox_Instance_5_Q2}), .b ({new_AGEMA_signal_1897, LED_128_Instance_SBox_Instance_5_Q3}), .clk (CLK), .r (Fresh[42]), .c ({new_AGEMA_signal_2007, LED_128_Instance_SBox_Instance_5_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .a ({new_AGEMA_signal_2006, LED_128_Instance_SBox_Instance_5_Q6}), .b ({new_AGEMA_signal_1898, LED_128_Instance_SBox_Instance_5_Q7}), .clk (CLK), .r (Fresh[43]), .c ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .a ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}), .b ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2079, LED_128_Instance_SBox_Instance_5_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .a ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}), .b ({new_AGEMA_signal_2079, LED_128_Instance_SBox_Instance_5_L7}), .c ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .a ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}), .b ({new_AGEMA_signal_2007, LED_128_Instance_SBox_Instance_5_T1}), .c ({new_AGEMA_signal_2041, LED_128_Instance_SBox_Instance_5_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .a ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_2041, LED_128_Instance_SBox_Instance_5_L8}), .c ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .a ({new_AGEMA_signal_1826, LED_128_Instance_SBox_Instance_5_L4}), .b ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .a ({new_AGEMA_signal_1944, LED_128_Instance_SBox_Instance_6_Q2}), .b ({new_AGEMA_signal_1829, LED_128_Instance_SBox_Instance_6_Q3}), .clk (CLK), .r (Fresh[44]), .c ({new_AGEMA_signal_1977, LED_128_Instance_SBox_Instance_6_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .a ({new_AGEMA_signal_1976, LED_128_Instance_SBox_Instance_6_Q6}), .b ({new_AGEMA_signal_1830, LED_128_Instance_SBox_Instance_6_Q7}), .clk (CLK), .r (Fresh[45]), .c ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .a ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}), .b ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2042, LED_128_Instance_SBox_Instance_6_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .a ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .b ({new_AGEMA_signal_2042, LED_128_Instance_SBox_Instance_6_L7}), .c ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .a ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}), .b ({new_AGEMA_signal_1977, LED_128_Instance_SBox_Instance_6_T1}), .c ({new_AGEMA_signal_2009, LED_128_Instance_SBox_Instance_6_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .a ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_2009, LED_128_Instance_SBox_Instance_6_L8}), .c ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .a ({new_AGEMA_signal_1764, LED_128_Instance_SBox_Instance_6_L4}), .b ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .a ({new_AGEMA_signal_1946, LED_128_Instance_SBox_Instance_7_Q2}), .b ({new_AGEMA_signal_1834, LED_128_Instance_SBox_Instance_7_Q3}), .clk (CLK), .r (Fresh[46]), .c ({new_AGEMA_signal_1979, LED_128_Instance_SBox_Instance_7_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .a ({new_AGEMA_signal_1978, LED_128_Instance_SBox_Instance_7_Q6}), .b ({new_AGEMA_signal_1835, LED_128_Instance_SBox_Instance_7_Q7}), .clk (CLK), .r (Fresh[47]), .c ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .a ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}), .b ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2045, LED_128_Instance_SBox_Instance_7_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .a ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .b ({new_AGEMA_signal_2045, LED_128_Instance_SBox_Instance_7_L7}), .c ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .a ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}), .b ({new_AGEMA_signal_1979, LED_128_Instance_SBox_Instance_7_T1}), .c ({new_AGEMA_signal_2011, LED_128_Instance_SBox_Instance_7_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .a ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_2011, LED_128_Instance_SBox_Instance_7_L8}), .c ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .a ({new_AGEMA_signal_1770, LED_128_Instance_SBox_Instance_7_L4}), .b ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .a ({new_AGEMA_signal_1980, LED_128_Instance_SBox_Instance_8_Q2}), .b ({new_AGEMA_signal_1906, LED_128_Instance_SBox_Instance_8_Q3}), .clk (CLK), .r (Fresh[48]), .c ({new_AGEMA_signal_2013, LED_128_Instance_SBox_Instance_8_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .a ({new_AGEMA_signal_2012, LED_128_Instance_SBox_Instance_8_Q6}), .b ({new_AGEMA_signal_1907, LED_128_Instance_SBox_Instance_8_Q7}), .clk (CLK), .r (Fresh[49]), .c ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .a ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}), .b ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2084, LED_128_Instance_SBox_Instance_8_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .a ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}), .b ({new_AGEMA_signal_2084, LED_128_Instance_SBox_Instance_8_L7}), .c ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .a ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}), .b ({new_AGEMA_signal_2013, LED_128_Instance_SBox_Instance_8_T1}), .c ({new_AGEMA_signal_2049, LED_128_Instance_SBox_Instance_8_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .a ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_2049, LED_128_Instance_SBox_Instance_8_L8}), .c ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .a ({new_AGEMA_signal_1840, LED_128_Instance_SBox_Instance_8_L4}), .b ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .a ({new_AGEMA_signal_1982, LED_128_Instance_SBox_Instance_9_Q2}), .b ({new_AGEMA_signal_1911, LED_128_Instance_SBox_Instance_9_Q3}), .clk (CLK), .r (Fresh[50]), .c ({new_AGEMA_signal_2015, LED_128_Instance_SBox_Instance_9_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .a ({new_AGEMA_signal_2014, LED_128_Instance_SBox_Instance_9_Q6}), .b ({new_AGEMA_signal_1912, LED_128_Instance_SBox_Instance_9_Q7}), .clk (CLK), .r (Fresh[51]), .c ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .a ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}), .b ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2087, LED_128_Instance_SBox_Instance_9_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .a ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}), .b ({new_AGEMA_signal_2087, LED_128_Instance_SBox_Instance_9_L7}), .c ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .a ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}), .b ({new_AGEMA_signal_2015, LED_128_Instance_SBox_Instance_9_T1}), .c ({new_AGEMA_signal_2051, LED_128_Instance_SBox_Instance_9_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .a ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_2051, LED_128_Instance_SBox_Instance_9_L8}), .c ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .a ({new_AGEMA_signal_1844, LED_128_Instance_SBox_Instance_9_L4}), .b ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .a ({new_AGEMA_signal_1952, LED_128_Instance_SBox_Instance_10_Q2}), .b ({new_AGEMA_signal_1847, LED_128_Instance_SBox_Instance_10_Q3}), .clk (CLK), .r (Fresh[52]), .c ({new_AGEMA_signal_1985, LED_128_Instance_SBox_Instance_10_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .a ({new_AGEMA_signal_1984, LED_128_Instance_SBox_Instance_10_Q6}), .b ({new_AGEMA_signal_1848, LED_128_Instance_SBox_Instance_10_Q7}), .clk (CLK), .r (Fresh[53]), .c ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .a ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}), .b ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2052, LED_128_Instance_SBox_Instance_10_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .a ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .b ({new_AGEMA_signal_2052, LED_128_Instance_SBox_Instance_10_L7}), .c ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .a ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}), .b ({new_AGEMA_signal_1985, LED_128_Instance_SBox_Instance_10_T1}), .c ({new_AGEMA_signal_2017, LED_128_Instance_SBox_Instance_10_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .a ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_2017, LED_128_Instance_SBox_Instance_10_L8}), .c ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .a ({new_AGEMA_signal_1779, LED_128_Instance_SBox_Instance_10_L4}), .b ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .a ({new_AGEMA_signal_1954, LED_128_Instance_SBox_Instance_11_Q2}), .b ({new_AGEMA_signal_1852, LED_128_Instance_SBox_Instance_11_Q3}), .clk (CLK), .r (Fresh[54]), .c ({new_AGEMA_signal_1987, LED_128_Instance_SBox_Instance_11_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .a ({new_AGEMA_signal_1986, LED_128_Instance_SBox_Instance_11_Q6}), .b ({new_AGEMA_signal_1853, LED_128_Instance_SBox_Instance_11_Q7}), .clk (CLK), .r (Fresh[55]), .c ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .a ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}), .b ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2055, LED_128_Instance_SBox_Instance_11_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .a ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .b ({new_AGEMA_signal_2055, LED_128_Instance_SBox_Instance_11_L7}), .c ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .a ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}), .b ({new_AGEMA_signal_1987, LED_128_Instance_SBox_Instance_11_T1}), .c ({new_AGEMA_signal_2019, LED_128_Instance_SBox_Instance_11_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .a ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_2019, LED_128_Instance_SBox_Instance_11_L8}), .c ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .a ({new_AGEMA_signal_1785, LED_128_Instance_SBox_Instance_11_L4}), .b ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .a ({new_AGEMA_signal_1988, LED_128_Instance_SBox_Instance_12_Q2}), .b ({new_AGEMA_signal_1920, LED_128_Instance_SBox_Instance_12_Q3}), .clk (CLK), .r (Fresh[56]), .c ({new_AGEMA_signal_2021, LED_128_Instance_SBox_Instance_12_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .a ({new_AGEMA_signal_2020, LED_128_Instance_SBox_Instance_12_Q6}), .b ({new_AGEMA_signal_1921, LED_128_Instance_SBox_Instance_12_Q7}), .clk (CLK), .r (Fresh[57]), .c ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .a ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}), .b ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2092, LED_128_Instance_SBox_Instance_12_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .a ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}), .b ({new_AGEMA_signal_2092, LED_128_Instance_SBox_Instance_12_L7}), .c ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .a ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}), .b ({new_AGEMA_signal_2021, LED_128_Instance_SBox_Instance_12_T1}), .c ({new_AGEMA_signal_2059, LED_128_Instance_SBox_Instance_12_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .a ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_2059, LED_128_Instance_SBox_Instance_12_L8}), .c ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .a ({new_AGEMA_signal_1860, LED_128_Instance_SBox_Instance_12_L4}), .b ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .a ({new_AGEMA_signal_1990, LED_128_Instance_SBox_Instance_13_Q2}), .b ({new_AGEMA_signal_1925, LED_128_Instance_SBox_Instance_13_Q3}), .clk (CLK), .r (Fresh[58]), .c ({new_AGEMA_signal_2023, LED_128_Instance_SBox_Instance_13_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .a ({new_AGEMA_signal_2022, LED_128_Instance_SBox_Instance_13_Q6}), .b ({new_AGEMA_signal_1926, LED_128_Instance_SBox_Instance_13_Q7}), .clk (CLK), .r (Fresh[59]), .c ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .a ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}), .b ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2095, LED_128_Instance_SBox_Instance_13_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .a ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}), .b ({new_AGEMA_signal_2095, LED_128_Instance_SBox_Instance_13_L7}), .c ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .a ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}), .b ({new_AGEMA_signal_2023, LED_128_Instance_SBox_Instance_13_T1}), .c ({new_AGEMA_signal_2061, LED_128_Instance_SBox_Instance_13_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .a ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_2061, LED_128_Instance_SBox_Instance_13_L8}), .c ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .a ({new_AGEMA_signal_1865, LED_128_Instance_SBox_Instance_13_L4}), .b ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .a ({new_AGEMA_signal_1960, LED_128_Instance_SBox_Instance_14_Q2}), .b ({new_AGEMA_signal_1868, LED_128_Instance_SBox_Instance_14_Q3}), .clk (CLK), .r (Fresh[60]), .c ({new_AGEMA_signal_1993, LED_128_Instance_SBox_Instance_14_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .a ({new_AGEMA_signal_1992, LED_128_Instance_SBox_Instance_14_Q6}), .b ({new_AGEMA_signal_1869, LED_128_Instance_SBox_Instance_14_Q7}), .clk (CLK), .r (Fresh[61]), .c ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .a ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}), .b ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2062, LED_128_Instance_SBox_Instance_14_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .a ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .b ({new_AGEMA_signal_2062, LED_128_Instance_SBox_Instance_14_L7}), .c ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .a ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}), .b ({new_AGEMA_signal_1993, LED_128_Instance_SBox_Instance_14_T1}), .c ({new_AGEMA_signal_2025, LED_128_Instance_SBox_Instance_14_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .a ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_2025, LED_128_Instance_SBox_Instance_14_L8}), .c ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .a ({new_AGEMA_signal_1792, LED_128_Instance_SBox_Instance_14_L4}), .b ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .a ({new_AGEMA_signal_1962, LED_128_Instance_SBox_Instance_15_Q2}), .b ({new_AGEMA_signal_1873, LED_128_Instance_SBox_Instance_15_Q3}), .clk (CLK), .r (Fresh[62]), .c ({new_AGEMA_signal_1995, LED_128_Instance_SBox_Instance_15_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .a ({new_AGEMA_signal_1994, LED_128_Instance_SBox_Instance_15_Q6}), .b ({new_AGEMA_signal_1874, LED_128_Instance_SBox_Instance_15_Q7}), .clk (CLK), .r (Fresh[63]), .c ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .a ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}), .b ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2065, LED_128_Instance_SBox_Instance_15_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .a ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .b ({new_AGEMA_signal_2065, LED_128_Instance_SBox_Instance_15_L7}), .c ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .a ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}), .b ({new_AGEMA_signal_1995, LED_128_Instance_SBox_Instance_15_T1}), .c ({new_AGEMA_signal_2027, LED_128_Instance_SBox_Instance_15_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .a ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_2027, LED_128_Instance_SBox_Instance_15_L8}), .c ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .a ({new_AGEMA_signal_1798, LED_128_Instance_SBox_Instance_15_L4}), .b ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U54 ( .a ({new_AGEMA_signal_2383, LED_128_Instance_MCS_Instance_0_n38}), .b ({new_AGEMA_signal_2244, LED_128_Instance_MCS_Instance_0_n37}), .c ({new_AGEMA_signal_2426, LED_128_Instance_mixcolumns_out[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U53 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2244, LED_128_Instance_MCS_Instance_0_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U52 ( .a ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}), .b ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .c ({new_AGEMA_signal_2383, LED_128_Instance_MCS_Instance_0_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U51 ( .a ({new_AGEMA_signal_2202, LED_128_Instance_MCS_Instance_0_n36}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U50 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_2202, LED_128_Instance_MCS_Instance_0_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U49 ( .a ({new_AGEMA_signal_2335, LED_128_Instance_MCS_Instance_0_n33}), .b ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}), .c ({new_AGEMA_signal_2427, LED_128_Instance_mixcolumns_out[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U48 ( .a ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2335, LED_128_Instance_MCS_Instance_0_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U47 ( .a ({new_AGEMA_signal_2486, LED_128_Instance_MCS_Instance_0_n32}), .b ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_2500, LED_128_Instance_mixcolumns_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U46 ( .a ({new_AGEMA_signal_2476, LED_128_Instance_MCS_Instance_0_n30}), .b ({new_AGEMA_signal_2284, LED_128_Instance_MCS_Instance_0_n29}), .c ({new_AGEMA_signal_2486, LED_128_Instance_MCS_Instance_0_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U45 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .c ({new_AGEMA_signal_2284, LED_128_Instance_MCS_Instance_0_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U44 ( .a ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}), .b ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_2476, LED_128_Instance_MCS_Instance_0_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U43 ( .a ({new_AGEMA_signal_2285, LED_128_Instance_MCS_Instance_0_n27}), .b ({new_AGEMA_signal_2245, LED_128_Instance_MCS_Instance_0_n26}), .c ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U42 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .c ({new_AGEMA_signal_2245, LED_128_Instance_MCS_Instance_0_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U41 ( .a ({new_AGEMA_signal_1931, LED_128_Instance_subcells_out[60]}), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_2285, LED_128_Instance_MCS_Instance_0_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U40 ( .a ({new_AGEMA_signal_2477, LED_128_Instance_MCS_Instance_0_n25}), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_2487, LED_128_Instance_mixcolumns_out[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U39 ( .a ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .b ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_2477, LED_128_Instance_MCS_Instance_0_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U38 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}), .c ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U37 ( .a ({new_AGEMA_signal_2384, LED_128_Instance_MCS_Instance_0_n24}), .b ({new_AGEMA_signal_2115, LED_128_Instance_MCS_Instance_0_n23}), .c ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U36 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2115, LED_128_Instance_MCS_Instance_0_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U35 ( .a ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .b ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .c ({new_AGEMA_signal_2384, LED_128_Instance_MCS_Instance_0_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U34 ( .a ({new_AGEMA_signal_2286, LED_128_Instance_MCS_Instance_0_n22}), .b ({new_AGEMA_signal_2172, LED_128_Instance_MCS_Instance_0_n21}), .c ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U33 ( .a ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2172, LED_128_Instance_MCS_Instance_0_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U32 ( .a ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .b ({new_AGEMA_signal_1943, LED_128_Instance_subcells_out[20]}), .c ({new_AGEMA_signal_2286, LED_128_Instance_MCS_Instance_0_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U31 ( .a ({new_AGEMA_signal_2203, LED_128_Instance_MCS_Instance_0_n19}), .b ({new_AGEMA_signal_2116, LED_128_Instance_MCS_Instance_0_n18}), .c ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U30 ( .a ({new_AGEMA_signal_1915, LED_128_Instance_subcells_out[40]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2116, LED_128_Instance_MCS_Instance_0_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U29 ( .a ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_2203, LED_128_Instance_MCS_Instance_0_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U28 ( .a ({new_AGEMA_signal_2140, LED_128_Instance_MCS_Instance_0_n16}), .b ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}), .c ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U27 ( .a ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}), .b ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2140, LED_128_Instance_MCS_Instance_0_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U26 ( .a ({new_AGEMA_signal_2339, LED_128_Instance_MCS_Instance_0_n15}), .b ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U25 ( .a ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U24 ( .a ({new_AGEMA_signal_2287, LED_128_Instance_MCS_Instance_0_n14}), .b ({new_AGEMA_signal_2117, LED_128_Instance_MCS_Instance_0_n13}), .c ({new_AGEMA_signal_2339, LED_128_Instance_MCS_Instance_0_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U23 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2117, LED_128_Instance_MCS_Instance_0_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U22 ( .a ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2287, LED_128_Instance_MCS_Instance_0_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U21 ( .a ({new_AGEMA_signal_2118, LED_128_Instance_MCS_Instance_0_n11}), .b ({new_AGEMA_signal_2247, LED_128_Instance_MCS_Instance_0_n10}), .c ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U20 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .c ({new_AGEMA_signal_2247, LED_128_Instance_MCS_Instance_0_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U19 ( .a ({new_AGEMA_signal_1915, LED_128_Instance_subcells_out[40]}), .b ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}), .c ({new_AGEMA_signal_2118, LED_128_Instance_MCS_Instance_0_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U18 ( .a ({new_AGEMA_signal_2204, LED_128_Instance_MCS_Instance_0_n9}), .b ({new_AGEMA_signal_2119, LED_128_Instance_MCS_Instance_0_n8}), .c ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U17 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2119, LED_128_Instance_MCS_Instance_0_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U16 ( .a ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}), .c ({new_AGEMA_signal_2204, LED_128_Instance_MCS_Instance_0_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U15 ( .a ({new_AGEMA_signal_2100, LED_128_Instance_MCS_Instance_0_n7}), .b ({new_AGEMA_signal_2141, LED_128_Instance_MCS_Instance_0_n6}), .c ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U14 ( .a ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}), .b ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2141, LED_128_Instance_MCS_Instance_0_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U13 ( .a ({new_AGEMA_signal_1933, LED_128_Instance_subcells_out[0]}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2100, LED_128_Instance_MCS_Instance_0_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U12 ( .a ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2340, LED_128_Instance_mixcolumns_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U11 ( .a ({new_AGEMA_signal_2142, LED_128_Instance_MCS_Instance_0_n4}), .b ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}), .c ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U10 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U9 ( .a ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}), .b ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}), .c ({new_AGEMA_signal_2142, LED_128_Instance_MCS_Instance_0_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U8 ( .a ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}), .b ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U7 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_1931, LED_128_Instance_subcells_out[60]}), .c ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U6 ( .a ({new_AGEMA_signal_2123, LED_128_Instance_MCS_Instance_0_n3}), .b ({new_AGEMA_signal_2122, LED_128_Instance_MCS_Instance_0_n2}), .c ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U5 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2122, LED_128_Instance_MCS_Instance_0_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U4 ( .a ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}), .b ({new_AGEMA_signal_1943, LED_128_Instance_subcells_out[20]}), .c ({new_AGEMA_signal_2123, LED_128_Instance_MCS_Instance_0_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U3 ( .a ({new_AGEMA_signal_2175, LED_128_Instance_MCS_Instance_0_n1}), .b ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .c ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U2 ( .a ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2070, LED_128_Instance_subcells_out[1]}), .c ({new_AGEMA_signal_2175, LED_128_Instance_MCS_Instance_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_0_U1 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}), .c ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U54 ( .a ({new_AGEMA_signal_2386, LED_128_Instance_MCS_Instance_1_n38}), .b ({new_AGEMA_signal_2206, LED_128_Instance_MCS_Instance_1_n37}), .c ({new_AGEMA_signal_2429, LED_128_Instance_mixcolumns_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U53 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2206, LED_128_Instance_MCS_Instance_1_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U52 ( .a ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}), .b ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .c ({new_AGEMA_signal_2386, LED_128_Instance_MCS_Instance_1_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U51 ( .a ({new_AGEMA_signal_2207, LED_128_Instance_MCS_Instance_1_n36}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U50 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_2207, LED_128_Instance_MCS_Instance_1_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U49 ( .a ({new_AGEMA_signal_2291, LED_128_Instance_MCS_Instance_1_n33}), .b ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}), .c ({new_AGEMA_signal_2387, LED_128_Instance_mixcolumns_out[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U48 ( .a ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2291, LED_128_Instance_MCS_Instance_1_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U47 ( .a ({new_AGEMA_signal_2488, LED_128_Instance_MCS_Instance_1_n32}), .b ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_2501, LED_128_Instance_mixcolumns_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U46 ( .a ({new_AGEMA_signal_2478, LED_128_Instance_MCS_Instance_1_n30}), .b ({new_AGEMA_signal_2292, LED_128_Instance_MCS_Instance_1_n29}), .c ({new_AGEMA_signal_2488, LED_128_Instance_MCS_Instance_1_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U45 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .c ({new_AGEMA_signal_2292, LED_128_Instance_MCS_Instance_1_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U44 ( .a ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}), .b ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_2478, LED_128_Instance_MCS_Instance_1_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U43 ( .a ({new_AGEMA_signal_2293, LED_128_Instance_MCS_Instance_1_n27}), .b ({new_AGEMA_signal_2208, LED_128_Instance_MCS_Instance_1_n26}), .c ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U42 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .c ({new_AGEMA_signal_2208, LED_128_Instance_MCS_Instance_1_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U41 ( .a ({new_AGEMA_signal_1957, LED_128_Instance_subcells_out[48]}), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_2293, LED_128_Instance_MCS_Instance_1_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U40 ( .a ({new_AGEMA_signal_2479, LED_128_Instance_MCS_Instance_1_n25}), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_2489, LED_128_Instance_mixcolumns_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U39 ( .a ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .b ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_2479, LED_128_Instance_MCS_Instance_1_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U38 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}), .c ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U37 ( .a ({new_AGEMA_signal_2388, LED_128_Instance_MCS_Instance_1_n24}), .b ({new_AGEMA_signal_2145, LED_128_Instance_MCS_Instance_1_n23}), .c ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U36 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2145, LED_128_Instance_MCS_Instance_1_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U35 ( .a ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .b ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .c ({new_AGEMA_signal_2388, LED_128_Instance_MCS_Instance_1_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U34 ( .a ({new_AGEMA_signal_2294, LED_128_Instance_MCS_Instance_1_n22}), .b ({new_AGEMA_signal_2146, LED_128_Instance_MCS_Instance_1_n21}), .c ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U33 ( .a ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2146, LED_128_Instance_MCS_Instance_1_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U32 ( .a ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .b ({new_AGEMA_signal_1901, LED_128_Instance_subcells_out[24]}), .c ({new_AGEMA_signal_2294, LED_128_Instance_MCS_Instance_1_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U31 ( .a ({new_AGEMA_signal_2209, LED_128_Instance_MCS_Instance_1_n19}), .b ({new_AGEMA_signal_2124, LED_128_Instance_MCS_Instance_1_n18}), .c ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U30 ( .a ({new_AGEMA_signal_1917, LED_128_Instance_subcells_out[44]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2124, LED_128_Instance_MCS_Instance_1_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U29 ( .a ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_2209, LED_128_Instance_MCS_Instance_1_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U28 ( .a ({new_AGEMA_signal_2147, LED_128_Instance_MCS_Instance_1_n16}), .b ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}), .c ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U27 ( .a ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}), .b ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2147, LED_128_Instance_MCS_Instance_1_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U26 ( .a ({new_AGEMA_signal_2296, LED_128_Instance_MCS_Instance_1_n15}), .b ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U25 ( .a ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U24 ( .a ({new_AGEMA_signal_2251, LED_128_Instance_MCS_Instance_1_n14}), .b ({new_AGEMA_signal_2125, LED_128_Instance_MCS_Instance_1_n13}), .c ({new_AGEMA_signal_2296, LED_128_Instance_MCS_Instance_1_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U23 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2125, LED_128_Instance_MCS_Instance_1_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U22 ( .a ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2251, LED_128_Instance_MCS_Instance_1_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U21 ( .a ({new_AGEMA_signal_2101, LED_128_Instance_MCS_Instance_1_n11}), .b ({new_AGEMA_signal_2210, LED_128_Instance_MCS_Instance_1_n10}), .c ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U20 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .c ({new_AGEMA_signal_2210, LED_128_Instance_MCS_Instance_1_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U19 ( .a ({new_AGEMA_signal_1917, LED_128_Instance_subcells_out[44]}), .b ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}), .c ({new_AGEMA_signal_2101, LED_128_Instance_MCS_Instance_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U18 ( .a ({new_AGEMA_signal_2211, LED_128_Instance_MCS_Instance_1_n9}), .b ({new_AGEMA_signal_2126, LED_128_Instance_MCS_Instance_1_n8}), .c ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U17 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2126, LED_128_Instance_MCS_Instance_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U16 ( .a ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}), .c ({new_AGEMA_signal_2211, LED_128_Instance_MCS_Instance_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U15 ( .a ({new_AGEMA_signal_2127, LED_128_Instance_MCS_Instance_1_n7}), .b ({new_AGEMA_signal_2148, LED_128_Instance_MCS_Instance_1_n6}), .c ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U14 ( .a ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}), .b ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2148, LED_128_Instance_MCS_Instance_1_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U13 ( .a ({new_AGEMA_signal_1935, LED_128_Instance_subcells_out[4]}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2127, LED_128_Instance_MCS_Instance_1_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U12 ( .a ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2297, LED_128_Instance_mixcolumns_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U11 ( .a ({new_AGEMA_signal_2128, LED_128_Instance_MCS_Instance_1_n4}), .b ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}), .c ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U10 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U9 ( .a ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}), .b ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}), .c ({new_AGEMA_signal_2128, LED_128_Instance_MCS_Instance_1_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U8 ( .a ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}), .b ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U7 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_1957, LED_128_Instance_subcells_out[48]}), .c ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U6 ( .a ({new_AGEMA_signal_2129, LED_128_Instance_MCS_Instance_1_n3}), .b ({new_AGEMA_signal_2150, LED_128_Instance_MCS_Instance_1_n2}), .c ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U5 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2150, LED_128_Instance_MCS_Instance_1_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U4 ( .a ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}), .b ({new_AGEMA_signal_1901, LED_128_Instance_subcells_out[24]}), .c ({new_AGEMA_signal_2129, LED_128_Instance_MCS_Instance_1_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U3 ( .a ({new_AGEMA_signal_2151, LED_128_Instance_MCS_Instance_1_n1}), .b ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .c ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U2 ( .a ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2073, LED_128_Instance_subcells_out[5]}), .c ({new_AGEMA_signal_2151, LED_128_Instance_MCS_Instance_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_1_U1 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}), .c ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U54 ( .a ({new_AGEMA_signal_2344, LED_128_Instance_MCS_Instance_2_n38}), .b ({new_AGEMA_signal_2213, LED_128_Instance_MCS_Instance_2_n37}), .c ({new_AGEMA_signal_2389, LED_128_Instance_mixcolumns_out[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U53 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2213, LED_128_Instance_MCS_Instance_2_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U52 ( .a ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}), .b ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .c ({new_AGEMA_signal_2344, LED_128_Instance_MCS_Instance_2_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U51 ( .a ({new_AGEMA_signal_2180, LED_128_Instance_MCS_Instance_2_n36}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U50 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_2180, LED_128_Instance_MCS_Instance_2_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U49 ( .a ({new_AGEMA_signal_2299, LED_128_Instance_MCS_Instance_2_n33}), .b ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}), .c ({new_AGEMA_signal_2390, LED_128_Instance_mixcolumns_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U48 ( .a ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2299, LED_128_Instance_MCS_Instance_2_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U47 ( .a ({new_AGEMA_signal_2480, LED_128_Instance_MCS_Instance_2_n32}), .b ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_2490, LED_128_Instance_mixcolumns_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U46 ( .a ({new_AGEMA_signal_2458, LED_128_Instance_MCS_Instance_2_n30}), .b ({new_AGEMA_signal_2255, LED_128_Instance_MCS_Instance_2_n29}), .c ({new_AGEMA_signal_2480, LED_128_Instance_MCS_Instance_2_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U45 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .c ({new_AGEMA_signal_2255, LED_128_Instance_MCS_Instance_2_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U44 ( .a ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}), .b ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_2458, LED_128_Instance_MCS_Instance_2_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U43 ( .a ({new_AGEMA_signal_2300, LED_128_Instance_MCS_Instance_2_n27}), .b ({new_AGEMA_signal_2214, LED_128_Instance_MCS_Instance_2_n26}), .c ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U42 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .c ({new_AGEMA_signal_2214, LED_128_Instance_MCS_Instance_2_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U41 ( .a ({new_AGEMA_signal_1959, LED_128_Instance_subcells_out[52]}), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_2300, LED_128_Instance_MCS_Instance_2_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U40 ( .a ({new_AGEMA_signal_2459, LED_128_Instance_MCS_Instance_2_n25}), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_2481, LED_128_Instance_mixcolumns_out[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U39 ( .a ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .b ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_2459, LED_128_Instance_MCS_Instance_2_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U38 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}), .c ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U37 ( .a ({new_AGEMA_signal_2346, LED_128_Instance_MCS_Instance_2_n24}), .b ({new_AGEMA_signal_2152, LED_128_Instance_MCS_Instance_2_n23}), .c ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U36 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2152, LED_128_Instance_MCS_Instance_2_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U35 ( .a ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .b ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .c ({new_AGEMA_signal_2346, LED_128_Instance_MCS_Instance_2_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U34 ( .a ({new_AGEMA_signal_2256, LED_128_Instance_MCS_Instance_2_n22}), .b ({new_AGEMA_signal_2153, LED_128_Instance_MCS_Instance_2_n21}), .c ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U33 ( .a ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2153, LED_128_Instance_MCS_Instance_2_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U32 ( .a ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .b ({new_AGEMA_signal_1903, LED_128_Instance_subcells_out[28]}), .c ({new_AGEMA_signal_2256, LED_128_Instance_MCS_Instance_2_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U31 ( .a ({new_AGEMA_signal_2181, LED_128_Instance_MCS_Instance_2_n19}), .b ({new_AGEMA_signal_2154, LED_128_Instance_MCS_Instance_2_n18}), .c ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U30 ( .a ({new_AGEMA_signal_1949, LED_128_Instance_subcells_out[32]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2154, LED_128_Instance_MCS_Instance_2_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U29 ( .a ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_2181, LED_128_Instance_MCS_Instance_2_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U28 ( .a ({new_AGEMA_signal_2131, LED_128_Instance_MCS_Instance_2_n16}), .b ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}), .c ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U27 ( .a ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}), .b ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2131, LED_128_Instance_MCS_Instance_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U26 ( .a ({new_AGEMA_signal_2303, LED_128_Instance_MCS_Instance_2_n15}), .b ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U25 ( .a ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U24 ( .a ({new_AGEMA_signal_2257, LED_128_Instance_MCS_Instance_2_n14}), .b ({new_AGEMA_signal_2156, LED_128_Instance_MCS_Instance_2_n13}), .c ({new_AGEMA_signal_2303, LED_128_Instance_MCS_Instance_2_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U23 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2156, LED_128_Instance_MCS_Instance_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U22 ( .a ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2257, LED_128_Instance_MCS_Instance_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U21 ( .a ({new_AGEMA_signal_2103, LED_128_Instance_MCS_Instance_2_n11}), .b ({new_AGEMA_signal_2216, LED_128_Instance_MCS_Instance_2_n10}), .c ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U20 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .c ({new_AGEMA_signal_2216, LED_128_Instance_MCS_Instance_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U19 ( .a ({new_AGEMA_signal_1949, LED_128_Instance_subcells_out[32]}), .b ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}), .c ({new_AGEMA_signal_2103, LED_128_Instance_MCS_Instance_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U18 ( .a ({new_AGEMA_signal_2217, LED_128_Instance_MCS_Instance_2_n9}), .b ({new_AGEMA_signal_2157, LED_128_Instance_MCS_Instance_2_n8}), .c ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U17 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2157, LED_128_Instance_MCS_Instance_2_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U16 ( .a ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}), .c ({new_AGEMA_signal_2217, LED_128_Instance_MCS_Instance_2_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U15 ( .a ({new_AGEMA_signal_2132, LED_128_Instance_MCS_Instance_2_n7}), .b ({new_AGEMA_signal_2158, LED_128_Instance_MCS_Instance_2_n6}), .c ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U14 ( .a ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}), .b ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2158, LED_128_Instance_MCS_Instance_2_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U13 ( .a ({new_AGEMA_signal_1887, LED_128_Instance_subcells_out[8]}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2132, LED_128_Instance_MCS_Instance_2_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U12 ( .a ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2304, LED_128_Instance_mixcolumns_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U11 ( .a ({new_AGEMA_signal_2159, LED_128_Instance_MCS_Instance_2_n4}), .b ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}), .c ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U10 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U9 ( .a ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}), .b ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}), .c ({new_AGEMA_signal_2159, LED_128_Instance_MCS_Instance_2_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U8 ( .a ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}), .b ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U7 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_1959, LED_128_Instance_subcells_out[52]}), .c ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U6 ( .a ({new_AGEMA_signal_2104, LED_128_Instance_MCS_Instance_2_n3}), .b ({new_AGEMA_signal_2161, LED_128_Instance_MCS_Instance_2_n2}), .c ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U5 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2161, LED_128_Instance_MCS_Instance_2_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U4 ( .a ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}), .b ({new_AGEMA_signal_1903, LED_128_Instance_subcells_out[28]}), .c ({new_AGEMA_signal_2104, LED_128_Instance_MCS_Instance_2_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U3 ( .a ({new_AGEMA_signal_2162, LED_128_Instance_MCS_Instance_2_n1}), .b ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .c ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U2 ( .a ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2034, LED_128_Instance_subcells_out[9]}), .c ({new_AGEMA_signal_2162, LED_128_Instance_MCS_Instance_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_2_U1 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}), .c ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U54 ( .a ({new_AGEMA_signal_2392, LED_128_Instance_MCS_Instance_3_n38}), .b ({new_AGEMA_signal_2261, LED_128_Instance_MCS_Instance_3_n37}), .c ({new_AGEMA_signal_2432, LED_128_Instance_mixcolumns_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U53 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2261, LED_128_Instance_MCS_Instance_3_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U52 ( .a ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}), .b ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .c ({new_AGEMA_signal_2392, LED_128_Instance_MCS_Instance_3_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U51 ( .a ({new_AGEMA_signal_2185, LED_128_Instance_MCS_Instance_3_n36}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U50 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_2185, LED_128_Instance_MCS_Instance_3_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U49 ( .a ({new_AGEMA_signal_2349, LED_128_Instance_MCS_Instance_3_n33}), .b ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}), .c ({new_AGEMA_signal_2433, LED_128_Instance_mixcolumns_out[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U48 ( .a ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2349, LED_128_Instance_MCS_Instance_3_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U47 ( .a ({new_AGEMA_signal_2482, LED_128_Instance_MCS_Instance_3_n32}), .b ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_2491, LED_128_Instance_mixcolumns_out[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U46 ( .a ({new_AGEMA_signal_2460, LED_128_Instance_MCS_Instance_3_n30}), .b ({new_AGEMA_signal_2262, LED_128_Instance_MCS_Instance_3_n29}), .c ({new_AGEMA_signal_2482, LED_128_Instance_MCS_Instance_3_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U45 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .c ({new_AGEMA_signal_2262, LED_128_Instance_MCS_Instance_3_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U44 ( .a ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}), .b ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_2460, LED_128_Instance_MCS_Instance_3_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U43 ( .a ({new_AGEMA_signal_2305, LED_128_Instance_MCS_Instance_3_n27}), .b ({new_AGEMA_signal_2263, LED_128_Instance_MCS_Instance_3_n26}), .c ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U42 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .c ({new_AGEMA_signal_2263, LED_128_Instance_MCS_Instance_3_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U41 ( .a ({new_AGEMA_signal_1929, LED_128_Instance_subcells_out[56]}), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_2305, LED_128_Instance_MCS_Instance_3_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U40 ( .a ({new_AGEMA_signal_2461, LED_128_Instance_MCS_Instance_3_n25}), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_2483, LED_128_Instance_mixcolumns_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U39 ( .a ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .b ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_2461, LED_128_Instance_MCS_Instance_3_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U38 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}), .c ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U37 ( .a ({new_AGEMA_signal_2351, LED_128_Instance_MCS_Instance_3_n24}), .b ({new_AGEMA_signal_2135, LED_128_Instance_MCS_Instance_3_n23}), .c ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U36 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2135, LED_128_Instance_MCS_Instance_3_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U35 ( .a ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .b ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .c ({new_AGEMA_signal_2351, LED_128_Instance_MCS_Instance_3_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U34 ( .a ({new_AGEMA_signal_2264, LED_128_Instance_MCS_Instance_3_n22}), .b ({new_AGEMA_signal_2186, LED_128_Instance_MCS_Instance_3_n21}), .c ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U33 ( .a ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2186, LED_128_Instance_MCS_Instance_3_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U32 ( .a ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .b ({new_AGEMA_signal_1941, LED_128_Instance_subcells_out[16]}), .c ({new_AGEMA_signal_2264, LED_128_Instance_MCS_Instance_3_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U31 ( .a ({new_AGEMA_signal_2187, LED_128_Instance_MCS_Instance_3_n19}), .b ({new_AGEMA_signal_2163, LED_128_Instance_MCS_Instance_3_n18}), .c ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U30 ( .a ({new_AGEMA_signal_1951, LED_128_Instance_subcells_out[36]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2163, LED_128_Instance_MCS_Instance_3_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U29 ( .a ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_2187, LED_128_Instance_MCS_Instance_3_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U28 ( .a ({new_AGEMA_signal_2136, LED_128_Instance_MCS_Instance_3_n16}), .b ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}), .c ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U27 ( .a ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}), .b ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2136, LED_128_Instance_MCS_Instance_3_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U26 ( .a ({new_AGEMA_signal_2353, LED_128_Instance_MCS_Instance_3_n15}), .b ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U25 ( .a ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U24 ( .a ({new_AGEMA_signal_2307, LED_128_Instance_MCS_Instance_3_n14}), .b ({new_AGEMA_signal_2165, LED_128_Instance_MCS_Instance_3_n13}), .c ({new_AGEMA_signal_2353, LED_128_Instance_MCS_Instance_3_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U23 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2165, LED_128_Instance_MCS_Instance_3_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U22 ( .a ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2307, LED_128_Instance_MCS_Instance_3_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U21 ( .a ({new_AGEMA_signal_2137, LED_128_Instance_MCS_Instance_3_n11}), .b ({new_AGEMA_signal_2265, LED_128_Instance_MCS_Instance_3_n10}), .c ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U20 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .c ({new_AGEMA_signal_2265, LED_128_Instance_MCS_Instance_3_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U19 ( .a ({new_AGEMA_signal_1951, LED_128_Instance_subcells_out[36]}), .b ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}), .c ({new_AGEMA_signal_2137, LED_128_Instance_MCS_Instance_3_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U18 ( .a ({new_AGEMA_signal_2220, LED_128_Instance_MCS_Instance_3_n9}), .b ({new_AGEMA_signal_2166, LED_128_Instance_MCS_Instance_3_n8}), .c ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U17 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2166, LED_128_Instance_MCS_Instance_3_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U16 ( .a ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}), .c ({new_AGEMA_signal_2220, LED_128_Instance_MCS_Instance_3_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U15 ( .a ({new_AGEMA_signal_2105, LED_128_Instance_MCS_Instance_3_n7}), .b ({new_AGEMA_signal_2167, LED_128_Instance_MCS_Instance_3_n6}), .c ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U14 ( .a ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}), .b ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2167, LED_128_Instance_MCS_Instance_3_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U13 ( .a ({new_AGEMA_signal_1889, LED_128_Instance_subcells_out[12]}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2105, LED_128_Instance_MCS_Instance_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U12 ( .a ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2354, LED_128_Instance_mixcolumns_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U11 ( .a ({new_AGEMA_signal_2168, LED_128_Instance_MCS_Instance_3_n4}), .b ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}), .c ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U10 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U9 ( .a ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}), .b ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}), .c ({new_AGEMA_signal_2168, LED_128_Instance_MCS_Instance_3_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U8 ( .a ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}), .b ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U7 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_1929, LED_128_Instance_subcells_out[56]}), .c ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U6 ( .a ({new_AGEMA_signal_2106, LED_128_Instance_MCS_Instance_3_n3}), .b ({new_AGEMA_signal_2169, LED_128_Instance_MCS_Instance_3_n2}), .c ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U5 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2169, LED_128_Instance_MCS_Instance_3_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U4 ( .a ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}), .b ({new_AGEMA_signal_1941, LED_128_Instance_subcells_out[16]}), .c ({new_AGEMA_signal_2106, LED_128_Instance_MCS_Instance_3_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U3 ( .a ({new_AGEMA_signal_2190, LED_128_Instance_MCS_Instance_3_n1}), .b ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .c ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U2 ( .a ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2037, LED_128_Instance_subcells_out[13]}), .c ({new_AGEMA_signal_2190, LED_128_Instance_MCS_Instance_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) LED_128_Instance_MCS_Instance_3_U1 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}), .c ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}) ) ;

    /* register cells */
    DFF_X1 LED_128_Instance_ks_reg_0__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N10), .Q (LED_128_Instance_ks_reg_0__Q), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_1__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N11), .Q (LED_128_Instance_n26), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_2__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N12), .Q (LED_128_Instance_n25), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_3__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N13), .Q (LED_128_Instance_n2), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_0__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N4), .Q (roundconstant[0]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_1__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N5), .Q (roundconstant[1]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_2__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N6), .Q (roundconstant[2]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_3__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N7), .Q (roundconstant[3]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_4__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N8), .Q (roundconstant[4]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_5__FF_FF ( .CK (clk_gated), .D (LED_128_Instance_N9), .Q (roundconstant[5]), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2201, LED_128_Instance_state1[0]}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2319, LED_128_Instance_state1[1]}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2227, LED_128_Instance_state1[2]}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2277, LED_128_Instance_state1[3]}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2229, LED_128_Instance_state1[4]}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2321, LED_128_Instance_state1[5]}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2231, LED_128_Instance_state1[6]}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2233, LED_128_Instance_state1[7]}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2235, LED_128_Instance_state1[8]}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2279, LED_128_Instance_state1[9]}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2237, LED_128_Instance_state1[10]}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2239, LED_128_Instance_state1[11]}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2241, LED_128_Instance_state1[12]}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2281, LED_128_Instance_state1[13]}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2243, LED_128_Instance_state1[14]}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2283, LED_128_Instance_state1[15]}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2368, LED_128_Instance_state1[16]}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2403, LED_128_Instance_state1[17]}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2405, LED_128_Instance_state1[18]}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2323, LED_128_Instance_state1[19]}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2325, LED_128_Instance_state1[20]}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2370, LED_128_Instance_state1[21]}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2407, LED_128_Instance_state1[22]}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2327, LED_128_Instance_state1[23]}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2329, LED_128_Instance_state1[24]}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2372, LED_128_Instance_state1[25]}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2374, LED_128_Instance_state1[26]}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2331, LED_128_Instance_state1[27]}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2376, LED_128_Instance_state1[28]}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2409, LED_128_Instance_state1[29]}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2378, LED_128_Instance_state1[30]}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2333, LED_128_Instance_state1[31]}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2411, LED_128_Instance_state1[32]}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2443, LED_128_Instance_state1[33]}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2413, LED_128_Instance_state1[34]}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2463, LED_128_Instance_state1[35]}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2415, LED_128_Instance_state1[36]}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2417, LED_128_Instance_state1[37]}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2380, LED_128_Instance_state1[38]}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2465, LED_128_Instance_state1[39]}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2419, LED_128_Instance_state1[40]}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2421, LED_128_Instance_state1[41]}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2382, LED_128_Instance_state1[42]}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2445, LED_128_Instance_state1[43]}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2423, LED_128_Instance_state1[44]}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2447, LED_128_Instance_state1[45]}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2425, LED_128_Instance_state1[46]}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2449, LED_128_Instance_state1[47]}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2505, LED_128_Instance_state1[48]}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2513, LED_128_Instance_state1[49]}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2467, LED_128_Instance_state1[50]}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2469, LED_128_Instance_state1[51]}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2507, LED_128_Instance_state1[52]}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2515, LED_128_Instance_state1[53]}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2451, LED_128_Instance_state1[54]}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2471, LED_128_Instance_state1[55]}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2497, LED_128_Instance_state1[56]}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2509, LED_128_Instance_state1[57]}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2453, LED_128_Instance_state1[58]}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2455, LED_128_Instance_state1[59]}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2499, LED_128_Instance_state1[60]}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2511, LED_128_Instance_state1[61]}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2473, LED_128_Instance_state1[62]}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) LED_128_Instance_cipherstate_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2475, LED_128_Instance_state1[63]}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 internal_done_reg_FF_FF ( .CK (clk_gated), .D (n15), .Q (OUT_done), .QN () ) ;
endmodule
