module PRESENT_Top(x, y);
 input [145:0] x;
 output [64:0] y;

 wire [1742:0] t;
  FX FX_inst(.x({t[614], t[613], t[612], t[611], t[610], t[609], t[608], t[607], t[606], t[605], t[604], t[603], t[602], t[601], t[600], t[599], t[598], t[597], t[596], t[595], t[594], t[593], t[592], t[591], t[590], t[589], t[588], t[587], t[586], t[585], t[584], t[583], t[582], t[581], t[580], t[579], t[578], t[577], t[576], t[575], t[574], t[573], t[572], t[571], t[570], t[569], t[568], t[567], t[566], t[565], t[564], t[563], t[562], t[561], t[560], t[559], t[558], t[557], t[556], t[555], t[554], t[553], t[552], t[551], t[550], t[549], t[548], t[547], t[546], t[545], t[544], t[543], t[542], t[541], t[540], t[539], t[538], t[537], t[536], t[535], t[534], t[533], t[532], t[531], t[530], t[529], t[528], t[527], t[526], t[525], t[524], t[523], t[522], t[521], t[520], t[519], t[518], t[517], t[516], t[515], t[514], t[513], t[512], t[511], t[510], t[509], t[508], t[507], t[506], t[505], t[504], t[503], t[502], t[501], t[500], t[499], t[498], t[497], t[496], t[495], t[494], t[493], t[492], t[491], t[490], t[489], t[488], t[487], t[486], t[485], t[484], t[483], t[482], t[481], t[480], t[479], t[478], t[477], t[476], t[475], t[474], t[473], t[472], t[471], t[470], t[469], t[468], t[467], t[466], t[465], t[464], t[463], t[462], t[461], t[460], t[459], t[458], t[457], t[456], t[455], t[454], t[453], t[452], t[451], t[450], t[449], t[448], t[447], t[446], t[445], t[444], t[443], t[442], t[441], t[440], t[439], t[438], t[437], t[436], t[435], t[434], t[433], t[432], t[431], t[430], t[429], t[428], t[427], t[426], t[425], t[424], t[423], t[422], t[421], t[420], t[419], t[418], t[417], t[416], t[415], t[414], t[413], t[412], t[411], t[410], t[409], t[408], t[407], t[406], t[405], t[404], t[403], t[402], t[401], t[400], t[399], t[398], t[397], t[396], t[395], t[394], t[393], t[392], t[391], t[390], t[389], t[388], t[387], t[386], t[385], t[384], t[383], t[382], t[381], t[380], t[379], t[378], t[377], t[376], t[375], t[374], t[373], t[372], t[371], t[370], t[369], t[368], t[367], t[366], t[365], t[364], t[363], t[362], t[361], t[360], t[359], t[358], t[357], t[356], t[355], t[354], t[353], t[352], t[351], t[350], t[349], t[348], t[347], t[346], t[345], t[344], t[343], t[342], t[341], t[340], t[339], t[338], t[337], t[336], t[335], t[334], t[333], t[332], t[331], t[330], t[329], t[328], t[327], t[326], t[325], t[324], t[323], t[322], t[321], t[320], t[319], t[318], t[317], t[316], t[315], t[314], t[313], t[312], t[311], t[310], t[309], t[308], t[307], t[306], t[305], t[304], t[303], t[302], t[301], t[300], t[299], t[298], t[297], t[296], t[295], t[294], t[293], t[292], t[291], t[290], t[289], t[288], t[287], t[286], t[285], t[284], t[283], t[282], t[281], t[280], t[279], t[278], t[277], t[276], t[275], t[274], t[273], t[272], t[271], t[270], t[269], t[268], t[267], t[266], t[265], t[264], t[263], t[262], t[261], t[260], t[259], t[258], t[257], t[256], t[255], t[254], t[253], t[252], t[251], t[250], t[249], t[248], t[247], t[246], t[245], t[244], t[243], t[242], t[241], t[240], t[239], t[238], t[237], t[236], t[235], t[234], t[233], t[232], t[231], t[230], t[229], t[228], t[227], t[226], t[225], t[224], t[223], t[222], t[221], t[220], t[219], t[218], t[217], t[216], t[215], t[214], t[213], t[212], t[211], t[210], t[209], t[208], t[207], t[206], t[205], t[204], t[203], t[202], t[201], t[200], t[199], t[198], t[197], t[196], t[195], t[194], t[193], t[192], t[191], t[190], t[189], t[188], t[187], t[186], t[185], t[184], t[183], t[182], t[181], t[180], t[179], t[178], t[177], t[176], t[175], t[174], t[173], t[172], t[171], t[170], t[169], t[168], t[167], t[166], t[165], t[164], t[163], t[162], t[161], t[160], t[159], t[158], t[157], t[156], t[155], t[154], t[153], t[152], t[151], t[150], t[149], t[148], t[147], t[146], t[145], t[144], t[143], t[142], t[141], t[140], t[139], t[138], t[137], t[136], t[135], t[134], t[133], t[132], t[131], t[130], t[129], t[128], t[127], t[126], t[125], t[124], t[123], t[122], t[121], t[120], t[119], t[118], t[117], t[116], t[115], t[114], t[113], t[112], t[111], t[110], t[109], t[108], t[107], t[106], t[105], t[104], t[103], t[102], t[101], t[100], t[99], t[98], t[97], t[96], t[95], t[94], t[93], t[92], t[91], t[90], t[89], t[88], t[87], t[86], t[85], t[84], t[83], t[82], t[81], t[80], t[79], t[78], t[77], t[76], t[75], t[74], t[73], t[72], t[71], t[70], t[69], t[68], t[67], t[66], t[65], t[64], t[63], t[62], t[61], t[60], t[59], t[58], t[57], t[56], t[55], t[54], t[53], t[52], t[51], t[50], t[49], t[48], t[47], t[46], t[45], t[44], t[43], t[42], t[41], t[40], t[39], t[38], t[37], t[36], t[35], t[34], t[33], t[32], t[31], t[30], t[29], t[28], t[27], t[26], t[25], t[24], t[23], t[22], t[21], t[20], t[19], t[18], t[17], t[16], t[15], t[14], t[13], t[12], t[11], t[10], t[9], t[8], t[7], t[6], t[5], t[4], t[3], t[2], t[1], t[0]}), .y({t[1055], t[1054], t[1053], t[1052], t[1051], t[1050], t[1049], t[1048], t[1047], t[1046], t[1045], t[1044], t[1043], t[1042], t[1041], t[1040], t[1039], t[1038], t[1037], t[1036], t[1035], t[1034], t[1033], t[1032], t[1031], t[1030], t[1029], t[1028], t[1027], t[1026], t[1025], t[1024], t[1023], t[1022], t[1021], t[1020], t[1019], t[1018], t[1017], t[1016], t[1015], t[1014], t[1013], t[1012], t[1011], t[1010], t[1009], t[1008], t[1007], t[1006], t[1005], t[1004], t[1003], t[1002], t[1001], t[1000], t[999], t[998], t[997], t[996], t[995], t[994], t[993], t[992], t[991], t[990], t[989], t[988], t[987], t[986], t[985], t[984], t[983], t[982], t[981], t[980], t[979], t[978], t[977], t[976], t[975], t[974], t[973], t[972], t[971], t[970], t[969], t[968], t[967], t[966], t[965], t[964], t[963], t[962], t[961], t[960], t[959], t[958], t[957], t[956], t[955], t[954], t[953], t[952], t[951], t[950], t[949], t[948], t[947], t[946], t[945], t[944], t[943], t[942], t[941], t[940], t[939], t[938], t[937], t[936], t[935], t[934], t[933], t[932], t[931], t[930], t[929], t[928], t[927], t[926], t[925], t[924], t[923], t[922], t[921], t[920], t[919], t[918], t[917], t[916], t[915], t[914], t[913], t[912], t[911], t[910], t[909], t[908], t[907], t[906], t[905], t[904], t[903], t[902], t[901], t[900], t[899], t[898], t[897], t[896], t[895], t[894], t[893], t[892], t[891], t[890], t[889], t[888], t[887], t[886], t[885], t[884], t[883], t[882], t[881], t[880], t[879], t[878], t[877], t[876], t[875], t[874], t[873], t[872], t[871], t[870], t[869], t[868], t[867], t[866], t[865], t[864], t[863], t[862], t[861], t[860], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[852], t[851], t[850], t[849], t[848], t[847], t[846], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[803], t[802], t[801], t[800], t[799], t[798], t[797], t[796], t[795], t[794], t[793], t[792], t[791], t[790], t[789], t[788], t[787], t[786], t[785], t[784], t[783], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[761], t[760], t[759], t[758], t[757], t[756], t[755], t[754], t[753], t[752], t[751], t[750], t[749], t[748], t[747], t[746], t[745], t[744], t[743], t[742], t[741], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[719], t[718], t[717], t[716], t[715], t[714], t[713], t[712], t[711], t[710], t[709], t[708], t[707], t[706], t[705], t[704], t[703], t[702], t[701], t[700], t[699], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[684], t[683], t[682], t[681], t[680], t[679], t[678], t[677], t[676], t[675], t[674], t[673], t[672], t[671], t[670], t[669], t[668], t[667], t[666], t[665], t[664], t[663], t[662], t[661], t[660], t[659], t[658], t[657], t[656], t[655], t[654], t[653], t[652], t[651], t[650], t[649], t[648], t[647], t[646], t[645], t[644], t[643], t[642], t[641], t[640], t[639], t[638], t[637], t[636], t[635], t[634], t[633], t[632], t[631], t[630], t[629], t[628], t[627], t[626], t[625], t[624], t[623], t[622], t[621], t[620], t[619], t[618], t[617], t[616], t[615]}));
  R1_ind R1_ind_inst(.x({t[136], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[168], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[144], t[747], t[746], t[745], t[744], t[743], t[742], t[741], x[60], x[61], x[62], x[63], x[56], x[57], x[58], x[59], x[52], x[53], x[54], x[55], x[48], x[49], x[50], x[51], x[44], x[45], x[46], x[47], x[40], x[41], x[42], x[43], x[36], x[37], x[38], x[39], x[32], x[33], x[34], x[35], x[28], x[29], x[30], x[31], t[152], t[754], t[753], t[752], t[751], t[750], t[749], t[748], x[24], x[25], x[26], x[27], x[20], x[21], x[22], x[23], x[16], x[17], x[18], x[19], x[12], x[13], x[14], x[15], x[8], x[9], x[10], x[11], x[4], x[5], x[6], x[7], x[0], x[1], x[2], x[3], t[128], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[160], t[761], t[760], t[759], t[758], t[757], t[756], t[755], x[140], x[141], x[142], x[143], x[136], t[318], x[137], t[319], x[138], t[320], x[139], t[322], t[873], t[872], t[871], t[870], t[869], t[868], t[867], x[132], t[329], x[133], t[330], x[134], t[331], x[135], t[333], t[880], t[879], t[878], t[877], t[876], t[875], t[874], t[64], t[677], t[676], t[675], t[674], t[673], t[672], t[671], x[128], t[340], x[129], t[341], x[130], t[342], x[131], t[344], t[887], t[886], t[885], t[884], t[883], t[882], t[881], t[40], t[656], t[655], t[654], t[653], t[652], t[651], t[650], x[124], t[351], t[72], t[684], t[683], t[682], t[681], t[680], t[679], t[678], x[125], t[352], t[48], t[663], t[662], t[661], t[660], t[659], t[658], t[657], x[126], t[353], t[56], t[670], t[669], t[668], t[667], t[666], t[665], t[664], x[127], t[355], t[894], t[893], t[892], t[891], t[890], t[889], t[888], x[120], t[362], x[121], t[363], x[122], t[364], x[123], t[120], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[366], t[901], t[900], t[899], t[898], t[897], t[896], t[895], x[116], t[373], x[117], t[374], x[118], t[375], x[119], t[377], t[908], t[907], t[906], t[905], t[904], t[903], t[902], x[112], t[384], x[113], t[385], x[114], t[386], x[115], t[388], t[915], t[914], t[913], t[912], t[911], t[910], t[909], x[108], t[395], x[109], t[396], x[110], t[397], x[111], t[399], t[922], t[921], t[920], t[919], t[918], t[917], t[916], x[104], t[406], x[105], t[407], x[106], t[408], x[107], t[410], t[929], t[928], t[927], t[926], t[925], t[924], t[923], x[100], t[417], x[101], t[418], x[102], t[419], x[103], t[421], t[936], t[935], t[934], t[933], t[932], t[931], t[930], x[96], t[494], x[97], t[495], x[98], t[496], x[99], t[192], t[789], t[788], t[787], t[786], t[785], t[784], t[783], t[498], t[985], t[984], t[983], t[982], t[981], t[980], t[979], x[92], t[505], x[93], t[506], x[94], t[507], x[95], t[184], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[509], t[992], t[991], t[990], t[989], t[988], t[987], t[986], x[88], t[516], x[89], t[517], x[90], t[518], x[91], t[520], t[999], t[998], t[997], t[996], t[995], t[994], t[993], x[84], t[527], x[85], t[528], x[86], t[529], x[87], t[531], t[1006], t[1005], t[1004], t[1003], t[1002], t[1001], t[1000], x[80], t[538], x[81], t[539], x[82], t[540], x[83], t[542], t[1013], t[1012], t[1011], t[1010], t[1009], t[1008], t[1007], x[76], t[549], x[77], t[550], x[78], t[551], x[79], t[553], t[1020], t[1019], t[1018], t[1017], t[1016], t[1015], t[1014], x[72], t[560], x[73], t[561], x[74], t[562], x[75], t[564], t[1027], t[1026], t[1025], t[1024], t[1023], t[1022], t[1021], x[68], t[571], x[69], t[572], x[70], t[573], x[71], t[575], t[1034], t[1033], t[1032], t[1031], t[1030], t[1029], t[1028], x[64], t[593], t[582], x[65], t[594], t[583], x[66], t[595], t[584], t[606], t[604], t[608], t[605], t[1055], t[1054], t[1053], t[1052], t[1051], t[1050], t[1049], x[67], x[145], t[200], t[796], t[795], t[794], t[793], t[792], t[791], t[790], t[176], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[597], t[1048], t[1047], t[1046], t[1045], t[1044], t[1043], t[1042], t[586], t[1041], t[1040], t[1039], t[1038], t[1037], t[1036], t[1035], t[96], t[705], t[704], t[703], t[702], t[701], t[700], t[699], t[104], t[712], t[711], t[710], t[709], t[708], t[707], t[706], t[88], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[80], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[24], t[642], t[641], t[640], t[639], t[638], t[637], t[636], t[32], t[649], t[648], t[647], t[646], t[645], t[644], t[643], t[16], t[635], t[634], t[633], t[632], t[631], t[630], t[629], t[8], t[628], t[627], t[626], t[625], t[624], t[623], t[622], t[112], t[719], t[718], t[717], t[716], t[715], t[714], t[713], t[487], t[485], t[484], t[483], t[978], t[977], t[976], t[975], t[974], t[973], t[972], t[476], t[474], t[473], t[472], t[971], t[970], t[969], t[968], t[967], t[966], t[965], t[465], t[463], t[462], t[461], t[964], t[963], t[962], t[961], t[960], t[959], t[958], t[454], t[452], t[451], t[450], t[957], t[956], t[955], t[954], t[953], t[952], t[951], t[443], t[441], t[440], t[439], t[950], t[949], t[948], t[947], t[946], t[945], t[944], t[432], t[430], t[429], t[428], t[943], t[942], t[941], t[940], t[939], t[938], t[937], t[311], t[309], t[308], t[307], t[866], t[865], t[864], t[863], t[862], t[861], t[860], t[300], t[298], t[297], t[296], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[289], t[287], t[286], t[285], t[852], t[851], t[850], t[849], t[848], t[847], t[846], t[278], t[276], t[275], t[274], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[267], t[265], t[264], t[263], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[256], t[254], t[253], t[252], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[245], t[243], t[242], t[241], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[234], t[232], t[231], t[230], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[223], t[221], t[220], t[219], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[212], t[210], t[209], t[208], t[803], t[802], t[801], t[800], t[799], t[798], t[797], t[0], t[621], t[620], t[619], t[618], t[617], t[616], t[615]}), .y({t[1294], t[1293], t[1292], t[1291], t[1290], t[1289], t[1288], t[1287], t[1286], t[1285], t[1284], t[1283], t[1282], t[1281], t[1280], t[1279], t[1278], t[1277], t[1276], t[1275], t[1274], t[1273], t[1272], t[1271], t[1270], t[1269], t[1268], t[1267], t[1266], t[1265], t[1264], t[1263], t[1262], t[1261], t[1260], t[1259], t[1258], t[1257], t[1256], t[1255], t[1254], t[1253], t[1252], t[1251], t[1250], t[1249], t[1248], t[1247], t[1246], t[1245], t[1244], t[1243], t[1242], t[1241], t[1240], t[1239], t[1238], t[1237], t[1236], t[1235], t[1234], t[1233], t[1232], t[1231], t[1230], t[1229], t[1228], t[1227], t[1226], t[1225], t[1224], t[1223], t[1222], t[1221], t[1220], t[1219], t[1218], t[1217], t[1216], t[1215], t[1214], t[1213], t[1212], t[1211], t[1210], t[1209], t[1208], t[1207], t[1206], t[1205], t[1204], t[1203], t[1202], t[1201], t[1200], t[1199], t[1198], t[1197], t[1196], t[1195], t[1194], t[1193], t[1192], t[1191], t[1190], t[1189], t[1188], t[1187], t[1186], t[1185], t[1184], t[1183], t[1182], t[1181], t[1180], t[1179], t[1178], t[1177], t[1176], t[1175], t[1174], t[1173], t[1172], t[1171], t[1170], t[1169], t[1168], t[1167], t[1166], t[1165], t[1164], t[1163], t[1162], t[1161], t[1160], t[1159], t[1158], t[1157], t[1156], t[1155], t[1154], t[1153], t[1152], t[1151], t[1150], t[1149], t[1148], t[1147], t[1146], t[1145], t[1144], t[1143], t[1142], t[1141], t[1140], t[1139], t[1138], t[1137], t[1136], t[1135], t[1134], t[1133], t[1132], t[1131], t[1130], t[1129], t[1128], t[1127], t[1126], t[1125], t[1124], t[1123], t[1122], t[1121], t[1120], t[1119], t[1118], t[1117], t[1116], t[1115], t[1114], t[1113], t[1112], t[1111], t[1110], t[1109], t[1108], t[1107], t[1106], t[1105], t[1104], t[1103], t[1102], t[1101], t[1100], t[1099], t[1098], t[1097], t[1096], t[1095], t[1094], t[1093], t[1092], t[1091], t[1090], t[1089], t[1088], t[1087], t[1086], t[1085], t[1084], t[1083], t[1082], t[1081], t[1080], t[1079], t[1078], t[1077], t[1076], t[1075], t[1074], t[1073], t[1072], t[1071], t[1070], t[1069], t[1068], t[1067], t[1066], t[1065], t[1064], t[1063], t[1062], t[1061], t[1060], t[1059], t[1058], t[1057], t[1056]}));
  R2_ind R2_ind_inst(.x({x[67], x[66], x[65], x[64], x[71], x[70], x[69], x[68], x[75], x[74], x[73], t[591], t[590], t[589], t[587], x[72], t[588], t[585], t[592], t[586], t[584], t[583], t[582], x[79], x[78], x[77], t[580], t[579], t[578], t[576], x[76], t[577], t[574], t[581], t[575], t[573], t[572], t[571], x[83], x[82], x[81], t[569], t[568], t[567], t[565], x[80], t[566], t[563], t[570], t[564], t[562], t[561], t[560], x[87], x[86], x[85], t[558], t[557], t[556], t[554], x[84], t[555], t[552], t[559], t[553], t[551], t[550], t[549], x[91], x[90], x[89], t[547], t[546], t[545], t[543], x[88], t[544], t[541], t[548], t[542], t[540], t[539], t[538], x[95], x[94], x[93], t[536], t[535], t[534], t[532], x[92], t[533], t[530], t[537], t[531], t[529], t[528], t[527], t[205], t[201], t[207], t[206], t[204], t[203], t[202], t[200], x[99], x[98], x[97], t[525], t[524], t[523], t[521], x[96], t[522], t[519], t[526], t[520], t[518], t[517], t[516], x[103], x[102], x[101], t[514], t[513], t[512], t[510], x[100], t[511], t[508], t[515], t[509], t[507], t[506], t[505], x[3], x[2], x[1], x[0], x[7], x[6], x[5], x[4], x[11], x[10], x[9], x[8], x[15], x[14], x[13], x[12], x[19], x[18], x[17], x[16], x[23], x[22], x[21], x[20], x[107], x[106], x[105], t[503], t[502], t[501], t[499], x[104], t[500], t[497], t[504], t[498], t[496], t[495], t[494], x[111], x[110], x[109], t[426], t[425], t[424], t[422], x[108], t[423], t[420], t[427], t[421], t[419], t[418], t[417], x[115], x[114], x[113], t[415], t[414], t[413], t[411], x[112], t[412], t[409], t[416], t[410], t[408], t[407], t[406], x[119], x[118], x[117], t[404], t[403], t[402], t[400], x[116], t[401], t[398], t[405], t[399], t[397], t[396], t[395], x[123], x[122], x[121], t[393], t[392], t[391], t[389], x[120], t[390], t[387], t[394], t[388], t[386], t[385], t[384], x[127], x[126], t[382], t[381], t[380], t[378], x[125], t[379], t[376], t[383], t[377], t[375], t[374], t[373], x[124], x[131], x[130], x[129], t[371], t[370], t[369], t[367], t[368], t[365], t[372], t[366], t[364], t[363], t[362], x[128], x[135], x[134], x[133], t[360], t[359], t[358], t[356], x[132], t[357], t[354], t[361], t[355], t[353], t[352], t[351], x[139], x[138], x[137], t[349], t[348], t[347], t[345], x[136], t[346], t[343], t[350], t[344], t[342], t[341], t[340], t[189], t[185], t[191], t[190], t[188], t[187], t[186], t[184], x[143], x[142], t[327], t[325], t[323], x[141], t[338], t[337], t[336], t[334], t[324], x[140], t[335], t[332], t[339], t[333], t[331], t[330], t[329], t[181], t[177], t[183], t[182], t[180], t[179], t[178], t[176], t[326], t[321], t[328], t[322], t[320], t[319], t[318], t[197], t[193], t[199], t[198], t[196], t[195], t[194], t[192], x[27], x[26], x[25], x[24], t[165], t[161], t[167], t[166], t[164], t[163], t[162], t[160], x[31], x[30], x[29], x[28], x[35], x[34], x[33], x[32], x[39], x[38], x[37], x[36], x[43], x[42], x[41], x[40], x[47], x[46], x[45], x[44], x[51], t[459], t[458], t[457], t[455], t[453], t[460], t[456], t[454], t[452], t[451], t[450], x[50], t[470], t[469], t[468], t[466], t[464], t[471], t[467], t[465], t[463], t[462], t[461], x[49], t[481], t[480], t[479], t[477], t[475], t[482], t[478], t[476], t[474], t[473], t[472], x[48], x[55], t[305], t[304], t[303], t[301], t[299], t[306], t[302], t[300], t[298], t[297], t[296], x[54], t[316], t[315], t[314], t[312], t[310], t[317], t[313], t[311], t[309], t[308], t[307], x[53], t[437], t[436], t[435], t[433], t[431], t[438], t[434], t[432], t[430], t[429], t[428], x[52], t[448], t[447], t[446], t[444], t[442], t[449], t[445], t[443], t[441], t[440], t[439], t[157], t[153], t[159], t[158], t[156], t[155], t[154], t[152], x[59], t[261], t[260], t[259], t[257], t[255], t[262], t[258], t[256], t[254], t[253], t[252], x[58], t[272], t[271], t[270], t[268], t[266], t[273], t[269], t[267], t[265], t[264], t[263], x[57], t[283], t[282], t[281], t[279], t[277], t[284], t[280], t[278], t[276], t[275], t[274], x[56], t[294], t[293], t[292], t[290], t[288], t[295], t[291], t[289], t[287], t[286], t[285], x[60], t[250], t[249], t[248], t[246], t[244], t[251], t[247], t[245], t[243], t[242], t[241], t[489], t[599], x[61], t[239], t[238], t[237], t[235], t[233], t[240], t[236], t[234], t[232], t[231], t[230], t[217], t[215], t[213], x[62], t[228], t[227], t[226], t[224], t[222], t[229], t[225], t[223], t[221], t[220], t[219], t[214], t[613], t[612], t[611], t[609], t[610], t[607], t[614], t[608], t[606], t[605], t[604], t[492], t[491], t[490], t[488], t[486], t[493], t[487], t[485], t[484], t[483], t[602], t[601], t[600], t[598], t[596], t[603], t[597], t[595], t[594], t[593], x[63], t[216], t[211], t[218], t[212], t[210], t[209], t[208], t[173], t[169], t[175], t[174], t[172], t[171], t[170], t[168], t[149], t[145], t[151], t[150], t[148], t[147], t[146], t[144], t[133], t[129], t[135], t[134], t[132], t[131], t[130], t[128], t[141], t[137], t[143], t[142], t[140], t[139], t[138], t[136], t[125], t[121], t[127], t[126], t[124], t[123], t[122], t[120], t[69], t[65], t[71], t[70], t[68], t[67], t[66], t[64], t[45], t[41], t[47], t[46], t[44], t[43], t[42], t[40], t[53], t[49], t[55], t[54], t[52], t[51], t[50], t[48], t[77], t[73], t[79], t[78], t[76], t[75], t[74], t[72], t[61], t[57], t[63], t[62], t[60], t[59], t[58], t[56], x[145], t[101], t[97], t[103], t[102], t[100], t[99], t[98], t[96], t[109], t[105], t[111], t[110], t[108], t[107], t[106], t[104], t[93], t[89], t[95], t[94], t[92], t[91], t[90], t[88], t[85], t[81], t[87], t[86], t[84], t[83], t[82], t[80], t[29], t[25], t[31], t[30], t[28], t[27], t[26], t[24], t[37], t[33], t[39], t[38], t[36], t[35], t[34], t[32], t[21], t[17], t[23], t[22], t[20], t[19], t[18], t[16], t[13], t[9], t[15], t[14], t[12], t[11], t[10], t[8], t[117], t[113], t[119], t[118], t[116], t[115], t[114], t[112], t[1], t[7], t[6], t[5], t[4], t[3], t[2], t[0]}), .y({t[1742], t[1741], t[1740], t[1739], t[1738], t[1737], t[1736], t[1735], t[1734], t[1733], t[1732], t[1731], t[1730], t[1729], t[1728], t[1727], t[1726], t[1725], t[1724], t[1723], t[1722], t[1721], t[1720], t[1719], t[1718], t[1717], t[1716], t[1715], t[1714], t[1713], t[1712], t[1711], t[1710], t[1709], t[1708], t[1707], t[1706], t[1705], t[1704], t[1703], t[1702], t[1701], t[1700], t[1699], t[1698], t[1697], t[1696], t[1695], t[1694], t[1693], t[1692], t[1691], t[1690], t[1689], t[1688], t[1687], t[1686], t[1685], t[1684], t[1683], t[1682], t[1681], t[1680], t[1679], t[1678], t[1677], t[1676], t[1675], t[1674], t[1673], t[1672], t[1671], t[1670], t[1669], t[1668], t[1667], t[1666], t[1665], t[1664], t[1663], t[1662], t[1661], t[1660], t[1659], t[1658], t[1657], t[1656], t[1655], t[1654], t[1653], t[1652], t[1651], t[1650], t[1649], t[1648], t[1647], t[1646], t[1645], t[1644], t[1643], t[1642], t[1641], t[1640], t[1639], t[1638], t[1637], t[1636], t[1635], t[1634], t[1633], t[1632], t[1631], t[1630], t[1629], t[1628], t[1627], t[1626], t[1625], t[1624], t[1623], t[1622], t[1621], t[1620], t[1619], t[1618], t[1617], t[1616], t[1615], t[1614], t[1613], t[1612], t[1611], t[1610], t[1609], t[1608], t[1607], t[1606], t[1605], t[1604], t[1603], t[1602], t[1601], t[1600], t[1599], t[1598], t[1597], t[1596], t[1595], t[1594], t[1593], t[1592], t[1591], t[1590], t[1589], t[1588], t[1587], t[1586], t[1585], t[1584], t[1583], t[1582], t[1581], t[1580], t[1579], t[1578], t[1577], t[1576], t[1575], t[1574], t[1573], t[1572], t[1571], t[1570], t[1569], t[1568], t[1567], t[1566], t[1565], t[1564], t[1563], t[1562], t[1561], t[1560], t[1559], t[1558], t[1557], t[1556], t[1555], t[1554], t[1553], t[1552], t[1551], t[1550], t[1549], t[1548], t[1547], t[1546], t[1545], t[1544], t[1543], t[1542], t[1541], t[1540], t[1539], t[1538], t[1537], t[1536], t[1535], t[1534], t[1533], t[1532], t[1531], t[1530], t[1529], t[1528], t[1527], t[1526], t[1525], t[1524], t[1523], t[1522], t[1521], t[1520], t[1519], t[1518], t[1517], t[1516], t[1515], t[1514], t[1513], t[1512], t[1511], t[1510], t[1509], t[1508], t[1507], t[1506], t[1505], t[1504], t[1503], t[1502], t[1501], t[1500], t[1499], t[1498], t[1497], t[1496], t[1495], t[1494], t[1493], t[1492], t[1491], t[1490], t[1489], t[1488], t[1487], t[1486], t[1485], t[1484], t[1483], t[1482], t[1481], t[1480], t[1479], t[1478], t[1477], t[1476], t[1475], t[1474], t[1473], t[1472], t[1471], t[1470], t[1469], t[1468], t[1467], t[1466], t[1465], t[1464], t[1463], t[1462], t[1461], t[1460], t[1459], t[1458], t[1457], t[1456], t[1455], t[1454], t[1453], t[1452], t[1451], t[1450], t[1449], t[1448], t[1447], t[1446], t[1445], t[1444], t[1443], t[1442], t[1441], t[1440], t[1439], t[1438], t[1437], t[1436], t[1435], t[1434], t[1433], t[1432], t[1431], t[1430], t[1429], t[1428], t[1427], t[1426], t[1425], t[1424], t[1423], t[1422], t[1421], t[1420], t[1419], t[1418], t[1417], t[1416], t[1415], t[1414], t[1413], t[1412], t[1411], t[1410], t[1409], t[1408], t[1407], t[1406], t[1405], t[1404], t[1403], t[1402], t[1401], t[1400], t[1399], t[1398], t[1397], t[1396], t[1395], t[1394], t[1393], t[1392], t[1391], t[1390], t[1389], t[1388], t[1387], t[1386], t[1385], t[1384], t[1383], t[1382], t[1381], t[1380], t[1379], t[1378], t[1377], t[1376], t[1375], t[1374], t[1373], t[1372], t[1371], t[1370], t[1369], t[1368], t[1367], t[1366], t[1365], t[1364], t[1363], t[1362], t[1361], t[1360], t[1359], t[1358], t[1357], t[1356], t[1355], t[1354], t[1353], t[1352], t[1351], t[1350], t[1349], t[1348], t[1347], t[1346], t[1345], t[1344], t[1343], t[1342], t[1341], t[1340], t[1339], t[1338], t[1337], t[1336], t[1335], t[1334], t[1333], t[1332], t[1331], t[1330], t[1329], t[1328], t[1327], t[1326], t[1325], t[1324], t[1323], t[1322], t[1321], t[1320], t[1319], t[1318], t[1317], t[1316], t[1315], t[1314], t[1313], t[1312], t[1311], t[1310], t[1309], t[1308], t[1307], t[1306], t[1305], t[1304], t[1303], t[1302], t[1301], t[1300], t[1299], t[1298], t[1297], t[1296], t[1295]}));
  Reg1 Reg1_inst(.x({t[1283], t[1285], t[1282], t[1284], t[1294], t[1289], t[1291], t[1226], t[1227], t[1228], t[1229], t[1230], t[1231], t[1232], t[1233], t[1234], t[1235], t[1236], t[1237], t[1238], t[1239], t[1240], t[1241], t[1242], t[1243], t[1244], t[1245], t[1246], t[1247], t[1248], t[1249], t[1250], t[1251], t[1252], t[1253], t[1254], t[1255], t[1256], t[1257], t[1258], t[1259], t[1260], t[1261], t[1202], t[1203], t[1204], t[1205], t[1206], t[1207], t[1208], t[1209], t[1210], t[1211], t[1212], t[1213], t[1214], t[1215], t[1216], t[1217], t[1218], t[1219], t[1220], t[1221], t[1222], t[1223], t[1224], t[1225], t[1265], t[1264], t[1263], t[1262], t[1280], t[1293], t[1281], t[1287], t[1292], t[1286], t[1162], t[1163], t[1164], t[1165], t[1166], t[1167], t[1168], t[1169], t[1170], t[1171], t[1172], t[1173], t[1174], t[1175], t[1176], t[1177], t[1178], t[1179], t[1180], t[1181], t[1182], t[1183], t[1184], t[1185], t[1186], t[1187], t[1188], t[1189], t[1190], t[1191], t[1192], t[1193], t[1194], t[1195], t[1196], t[1197], t[1122], t[1123], t[1124], t[1125], t[1126], t[1127], t[1128], t[1129], t[1130], t[1131], t[1132], t[1133], t[1134], t[1135], t[1136], t[1137], t[1138], t[1139], t[1140], t[1141], t[1142], t[1143], t[1144], t[1145], t[1146], t[1147], t[1148], t[1149], t[1150], t[1151], t[1152], t[1153], t[1154], t[1155], t[1156], t[1157], t[1158], t[1159], t[1160], t[1161], t[1198], t[1199], t[1200], t[1201], t[1270], t[1269], t[1267], t[1268], t[1272], t[1275], t[1274], t[1273], t[1271], t[1278], t[1276], t[1277], t[1266], t[1121], t[1279], t[1290], t[1288], x[144]}), .y({t[608], t[606], t[605], t[604], t[597], t[595], t[594], t[593], t[586], t[584], t[583], t[582], t[575], t[573], t[572], t[571], t[564], t[562], t[561], t[560], t[553], t[551], t[550], t[549], t[542], t[540], t[539], t[538], t[531], t[529], t[528], t[527], t[520], t[518], t[517], t[516], t[509], t[507], t[506], t[505], t[498], t[496], t[495], t[494], t[487], t[485], t[484], t[483], t[476], t[474], t[473], t[472], t[465], t[463], t[462], t[461], t[454], t[452], t[451], t[450], t[443], t[441], t[440], t[439], t[432], t[430], t[429], t[428], t[421], t[419], t[418], t[417], t[410], t[408], t[407], t[406], t[399], t[397], t[396], t[395], t[388], t[386], t[385], t[384], t[377], t[375], t[374], t[373], t[366], t[364], t[363], t[362], t[355], t[353], t[352], t[351], t[344], t[342], t[341], t[340], t[333], t[331], t[330], t[329], t[322], t[320], t[319], t[318], t[311], t[309], t[308], t[307], t[300], t[298], t[297], t[296], t[289], t[287], t[286], t[285], t[278], t[276], t[275], t[274], t[267], t[265], t[264], t[263], t[256], t[254], t[253], t[252], t[245], t[243], t[242], t[241], t[234], t[232], t[231], t[230], t[223], t[221], t[220], t[219], t[212], t[210], t[209], t[208], t[200], t[192], t[184], t[176], t[168], t[160], t[152], t[144], t[136], t[128], t[120], t[112], t[104], t[96], t[88], t[80], t[72], t[64], t[56], t[48], t[40], t[32], t[24], t[16], t[8], t[0]}));
  Reg2 Reg2_inst(.x({t[1742], t[1741], t[1740], t[1739], t[1738], t[1737], t[1736], t[1427], t[1426], t[1425], t[1424], t[1423], t[1422], t[1421], t[1448], t[1447], t[1446], t[1445], t[1444], t[1443], t[1442], t[1441], t[1440], t[1439], t[1438], t[1437], t[1436], t[1435], t[1553], t[1552], t[1551], t[1550], t[1549], t[1548], t[1547], t[1546], t[1545], t[1544], t[1543], t[1542], t[1541], t[1540], t[1539], t[1538], t[1537], t[1536], t[1535], t[1534], t[1533], t[1532], t[1531], t[1530], t[1529], t[1528], t[1527], t[1526], t[1525], t[1524], t[1523], t[1522], t[1521], t[1520], t[1519], t[1518], t[1517], t[1516], t[1515], t[1514], t[1513], t[1512], t[1511], t[1510], t[1509], t[1508], t[1507], t[1506], t[1505], t[1504], t[1503], t[1502], t[1501], t[1500], t[1499], t[1498], t[1497], t[1496], t[1495], t[1494], t[1493], t[1492], t[1491], t[1665], t[1664], t[1663], t[1662], t[1661], t[1660], t[1659], t[1658], t[1657], t[1656], t[1655], t[1654], t[1653], t[1652], t[1651], t[1650], t[1649], t[1648], t[1647], t[1646], t[1645], t[1644], t[1643], t[1642], t[1641], t[1640], t[1639], t[1638], t[1637], t[1636], t[1635], t[1634], t[1633], t[1632], t[1631], t[1630], t[1629], t[1628], t[1627], t[1626], t[1625], t[1624], t[1490], t[1489], t[1488], t[1487], t[1486], t[1485], t[1484], t[1462], t[1461], t[1460], t[1459], t[1458], t[1457], t[1456], t[1455], t[1454], t[1453], t[1452], t[1451], t[1450], t[1449], t[1483], t[1482], t[1481], t[1480], t[1479], t[1478], t[1477], t[1476], t[1475], t[1474], t[1473], t[1472], t[1471], t[1470], t[1434], t[1433], t[1432], t[1431], t[1430], t[1429], t[1428], t[1469], t[1468], t[1467], t[1466], t[1465], t[1464], t[1463], t[1623], t[1622], t[1621], t[1620], t[1619], t[1618], t[1617], t[1616], t[1615], t[1614], t[1613], t[1612], t[1611], t[1610], t[1609], t[1608], t[1607], t[1606], t[1605], t[1604], t[1603], t[1602], t[1601], t[1600], t[1599], t[1598], t[1597], t[1596], t[1595], t[1594], t[1593], t[1592], t[1591], t[1590], t[1589], t[1588], t[1587], t[1586], t[1585], t[1584], t[1583], t[1582], t[1581], t[1580], t[1579], t[1578], t[1577], t[1576], t[1575], t[1574], t[1573], t[1572], t[1571], t[1570], t[1569], t[1568], t[1567], t[1566], t[1565], t[1564], t[1563], t[1562], t[1561], t[1735], t[1734], t[1733], t[1732], t[1731], t[1730], t[1729], t[1728], t[1727], t[1726], t[1725], t[1724], t[1723], t[1722], t[1721], t[1720], t[1719], t[1718], t[1717], t[1716], t[1715], t[1714], t[1713], t[1712], t[1711], t[1710], t[1709], t[1708], t[1707], t[1706], t[1705], t[1704], t[1703], t[1702], t[1701], t[1700], t[1699], t[1698], t[1697], t[1696], t[1695], t[1694], t[1693], t[1692], t[1691], t[1690], t[1689], t[1688], t[1687], t[1686], t[1685], t[1684], t[1683], t[1682], t[1681], t[1680], t[1679], t[1678], t[1677], t[1676], t[1675], t[1674], t[1673], t[1672], t[1671], t[1670], t[1669], t[1668], t[1667], t[1666], t[1560], t[1559], t[1558], t[1557], t[1556], t[1555], t[1554], t[1399], t[1398], t[1397], t[1396], t[1395], t[1394], t[1393], t[1392], t[1391], t[1390], t[1389], t[1388], t[1387], t[1386], t[1385], t[1384], t[1383], t[1382], t[1381], t[1380], t[1379], t[1378], t[1377], t[1376], t[1375], t[1374], t[1373], t[1372], t[1371], t[1370], t[1369], t[1368], t[1367], t[1366], t[1365], t[1364], t[1363], t[1362], t[1361], t[1360], t[1359], t[1358], t[1357], t[1356], t[1355], t[1354], t[1353], t[1352], t[1351], t[1350], t[1349], t[1348], t[1347], t[1346], t[1345], t[1344], t[1343], t[1342], t[1341], t[1340], t[1339], t[1338], t[1337], t[1336], t[1335], t[1334], t[1333], t[1332], t[1331], t[1330], t[1329], t[1328], t[1327], t[1326], t[1325], t[1324], t[1323], t[1322], t[1321], t[1320], t[1319], t[1318], t[1317], t[1316], t[1315], t[1314], t[1313], t[1312], t[1311], t[1310], t[1309], t[1308], t[1307], t[1306], t[1305], t[1304], t[1303], t[1302], t[1406], t[1405], t[1404], t[1403], t[1402], t[1401], t[1400], t[1420], t[1419], t[1418], t[1417], t[1416], t[1415], t[1414], t[1413], t[1412], t[1411], t[1410], t[1409], t[1408], t[1407], x[144]}), .y({t[614], t[613], t[612], t[611], t[610], t[609], t[607], t[603], t[602], t[601], t[600], t[599], t[598], t[596], t[592], t[591], t[590], t[589], t[588], t[587], t[585], t[581], t[580], t[579], t[578], t[577], t[576], t[574], t[570], t[569], t[568], t[567], t[566], t[565], t[563], t[559], t[558], t[557], t[556], t[555], t[554], t[552], t[548], t[547], t[546], t[545], t[544], t[543], t[541], t[537], t[536], t[535], t[534], t[533], t[532], t[530], t[526], t[525], t[524], t[523], t[522], t[521], t[519], t[515], t[514], t[513], t[512], t[511], t[510], t[508], t[504], t[503], t[502], t[501], t[500], t[499], t[497], t[493], t[492], t[491], t[490], t[489], t[488], t[486], t[482], t[481], t[480], t[479], t[478], t[477], t[475], t[471], t[470], t[469], t[468], t[467], t[466], t[464], t[460], t[459], t[458], t[457], t[456], t[455], t[453], t[449], t[448], t[447], t[446], t[445], t[444], t[442], t[438], t[437], t[436], t[435], t[434], t[433], t[431], t[427], t[426], t[425], t[424], t[423], t[422], t[420], t[416], t[415], t[414], t[413], t[412], t[411], t[409], t[405], t[404], t[403], t[402], t[401], t[400], t[398], t[394], t[393], t[392], t[391], t[390], t[389], t[387], t[383], t[382], t[381], t[380], t[379], t[378], t[376], t[372], t[371], t[370], t[369], t[368], t[367], t[365], t[361], t[360], t[359], t[358], t[357], t[356], t[354], t[350], t[349], t[348], t[347], t[346], t[345], t[343], t[339], t[338], t[337], t[336], t[335], t[334], t[332], t[328], t[327], t[326], t[325], t[324], t[323], t[321], t[317], t[316], t[315], t[314], t[313], t[312], t[310], t[306], t[305], t[304], t[303], t[302], t[301], t[299], t[295], t[294], t[293], t[292], t[291], t[290], t[288], t[284], t[283], t[282], t[281], t[280], t[279], t[277], t[273], t[272], t[271], t[270], t[269], t[268], t[266], t[262], t[261], t[260], t[259], t[258], t[257], t[255], t[251], t[250], t[249], t[248], t[247], t[246], t[244], t[240], t[239], t[238], t[237], t[236], t[235], t[233], t[229], t[228], t[227], t[226], t[225], t[224], t[222], t[218], t[217], t[216], t[215], t[214], t[213], t[211], t[207], t[206], t[205], t[204], t[203], t[202], t[201], t[199], t[198], t[197], t[196], t[195], t[194], t[193], t[191], t[190], t[189], t[188], t[187], t[186], t[185], t[183], t[182], t[181], t[180], t[179], t[178], t[177], t[175], t[174], t[173], t[172], t[171], t[170], t[169], t[167], t[166], t[165], t[164], t[163], t[162], t[161], t[159], t[158], t[157], t[156], t[155], t[154], t[153], t[151], t[150], t[149], t[148], t[147], t[146], t[145], t[143], t[142], t[141], t[140], t[139], t[138], t[137], t[135], t[134], t[133], t[132], t[131], t[130], t[129], t[127], t[126], t[125], t[124], t[123], t[122], t[121], t[119], t[118], t[117], t[116], t[115], t[114], t[113], t[111], t[110], t[109], t[108], t[107], t[106], t[105], t[103], t[102], t[101], t[100], t[99], t[98], t[97], t[95], t[94], t[93], t[92], t[91], t[90], t[89], t[87], t[86], t[85], t[84], t[83], t[82], t[81], t[79], t[78], t[77], t[76], t[75], t[74], t[73], t[71], t[70], t[69], t[68], t[67], t[66], t[65], t[63], t[62], t[61], t[60], t[59], t[58], t[57], t[55], t[54], t[53], t[52], t[51], t[50], t[49], t[47], t[46], t[45], t[44], t[43], t[42], t[41], t[39], t[38], t[37], t[36], t[35], t[34], t[33], t[31], t[30], t[29], t[28], t[27], t[26], t[25], t[23], t[22], t[21], t[20], t[19], t[18], t[17], t[15], t[14], t[13], t[12], t[11], t[10], t[9], t[7], t[6], t[5], t[4], t[3], t[2], t[1]}));
  multiplexer #(.WIDTH(65)) multiplexer_inst(.s({t[1295], t[1296], t[1297], t[1298], t[1299], t[1300], t[1301], t[1056]}), .d({t[1117], t[1118], t[1119], t[1120], t[1113], t[1114], t[1115], t[1116], t[1109], t[1110], t[1111], t[1112], t[1105], t[1106], t[1107], t[1108], t[1101], t[1102], t[1103], t[1104], t[1097], t[1098], t[1099], t[1100], t[1093], t[1094], t[1095], t[1096], t[1089], t[1090], t[1091], t[1092], t[1085], t[1086], t[1087], t[1088], t[1081], t[1082], t[1083], t[1084], t[1077], t[1078], t[1079], t[1080], t[1073], t[1074], t[1075], t[1076], t[1069], t[1070], t[1071], t[1072], t[1065], t[1066], t[1067], t[1068], t[1061], t[1062], t[1063], t[1064], t[1060], t[1059], t[1058], t[1057], t[1295]}), .q({y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], y[8], y[9], y[10], y[11], y[12], y[13], y[14], y[15], y[16], y[17], y[18], y[19], y[20], y[21], y[22], y[23], y[24], y[25], y[26], y[27], y[28], y[29], y[30], y[31], y[32], y[33], y[34], y[35], y[36], y[37], y[38], y[39], y[40], y[41], y[42], y[43], y[44], y[45], y[46], y[47], y[48], y[49], y[50], y[51], y[52], y[53], y[54], y[55], y[56], y[57], y[58], y[59], y[60], y[61], y[62], y[63], y[64]}));
endmodule

module register_stage(clk, D, Q);
  parameter WIDTH = 8;
  input clk;
  input [WIDTH-1:0] D;
  output [WIDTH-1:0] Q;

  reg [WIDTH-1:0] s_current_state;
  wire [WIDTH-1:0] s_next_state;
  assign s_next_state = D;
  always @ (posedge clk)
  begin
      s_current_state <= s_next_state;
  end
  assign Q = s_current_state;
endmodule

module multiplexer(s, d, q);
  parameter WIDTH = 8;
  input [7:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  muxtree #(.WIDTH(65)) inst_0(.s(s), .d({d[0],d[1],d[2],d[3],d[4],d[5],d[6],d[7],d[8],d[9],d[10],d[11],d[12],d[13],d[14],d[15],d[16],d[17],d[18],d[19],d[20],d[21],d[22],d[23],d[24],d[25],d[26],d[27],d[28],d[29],d[30],d[31],d[32],d[33],d[34],d[35],d[36],d[37],d[38],d[39],d[40],d[41],d[42],d[43],d[44],d[45],d[46],d[47],d[48],d[49],d[50],d[51],d[52],d[53],d[54],d[55],d[56],d[57],d[58],d[59],d[60],d[61],d[62],d[63],d[64]}), .q({q[0],q[1],q[2],q[3],q[4],q[5],q[6],q[7],q[8],q[9],q[10],q[11],q[12],q[13],q[14],q[15],q[16],q[17],q[18],q[19],q[20],q[21],q[22],q[23],q[24],q[25],q[26],q[27],q[28],q[29],q[30],q[31],q[32],q[33],q[34],q[35],q[36],q[37],q[38],q[39],q[40],q[41],q[42],q[43],q[44],q[45],q[46],q[47],q[48],q[49],q[50],q[51],q[52],q[53],q[54],q[55],q[56],q[57],q[58],q[59],q[60],q[61],q[62],q[63],q[64]}));
endmodule

module muxtree(s, d, q);
  parameter WIDTH = 8;
  input [7:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  wire [WIDTH-1:0] v0_0;
  wire [WIDTH-1:0] v0_1;
  wire [WIDTH-1:0] v1_0;
  wire [WIDTH-1:0] v1_1;
  wire [WIDTH-1:0] v1_2;
  wire [WIDTH-1:0] v1_3;
  wire [WIDTH-1:0] v2_0;
  wire [WIDTH-1:0] v2_1;
  wire [WIDTH-1:0] v2_2;
  wire [WIDTH-1:0] v2_3;
  wire [WIDTH-1:0] v2_4;
  wire [WIDTH-1:0] v2_5;
  wire [WIDTH-1:0] v2_6;
  wire [WIDTH-1:0] v2_7;
  wire [WIDTH-1:0] v3_0;
  wire [WIDTH-1:0] v3_1;
  wire [WIDTH-1:0] v3_2;
  wire [WIDTH-1:0] v3_3;
  wire [WIDTH-1:0] v3_4;
  wire [WIDTH-1:0] v3_5;
  wire [WIDTH-1:0] v3_6;
  wire [WIDTH-1:0] v3_7;
  wire [WIDTH-1:0] v3_8;
  wire [WIDTH-1:0] v3_9;
  wire [WIDTH-1:0] v3_10;
  wire [WIDTH-1:0] v3_11;
  wire [WIDTH-1:0] v3_12;
  wire [WIDTH-1:0] v3_13;
  wire [WIDTH-1:0] v3_14;
  wire [WIDTH-1:0] v3_15;
  wire [WIDTH-1:0] v4_0;
  wire [WIDTH-1:0] v4_1;
  wire [WIDTH-1:0] v4_2;
  wire [WIDTH-1:0] v4_3;
  wire [WIDTH-1:0] v4_4;
  wire [WIDTH-1:0] v4_5;
  wire [WIDTH-1:0] v4_6;
  wire [WIDTH-1:0] v4_7;
  wire [WIDTH-1:0] v4_8;
  wire [WIDTH-1:0] v4_9;
  wire [WIDTH-1:0] v4_10;
  wire [WIDTH-1:0] v4_11;
  wire [WIDTH-1:0] v4_12;
  wire [WIDTH-1:0] v4_13;
  wire [WIDTH-1:0] v4_14;
  wire [WIDTH-1:0] v4_15;
  wire [WIDTH-1:0] v4_16;
  wire [WIDTH-1:0] v4_17;
  wire [WIDTH-1:0] v4_18;
  wire [WIDTH-1:0] v4_19;
  wire [WIDTH-1:0] v4_20;
  wire [WIDTH-1:0] v4_21;
  wire [WIDTH-1:0] v4_22;
  wire [WIDTH-1:0] v4_23;
  wire [WIDTH-1:0] v4_24;
  wire [WIDTH-1:0] v4_25;
  wire [WIDTH-1:0] v4_26;
  wire [WIDTH-1:0] v4_27;
  wire [WIDTH-1:0] v4_28;
  wire [WIDTH-1:0] v4_29;
  wire [WIDTH-1:0] v4_30;
  wire [WIDTH-1:0] v4_31;
  wire [WIDTH-1:0] v5_0;
  wire [WIDTH-1:0] v5_1;
  wire [WIDTH-1:0] v5_2;
  wire [WIDTH-1:0] v5_3;
  wire [WIDTH-1:0] v5_4;
  wire [WIDTH-1:0] v5_5;
  wire [WIDTH-1:0] v5_6;
  wire [WIDTH-1:0] v5_7;
  wire [WIDTH-1:0] v5_8;
  wire [WIDTH-1:0] v5_9;
  wire [WIDTH-1:0] v5_10;
  wire [WIDTH-1:0] v5_11;
  wire [WIDTH-1:0] v5_12;
  wire [WIDTH-1:0] v5_13;
  wire [WIDTH-1:0] v5_14;
  wire [WIDTH-1:0] v5_15;
  wire [WIDTH-1:0] v5_16;
  wire [WIDTH-1:0] v5_17;
  wire [WIDTH-1:0] v5_18;
  wire [WIDTH-1:0] v5_19;
  wire [WIDTH-1:0] v5_20;
  wire [WIDTH-1:0] v5_21;
  wire [WIDTH-1:0] v5_22;
  wire [WIDTH-1:0] v5_23;
  wire [WIDTH-1:0] v5_24;
  wire [WIDTH-1:0] v5_25;
  wire [WIDTH-1:0] v5_26;
  wire [WIDTH-1:0] v5_27;
  wire [WIDTH-1:0] v5_28;
  wire [WIDTH-1:0] v5_29;
  wire [WIDTH-1:0] v5_30;
  wire [WIDTH-1:0] v5_31;
  wire [WIDTH-1:0] v5_32;
  wire [WIDTH-1:0] v5_33;
  wire [WIDTH-1:0] v5_34;
  wire [WIDTH-1:0] v5_35;
  wire [WIDTH-1:0] v5_36;
  wire [WIDTH-1:0] v5_37;
  wire [WIDTH-1:0] v5_38;
  wire [WIDTH-1:0] v5_39;
  wire [WIDTH-1:0] v5_40;
  wire [WIDTH-1:0] v5_41;
  wire [WIDTH-1:0] v5_42;
  wire [WIDTH-1:0] v5_43;
  wire [WIDTH-1:0] v5_44;
  wire [WIDTH-1:0] v5_45;
  wire [WIDTH-1:0] v5_46;
  wire [WIDTH-1:0] v5_47;
  wire [WIDTH-1:0] v5_48;
  wire [WIDTH-1:0] v5_49;
  wire [WIDTH-1:0] v5_50;
  wire [WIDTH-1:0] v5_51;
  wire [WIDTH-1:0] v5_52;
  wire [WIDTH-1:0] v5_53;
  wire [WIDTH-1:0] v5_54;
  wire [WIDTH-1:0] v5_55;
  wire [WIDTH-1:0] v5_56;
  wire [WIDTH-1:0] v5_57;
  wire [WIDTH-1:0] v5_58;
  wire [WIDTH-1:0] v5_59;
  wire [WIDTH-1:0] v5_60;
  wire [WIDTH-1:0] v5_61;
  wire [WIDTH-1:0] v5_62;
  wire [WIDTH-1:0] v5_63;
  wire [WIDTH-1:0] v6_0;
  wire [WIDTH-1:0] v6_1;
  wire [WIDTH-1:0] v6_2;
  wire [WIDTH-1:0] v6_3;
  wire [WIDTH-1:0] v6_4;
  wire [WIDTH-1:0] v6_5;
  wire [WIDTH-1:0] v6_6;
  wire [WIDTH-1:0] v6_7;
  wire [WIDTH-1:0] v6_8;
  wire [WIDTH-1:0] v6_9;
  wire [WIDTH-1:0] v6_10;
  wire [WIDTH-1:0] v6_11;
  wire [WIDTH-1:0] v6_12;
  wire [WIDTH-1:0] v6_13;
  wire [WIDTH-1:0] v6_14;
  wire [WIDTH-1:0] v6_15;
  wire [WIDTH-1:0] v6_16;
  wire [WIDTH-1:0] v6_17;
  wire [WIDTH-1:0] v6_18;
  wire [WIDTH-1:0] v6_19;
  wire [WIDTH-1:0] v6_20;
  wire [WIDTH-1:0] v6_21;
  wire [WIDTH-1:0] v6_22;
  wire [WIDTH-1:0] v6_23;
  wire [WIDTH-1:0] v6_24;
  wire [WIDTH-1:0] v6_25;
  wire [WIDTH-1:0] v6_26;
  wire [WIDTH-1:0] v6_27;
  wire [WIDTH-1:0] v6_28;
  wire [WIDTH-1:0] v6_29;
  wire [WIDTH-1:0] v6_30;
  wire [WIDTH-1:0] v6_31;
  wire [WIDTH-1:0] v6_32;
  wire [WIDTH-1:0] v6_33;
  wire [WIDTH-1:0] v6_34;
  wire [WIDTH-1:0] v6_35;
  wire [WIDTH-1:0] v6_36;
  wire [WIDTH-1:0] v6_37;
  wire [WIDTH-1:0] v6_38;
  wire [WIDTH-1:0] v6_39;
  wire [WIDTH-1:0] v6_40;
  wire [WIDTH-1:0] v6_41;
  wire [WIDTH-1:0] v6_42;
  wire [WIDTH-1:0] v6_43;
  wire [WIDTH-1:0] v6_44;
  wire [WIDTH-1:0] v6_45;
  wire [WIDTH-1:0] v6_46;
  wire [WIDTH-1:0] v6_47;
  wire [WIDTH-1:0] v6_48;
  wire [WIDTH-1:0] v6_49;
  wire [WIDTH-1:0] v6_50;
  wire [WIDTH-1:0] v6_51;
  wire [WIDTH-1:0] v6_52;
  wire [WIDTH-1:0] v6_53;
  wire [WIDTH-1:0] v6_54;
  wire [WIDTH-1:0] v6_55;
  wire [WIDTH-1:0] v6_56;
  wire [WIDTH-1:0] v6_57;
  wire [WIDTH-1:0] v6_58;
  wire [WIDTH-1:0] v6_59;
  wire [WIDTH-1:0] v6_60;
  wire [WIDTH-1:0] v6_61;
  wire [WIDTH-1:0] v6_62;
  wire [WIDTH-1:0] v6_63;
  wire [WIDTH-1:0] v6_64;
  wire [WIDTH-1:0] v6_65;
  wire [WIDTH-1:0] v6_66;
  wire [WIDTH-1:0] v6_67;
  wire [WIDTH-1:0] v6_68;
  wire [WIDTH-1:0] v6_69;
  wire [WIDTH-1:0] v6_70;
  wire [WIDTH-1:0] v6_71;
  wire [WIDTH-1:0] v6_72;
  wire [WIDTH-1:0] v6_73;
  wire [WIDTH-1:0] v6_74;
  wire [WIDTH-1:0] v6_75;
  wire [WIDTH-1:0] v6_76;
  wire [WIDTH-1:0] v6_77;
  wire [WIDTH-1:0] v6_78;
  wire [WIDTH-1:0] v6_79;
  wire [WIDTH-1:0] v6_80;
  wire [WIDTH-1:0] v6_81;
  wire [WIDTH-1:0] v6_82;
  wire [WIDTH-1:0] v6_83;
  wire [WIDTH-1:0] v6_84;
  wire [WIDTH-1:0] v6_85;
  wire [WIDTH-1:0] v6_86;
  wire [WIDTH-1:0] v6_87;
  wire [WIDTH-1:0] v6_88;
  wire [WIDTH-1:0] v6_89;
  wire [WIDTH-1:0] v6_90;
  wire [WIDTH-1:0] v6_91;
  wire [WIDTH-1:0] v6_92;
  wire [WIDTH-1:0] v6_93;
  wire [WIDTH-1:0] v6_94;
  wire [WIDTH-1:0] v6_95;
  wire [WIDTH-1:0] v6_96;
  wire [WIDTH-1:0] v6_97;
  wire [WIDTH-1:0] v6_98;
  wire [WIDTH-1:0] v6_99;
  wire [WIDTH-1:0] v6_100;
  wire [WIDTH-1:0] v6_101;
  wire [WIDTH-1:0] v6_102;
  wire [WIDTH-1:0] v6_103;
  wire [WIDTH-1:0] v6_104;
  wire [WIDTH-1:0] v6_105;
  wire [WIDTH-1:0] v6_106;
  wire [WIDTH-1:0] v6_107;
  wire [WIDTH-1:0] v6_108;
  wire [WIDTH-1:0] v6_109;
  wire [WIDTH-1:0] v6_110;
  wire [WIDTH-1:0] v6_111;
  wire [WIDTH-1:0] v6_112;
  wire [WIDTH-1:0] v6_113;
  wire [WIDTH-1:0] v6_114;
  wire [WIDTH-1:0] v6_115;
  wire [WIDTH-1:0] v6_116;
  wire [WIDTH-1:0] v6_117;
  wire [WIDTH-1:0] v6_118;
  wire [WIDTH-1:0] v6_119;
  wire [WIDTH-1:0] v6_120;
  wire [WIDTH-1:0] v6_121;
  wire [WIDTH-1:0] v6_122;
  wire [WIDTH-1:0] v6_123;
  wire [WIDTH-1:0] v6_124;
  wire [WIDTH-1:0] v6_125;
  wire [WIDTH-1:0] v6_126;
  wire [WIDTH-1:0] v6_127;

  assign q = s[0] ? v0_1 : {WIDTH{1'b0}};

  assign v0_0 = s[1] ? {WIDTH{1'b0}} : v1_0;
  assign v0_1 = s[1] ? {WIDTH{1'b0}} : v1_2;

  assign v1_0 = s[2] ? {WIDTH{1'b0}} : v2_0;
  assign v1_1 = s[2] ? {WIDTH{1'b0}} : v2_2;
  assign v1_2 = s[2] ? {WIDTH{1'b0}} : v2_4;
  assign v1_3 = s[2] ? {WIDTH{1'b0}} : v2_6;

  assign v2_0 = s[3] ? {WIDTH{1'b0}} : v3_0;
  assign v2_1 = s[3] ? {WIDTH{1'b0}} : v3_2;
  assign v2_2 = s[3] ? {WIDTH{1'b0}} : v3_4;
  assign v2_3 = s[3] ? {WIDTH{1'b0}} : v3_6;
  assign v2_4 = s[3] ? {WIDTH{1'b0}} : v3_8;
  assign v2_5 = s[3] ? {WIDTH{1'b0}} : v3_10;
  assign v2_6 = s[3] ? {WIDTH{1'b0}} : v3_12;
  assign v2_7 = s[3] ? {WIDTH{1'b0}} : v3_14;

  assign v3_0 = s[4] ? v4_1 : {WIDTH{1'b0}};
  assign v3_1 = s[4] ? v4_3 : {WIDTH{1'b0}};
  assign v3_2 = s[4] ? v4_5 : {WIDTH{1'b0}};
  assign v3_3 = s[4] ? v4_7 : {WIDTH{1'b0}};
  assign v3_4 = s[4] ? v4_9 : {WIDTH{1'b0}};
  assign v3_5 = s[4] ? v4_11 : {WIDTH{1'b0}};
  assign v3_6 = s[4] ? v4_13 : {WIDTH{1'b0}};
  assign v3_7 = s[4] ? v4_15 : {WIDTH{1'b0}};
  assign v3_8 = s[4] ? v4_17 : {WIDTH{1'b0}};
  assign v3_9 = s[4] ? v4_19 : {WIDTH{1'b0}};
  assign v3_10 = s[4] ? v4_21 : {WIDTH{1'b0}};
  assign v3_11 = s[4] ? v4_23 : {WIDTH{1'b0}};
  assign v3_12 = s[4] ? v4_25 : {WIDTH{1'b0}};
  assign v3_13 = s[4] ? v4_27 : {WIDTH{1'b0}};
  assign v3_14 = s[4] ? v4_29 : {WIDTH{1'b0}};
  assign v3_15 = s[4] ? v4_31 : {WIDTH{1'b0}};

  assign v4_0 = s[5] ? v5_1 : {WIDTH{1'b0}};
  assign v4_1 = s[5] ? v5_3 : {WIDTH{1'b0}};
  assign v4_2 = s[5] ? v5_5 : {WIDTH{1'b0}};
  assign v4_3 = s[5] ? v5_7 : {WIDTH{1'b0}};
  assign v4_4 = s[5] ? v5_9 : {WIDTH{1'b0}};
  assign v4_5 = s[5] ? v5_11 : {WIDTH{1'b0}};
  assign v4_6 = s[5] ? v5_13 : {WIDTH{1'b0}};
  assign v4_7 = s[5] ? v5_15 : {WIDTH{1'b0}};
  assign v4_8 = s[5] ? v5_17 : {WIDTH{1'b0}};
  assign v4_9 = s[5] ? v5_19 : {WIDTH{1'b0}};
  assign v4_10 = s[5] ? v5_21 : {WIDTH{1'b0}};
  assign v4_11 = s[5] ? v5_23 : {WIDTH{1'b0}};
  assign v4_12 = s[5] ? v5_25 : {WIDTH{1'b0}};
  assign v4_13 = s[5] ? v5_27 : {WIDTH{1'b0}};
  assign v4_14 = s[5] ? v5_29 : {WIDTH{1'b0}};
  assign v4_15 = s[5] ? v5_31 : {WIDTH{1'b0}};
  assign v4_16 = s[5] ? v5_33 : {WIDTH{1'b0}};
  assign v4_17 = s[5] ? v5_35 : {WIDTH{1'b0}};
  assign v4_18 = s[5] ? v5_37 : {WIDTH{1'b0}};
  assign v4_19 = s[5] ? v5_39 : {WIDTH{1'b0}};
  assign v4_20 = s[5] ? v5_41 : {WIDTH{1'b0}};
  assign v4_21 = s[5] ? v5_43 : {WIDTH{1'b0}};
  assign v4_22 = s[5] ? v5_45 : {WIDTH{1'b0}};
  assign v4_23 = s[5] ? v5_47 : {WIDTH{1'b0}};
  assign v4_24 = s[5] ? v5_49 : {WIDTH{1'b0}};
  assign v4_25 = s[5] ? v5_51 : {WIDTH{1'b0}};
  assign v4_26 = s[5] ? v5_53 : {WIDTH{1'b0}};
  assign v4_27 = s[5] ? v5_55 : {WIDTH{1'b0}};
  assign v4_28 = s[5] ? v5_57 : {WIDTH{1'b0}};
  assign v4_29 = s[5] ? v5_59 : {WIDTH{1'b0}};
  assign v4_30 = s[5] ? v5_61 : {WIDTH{1'b0}};
  assign v4_31 = s[5] ? v5_63 : {WIDTH{1'b0}};

  assign v5_0 = s[6] ? v6_1 : {WIDTH{1'b0}};
  assign v5_1 = s[6] ? v6_3 : {WIDTH{1'b0}};
  assign v5_2 = s[6] ? v6_5 : {WIDTH{1'b0}};
  assign v5_3 = s[6] ? v6_7 : {WIDTH{1'b0}};
  assign v5_4 = s[6] ? v6_9 : {WIDTH{1'b0}};
  assign v5_5 = s[6] ? v6_11 : {WIDTH{1'b0}};
  assign v5_6 = s[6] ? v6_13 : {WIDTH{1'b0}};
  assign v5_7 = s[6] ? v6_15 : {WIDTH{1'b0}};
  assign v5_8 = s[6] ? v6_17 : {WIDTH{1'b0}};
  assign v5_9 = s[6] ? v6_19 : {WIDTH{1'b0}};
  assign v5_10 = s[6] ? v6_21 : {WIDTH{1'b0}};
  assign v5_11 = s[6] ? v6_23 : {WIDTH{1'b0}};
  assign v5_12 = s[6] ? v6_25 : {WIDTH{1'b0}};
  assign v5_13 = s[6] ? v6_27 : {WIDTH{1'b0}};
  assign v5_14 = s[6] ? v6_29 : {WIDTH{1'b0}};
  assign v5_15 = s[6] ? v6_31 : {WIDTH{1'b0}};
  assign v5_16 = s[6] ? v6_33 : {WIDTH{1'b0}};
  assign v5_17 = s[6] ? v6_35 : {WIDTH{1'b0}};
  assign v5_18 = s[6] ? v6_37 : {WIDTH{1'b0}};
  assign v5_19 = s[6] ? v6_39 : {WIDTH{1'b0}};
  assign v5_20 = s[6] ? v6_41 : {WIDTH{1'b0}};
  assign v5_21 = s[6] ? v6_43 : {WIDTH{1'b0}};
  assign v5_22 = s[6] ? v6_45 : {WIDTH{1'b0}};
  assign v5_23 = s[6] ? v6_47 : {WIDTH{1'b0}};
  assign v5_24 = s[6] ? v6_49 : {WIDTH{1'b0}};
  assign v5_25 = s[6] ? v6_51 : {WIDTH{1'b0}};
  assign v5_26 = s[6] ? v6_53 : {WIDTH{1'b0}};
  assign v5_27 = s[6] ? v6_55 : {WIDTH{1'b0}};
  assign v5_28 = s[6] ? v6_57 : {WIDTH{1'b0}};
  assign v5_29 = s[6] ? v6_59 : {WIDTH{1'b0}};
  assign v5_30 = s[6] ? v6_61 : {WIDTH{1'b0}};
  assign v5_31 = s[6] ? v6_63 : {WIDTH{1'b0}};
  assign v5_32 = s[6] ? v6_65 : {WIDTH{1'b0}};
  assign v5_33 = s[6] ? v6_67 : {WIDTH{1'b0}};
  assign v5_34 = s[6] ? v6_69 : {WIDTH{1'b0}};
  assign v5_35 = s[6] ? v6_71 : {WIDTH{1'b0}};
  assign v5_36 = s[6] ? v6_73 : {WIDTH{1'b0}};
  assign v5_37 = s[6] ? v6_75 : {WIDTH{1'b0}};
  assign v5_38 = s[6] ? v6_77 : {WIDTH{1'b0}};
  assign v5_39 = s[6] ? v6_79 : {WIDTH{1'b0}};
  assign v5_40 = s[6] ? v6_81 : {WIDTH{1'b0}};
  assign v5_41 = s[6] ? v6_83 : {WIDTH{1'b0}};
  assign v5_42 = s[6] ? v6_85 : {WIDTH{1'b0}};
  assign v5_43 = s[6] ? v6_87 : {WIDTH{1'b0}};
  assign v5_44 = s[6] ? v6_89 : {WIDTH{1'b0}};
  assign v5_45 = s[6] ? v6_91 : {WIDTH{1'b0}};
  assign v5_46 = s[6] ? v6_93 : {WIDTH{1'b0}};
  assign v5_47 = s[6] ? v6_95 : {WIDTH{1'b0}};
  assign v5_48 = s[6] ? v6_97 : {WIDTH{1'b0}};
  assign v5_49 = s[6] ? v6_99 : {WIDTH{1'b0}};
  assign v5_50 = s[6] ? v6_101 : {WIDTH{1'b0}};
  assign v5_51 = s[6] ? v6_103 : {WIDTH{1'b0}};
  assign v5_52 = s[6] ? v6_105 : {WIDTH{1'b0}};
  assign v5_53 = s[6] ? v6_107 : {WIDTH{1'b0}};
  assign v5_54 = s[6] ? v6_109 : {WIDTH{1'b0}};
  assign v5_55 = s[6] ? v6_111 : {WIDTH{1'b0}};
  assign v5_56 = s[6] ? v6_113 : {WIDTH{1'b0}};
  assign v5_57 = s[6] ? v6_115 : {WIDTH{1'b0}};
  assign v5_58 = s[6] ? v6_117 : {WIDTH{1'b0}};
  assign v5_59 = s[6] ? v6_119 : {WIDTH{1'b0}};
  assign v5_60 = s[6] ? v6_121 : {WIDTH{1'b0}};
  assign v5_61 = s[6] ? v6_123 : {WIDTH{1'b0}};
  assign v5_62 = s[6] ? v6_125 : {WIDTH{1'b0}};
  assign v5_63 = s[6] ? v6_127 : {WIDTH{1'b0}};

  assign v6_0 = {WIDTH{1'b0}};
  assign v6_1 = {WIDTH{1'b0}};
  assign v6_2 = {WIDTH{1'b0}};
  assign v6_3 = {WIDTH{1'b0}};
  assign v6_4 = {WIDTH{1'b0}};
  assign v6_5 = {WIDTH{1'b0}};
  assign v6_6 = {WIDTH{1'b0}};
  assign v6_7 = {WIDTH{1'b0}};
  assign v6_8 = {WIDTH{1'b0}};
  assign v6_9 = {WIDTH{1'b0}};
  assign v6_10 = {WIDTH{1'b0}};
  assign v6_11 = {WIDTH{1'b0}};
  assign v6_12 = {WIDTH{1'b0}};
  assign v6_13 = {WIDTH{1'b0}};
  assign v6_14 = {WIDTH{1'b0}};
  assign v6_15 = {WIDTH{1'b0}};
  assign v6_16 = {WIDTH{1'b0}};
  assign v6_17 = {WIDTH{1'b0}};
  assign v6_18 = {WIDTH{1'b0}};
  assign v6_19 = {WIDTH{1'b0}};
  assign v6_20 = {WIDTH{1'b0}};
  assign v6_21 = {WIDTH{1'b0}};
  assign v6_22 = {WIDTH{1'b0}};
  assign v6_23 = {WIDTH{1'b0}};
  assign v6_24 = {WIDTH{1'b0}};
  assign v6_25 = {WIDTH{1'b0}};
  assign v6_26 = {WIDTH{1'b0}};
  assign v6_27 = {WIDTH{1'b0}};
  assign v6_28 = {WIDTH{1'b0}};
  assign v6_29 = {WIDTH{1'b0}};
  assign v6_30 = {WIDTH{1'b0}};
  assign v6_31 = {WIDTH{1'b0}};
  assign v6_32 = {WIDTH{1'b0}};
  assign v6_33 = {WIDTH{1'b0}};
  assign v6_34 = {WIDTH{1'b0}};
  assign v6_35 = {WIDTH{1'b0}};
  assign v6_36 = {WIDTH{1'b0}};
  assign v6_37 = {WIDTH{1'b0}};
  assign v6_38 = {WIDTH{1'b0}};
  assign v6_39 = {WIDTH{1'b0}};
  assign v6_40 = {WIDTH{1'b0}};
  assign v6_41 = {WIDTH{1'b0}};
  assign v6_42 = {WIDTH{1'b0}};
  assign v6_43 = {WIDTH{1'b0}};
  assign v6_44 = {WIDTH{1'b0}};
  assign v6_45 = {WIDTH{1'b0}};
  assign v6_46 = {WIDTH{1'b0}};
  assign v6_47 = {WIDTH{1'b0}};
  assign v6_48 = {WIDTH{1'b0}};
  assign v6_49 = {WIDTH{1'b0}};
  assign v6_50 = {WIDTH{1'b0}};
  assign v6_51 = {WIDTH{1'b0}};
  assign v6_52 = {WIDTH{1'b0}};
  assign v6_53 = {WIDTH{1'b0}};
  assign v6_54 = {WIDTH{1'b0}};
  assign v6_55 = {WIDTH{1'b0}};
  assign v6_56 = {WIDTH{1'b0}};
  assign v6_57 = {WIDTH{1'b0}};
  assign v6_58 = {WIDTH{1'b0}};
  assign v6_59 = {WIDTH{1'b0}};
  assign v6_60 = {WIDTH{1'b0}};
  assign v6_61 = {WIDTH{1'b0}};
  assign v6_62 = {WIDTH{1'b0}};
  assign v6_63 = {WIDTH{1'b0}};
  assign v6_64 = {WIDTH{1'b0}};
  assign v6_65 = {WIDTH{1'b0}};
  assign v6_66 = {WIDTH{1'b0}};
  assign v6_67 = {WIDTH{1'b0}};
  assign v6_68 = {WIDTH{1'b0}};
  assign v6_69 = {WIDTH{1'b0}};
  assign v6_70 = {WIDTH{1'b0}};
  assign v6_71 = s[7] ? d : {WIDTH{1'b0}};
  assign v6_72 = {WIDTH{1'b0}};
  assign v6_73 = {WIDTH{1'b0}};
  assign v6_74 = {WIDTH{1'b0}};
  assign v6_75 = {WIDTH{1'b0}};
  assign v6_76 = {WIDTH{1'b0}};
  assign v6_77 = {WIDTH{1'b0}};
  assign v6_78 = {WIDTH{1'b0}};
  assign v6_79 = {WIDTH{1'b0}};
  assign v6_80 = {WIDTH{1'b0}};
  assign v6_81 = {WIDTH{1'b0}};
  assign v6_82 = {WIDTH{1'b0}};
  assign v6_83 = {WIDTH{1'b0}};
  assign v6_84 = {WIDTH{1'b0}};
  assign v6_85 = {WIDTH{1'b0}};
  assign v6_86 = {WIDTH{1'b0}};
  assign v6_87 = {WIDTH{1'b0}};
  assign v6_88 = {WIDTH{1'b0}};
  assign v6_89 = {WIDTH{1'b0}};
  assign v6_90 = {WIDTH{1'b0}};
  assign v6_91 = {WIDTH{1'b0}};
  assign v6_92 = {WIDTH{1'b0}};
  assign v6_93 = {WIDTH{1'b0}};
  assign v6_94 = {WIDTH{1'b0}};
  assign v6_95 = {WIDTH{1'b0}};
  assign v6_96 = {WIDTH{1'b0}};
  assign v6_97 = {WIDTH{1'b0}};
  assign v6_98 = {WIDTH{1'b0}};
  assign v6_99 = {WIDTH{1'b0}};
  assign v6_100 = {WIDTH{1'b0}};
  assign v6_101 = {WIDTH{1'b0}};
  assign v6_102 = {WIDTH{1'b0}};
  assign v6_103 = {WIDTH{1'b0}};
  assign v6_104 = {WIDTH{1'b0}};
  assign v6_105 = {WIDTH{1'b0}};
  assign v6_106 = {WIDTH{1'b0}};
  assign v6_107 = {WIDTH{1'b0}};
  assign v6_108 = {WIDTH{1'b0}};
  assign v6_109 = {WIDTH{1'b0}};
  assign v6_110 = {WIDTH{1'b0}};
  assign v6_111 = {WIDTH{1'b0}};
  assign v6_112 = {WIDTH{1'b0}};
  assign v6_113 = {WIDTH{1'b0}};
  assign v6_114 = {WIDTH{1'b0}};
  assign v6_115 = {WIDTH{1'b0}};
  assign v6_116 = {WIDTH{1'b0}};
  assign v6_117 = {WIDTH{1'b0}};
  assign v6_118 = {WIDTH{1'b0}};
  assign v6_119 = {WIDTH{1'b0}};
  assign v6_120 = {WIDTH{1'b0}};
  assign v6_121 = {WIDTH{1'b0}};
  assign v6_122 = {WIDTH{1'b0}};
  assign v6_123 = {WIDTH{1'b0}};
  assign v6_124 = {WIDTH{1'b0}};
  assign v6_125 = {WIDTH{1'b0}};
  assign v6_126 = {WIDTH{1'b0}};
  assign v6_127 = {WIDTH{1'b0}};

endmodule

