/* modified netlist. Source: module SkinnyTop in file ../CaseStudies/06_Skinny64_64_round_based_encryption/FPGA_based/SkinnyTop_synthesis.v */
/* clock gating is added to the circuit, the latency increased 1 time(s)  */

module SkinnyTop_GHPCLL_ClockGating_d1 (clk, rst, Plaintext_s0, Key_s0, Key_s1, Plaintext_s1, Fresh, done, Ciphertext_s0, Ciphertext_s1, Synch);
    input clk ;
    input rst ;
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [1023:0] Fresh ;
    output done ;
    output [63:0] Ciphertext_s0 ;
    output [63:0] Ciphertext_s1 ;
    output Synch ;
    wire \FSMReg/s_current_state_sliced_sliced_0_290 ;
    wire \FSMReg/s_current_state_sliced_sliced_sliced_0_291 ;
    wire \FSMReg/s_current_state_sliced_sliced_sliced_1_292 ;
    wire \FSMReg/s_current_state_sliced_3_293 ;
    wire \FSMReg/s_current_state_sliced_sliced_sliced_2_294 ;
    wire [5:0] \FSMUpdate ;
    wire \FSM<0>_inv ;
    wire \FSM<1>_inv ;
    wire \FSM<2>_inv ;
    wire \FSM<3>_inv ;
    wire \FSM<4>_inv ;
    wire \FSM<5>_inv ;
    wire N01 ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire [63:0] StateRegInput ;
    wire [63:0] \TweakeyGeneration/StateReg/s_current_state ;
    wire [0:0] \FSMReg/s_current_state ;
    wire [5:0] FSMSelected ;
    wire [63:0] SubCellOutput ;
    wire [63:0] \TweakeyGeneration/StateRegInput ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_699 ;
    wire new_AGEMA_signal_700 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_713 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_721 ;
    wire new_AGEMA_signal_722 ;
    wire new_AGEMA_signal_723 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_729 ;
    wire new_AGEMA_signal_730 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_739 ;
    wire new_AGEMA_signal_740 ;
    wire new_AGEMA_signal_745 ;
    wire new_AGEMA_signal_746 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_753 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_762 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_769 ;
    wire new_AGEMA_signal_770 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_801 ;
    wire new_AGEMA_signal_802 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_808 ;
    wire new_AGEMA_signal_810 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1128 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[1].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMReg/s_current_state [0]), .O (FSMSelected[1]) ) ;
    LUT2 #( .INIT ( 4'hE ) ) \FSMMUX/GEN[0].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMUpdate [0]), .O (FSMSelected[0]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[4].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMReg/s_current_state_sliced_sliced_sliced_1_292 ), .O (FSMSelected[4]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[2].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMUpdate [2]), .O (FSMSelected[2]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[3].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMReg/s_current_state_sliced_3_293 ), .O (FSMSelected[3]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[5].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMUpdate [5]), .O (FSMSelected[5]) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[0].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_805, \TweakeyGeneration/StateReg/s_current_state [32]}), .I2 ({Key_s1[0], Key_s0[0]}), .O ({new_AGEMA_signal_807, \TweakeyGeneration/StateRegInput [0]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[1].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_808, \TweakeyGeneration/StateReg/s_current_state [33]}), .I2 ({Key_s1[1], Key_s0[1]}), .O ({new_AGEMA_signal_810, \TweakeyGeneration/StateRegInput [1]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[2].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_811, \TweakeyGeneration/StateReg/s_current_state [34]}), .I2 ({Key_s1[2], Key_s0[2]}), .O ({new_AGEMA_signal_813, \TweakeyGeneration/StateRegInput [2]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[3].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_814, \TweakeyGeneration/StateReg/s_current_state [35]}), .I2 ({Key_s1[3], Key_s0[3]}), .O ({new_AGEMA_signal_816, \TweakeyGeneration/StateRegInput [3]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[4].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_817, \TweakeyGeneration/StateReg/s_current_state [36]}), .I2 ({Key_s1[4], Key_s0[4]}), .O ({new_AGEMA_signal_819, \TweakeyGeneration/StateRegInput [4]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[5].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_820, \TweakeyGeneration/StateReg/s_current_state [37]}), .I2 ({Key_s1[5], Key_s0[5]}), .O ({new_AGEMA_signal_822, \TweakeyGeneration/StateRegInput [5]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[6].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_823, \TweakeyGeneration/StateReg/s_current_state [38]}), .I2 ({Key_s1[6], Key_s0[6]}), .O ({new_AGEMA_signal_825, \TweakeyGeneration/StateRegInput [6]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[7].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_826, \TweakeyGeneration/StateReg/s_current_state [39]}), .I2 ({Key_s1[7], Key_s0[7]}), .O ({new_AGEMA_signal_828, \TweakeyGeneration/StateRegInput [7]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[8].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_829, \TweakeyGeneration/StateReg/s_current_state [40]}), .I2 ({Key_s1[8], Key_s0[8]}), .O ({new_AGEMA_signal_831, \TweakeyGeneration/StateRegInput [8]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[9].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_832, \TweakeyGeneration/StateReg/s_current_state [41]}), .I2 ({Key_s1[9], Key_s0[9]}), .O ({new_AGEMA_signal_834, \TweakeyGeneration/StateRegInput [9]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[10].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_835, \TweakeyGeneration/StateReg/s_current_state [42]}), .I2 ({Key_s1[10], Key_s0[10]}), .O ({new_AGEMA_signal_837, \TweakeyGeneration/StateRegInput [10]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[11].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_838, \TweakeyGeneration/StateReg/s_current_state [43]}), .I2 ({Key_s1[11], Key_s0[11]}), .O ({new_AGEMA_signal_840, \TweakeyGeneration/StateRegInput [11]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[12].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_841, \TweakeyGeneration/StateReg/s_current_state [44]}), .I2 ({Key_s1[12], Key_s0[12]}), .O ({new_AGEMA_signal_843, \TweakeyGeneration/StateRegInput [12]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[13].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_844, \TweakeyGeneration/StateReg/s_current_state [45]}), .I2 ({Key_s1[13], Key_s0[13]}), .O ({new_AGEMA_signal_846, \TweakeyGeneration/StateRegInput [13]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[14].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_847, \TweakeyGeneration/StateReg/s_current_state [46]}), .I2 ({Key_s1[14], Key_s0[14]}), .O ({new_AGEMA_signal_849, \TweakeyGeneration/StateRegInput [14]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[15].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_850, \TweakeyGeneration/StateReg/s_current_state [47]}), .I2 ({Key_s1[15], Key_s0[15]}), .O ({new_AGEMA_signal_852, \TweakeyGeneration/StateRegInput [15]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[16].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_853, \TweakeyGeneration/StateReg/s_current_state [48]}), .I2 ({Key_s1[16], Key_s0[16]}), .O ({new_AGEMA_signal_855, \TweakeyGeneration/StateRegInput [16]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[17].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_856, \TweakeyGeneration/StateReg/s_current_state [49]}), .I2 ({Key_s1[17], Key_s0[17]}), .O ({new_AGEMA_signal_858, \TweakeyGeneration/StateRegInput [17]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[18].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_859, \TweakeyGeneration/StateReg/s_current_state [50]}), .I2 ({Key_s1[18], Key_s0[18]}), .O ({new_AGEMA_signal_861, \TweakeyGeneration/StateRegInput [18]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[19].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_862, \TweakeyGeneration/StateReg/s_current_state [51]}), .I2 ({Key_s1[19], Key_s0[19]}), .O ({new_AGEMA_signal_864, \TweakeyGeneration/StateRegInput [19]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[20].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_865, \TweakeyGeneration/StateReg/s_current_state [52]}), .I2 ({Key_s1[20], Key_s0[20]}), .O ({new_AGEMA_signal_867, \TweakeyGeneration/StateRegInput [20]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[21].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_868, \TweakeyGeneration/StateReg/s_current_state [53]}), .I2 ({Key_s1[21], Key_s0[21]}), .O ({new_AGEMA_signal_870, \TweakeyGeneration/StateRegInput [21]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[22].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_871, \TweakeyGeneration/StateReg/s_current_state [54]}), .I2 ({Key_s1[22], Key_s0[22]}), .O ({new_AGEMA_signal_873, \TweakeyGeneration/StateRegInput [22]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[23].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_874, \TweakeyGeneration/StateReg/s_current_state [55]}), .I2 ({Key_s1[23], Key_s0[23]}), .O ({new_AGEMA_signal_876, \TweakeyGeneration/StateRegInput [23]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[24].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_877, \TweakeyGeneration/StateReg/s_current_state [56]}), .I2 ({Key_s1[24], Key_s0[24]}), .O ({new_AGEMA_signal_879, \TweakeyGeneration/StateRegInput [24]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[25].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_880, \TweakeyGeneration/StateReg/s_current_state [57]}), .I2 ({Key_s1[25], Key_s0[25]}), .O ({new_AGEMA_signal_882, \TweakeyGeneration/StateRegInput [25]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[26].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_883, \TweakeyGeneration/StateReg/s_current_state [58]}), .I2 ({Key_s1[26], Key_s0[26]}), .O ({new_AGEMA_signal_885, \TweakeyGeneration/StateRegInput [26]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[27].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_886, \TweakeyGeneration/StateReg/s_current_state [59]}), .I2 ({Key_s1[27], Key_s0[27]}), .O ({new_AGEMA_signal_888, \TweakeyGeneration/StateRegInput [27]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[28].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_889, \TweakeyGeneration/StateReg/s_current_state [60]}), .I2 ({Key_s1[28], Key_s0[28]}), .O ({new_AGEMA_signal_891, \TweakeyGeneration/StateRegInput [28]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[29].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_892, \TweakeyGeneration/StateReg/s_current_state [61]}), .I2 ({Key_s1[29], Key_s0[29]}), .O ({new_AGEMA_signal_894, \TweakeyGeneration/StateRegInput [29]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[30].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_895, \TweakeyGeneration/StateReg/s_current_state [62]}), .I2 ({Key_s1[30], Key_s0[30]}), .O ({new_AGEMA_signal_897, \TweakeyGeneration/StateRegInput [30]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[31].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_898, \TweakeyGeneration/StateReg/s_current_state [63]}), .I2 ({Key_s1[31], Key_s0[31]}), .O ({new_AGEMA_signal_900, \TweakeyGeneration/StateRegInput [31]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[32].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_901, \TweakeyGeneration/StateReg/s_current_state [16]}), .I2 ({Key_s1[32], Key_s0[32]}), .O ({new_AGEMA_signal_903, \TweakeyGeneration/StateRegInput [32]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[33].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_904, \TweakeyGeneration/StateReg/s_current_state [17]}), .I2 ({Key_s1[33], Key_s0[33]}), .O ({new_AGEMA_signal_906, \TweakeyGeneration/StateRegInput [33]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[34].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_907, \TweakeyGeneration/StateReg/s_current_state [18]}), .I2 ({Key_s1[34], Key_s0[34]}), .O ({new_AGEMA_signal_909, \TweakeyGeneration/StateRegInput [34]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[35].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_910, \TweakeyGeneration/StateReg/s_current_state [19]}), .I2 ({Key_s1[35], Key_s0[35]}), .O ({new_AGEMA_signal_912, \TweakeyGeneration/StateRegInput [35]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[36].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_913, \TweakeyGeneration/StateReg/s_current_state [12]}), .I2 ({Key_s1[36], Key_s0[36]}), .O ({new_AGEMA_signal_915, \TweakeyGeneration/StateRegInput [36]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[37].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_916, \TweakeyGeneration/StateReg/s_current_state [13]}), .I2 ({Key_s1[37], Key_s0[37]}), .O ({new_AGEMA_signal_918, \TweakeyGeneration/StateRegInput [37]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[38].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_919, \TweakeyGeneration/StateReg/s_current_state [14]}), .I2 ({Key_s1[38], Key_s0[38]}), .O ({new_AGEMA_signal_921, \TweakeyGeneration/StateRegInput [38]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[39].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_922, \TweakeyGeneration/StateReg/s_current_state [15]}), .I2 ({Key_s1[39], Key_s0[39]}), .O ({new_AGEMA_signal_924, \TweakeyGeneration/StateRegInput [39]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[40].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_925, \TweakeyGeneration/StateReg/s_current_state [4]}), .I2 ({Key_s1[40], Key_s0[40]}), .O ({new_AGEMA_signal_927, \TweakeyGeneration/StateRegInput [40]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[41].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_928, \TweakeyGeneration/StateReg/s_current_state [5]}), .I2 ({Key_s1[41], Key_s0[41]}), .O ({new_AGEMA_signal_930, \TweakeyGeneration/StateRegInput [41]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[42].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_931, \TweakeyGeneration/StateReg/s_current_state [6]}), .I2 ({Key_s1[42], Key_s0[42]}), .O ({new_AGEMA_signal_933, \TweakeyGeneration/StateRegInput [42]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[43].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_934, \TweakeyGeneration/StateReg/s_current_state [7]}), .I2 ({Key_s1[43], Key_s0[43]}), .O ({new_AGEMA_signal_936, \TweakeyGeneration/StateRegInput [43]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[44].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_937, \TweakeyGeneration/StateReg/s_current_state [20]}), .I2 ({Key_s1[44], Key_s0[44]}), .O ({new_AGEMA_signal_939, \TweakeyGeneration/StateRegInput [44]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[45].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_940, \TweakeyGeneration/StateReg/s_current_state [21]}), .I2 ({Key_s1[45], Key_s0[45]}), .O ({new_AGEMA_signal_942, \TweakeyGeneration/StateRegInput [45]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[46].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_943, \TweakeyGeneration/StateReg/s_current_state [22]}), .I2 ({Key_s1[46], Key_s0[46]}), .O ({new_AGEMA_signal_945, \TweakeyGeneration/StateRegInput [46]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[47].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_946, \TweakeyGeneration/StateReg/s_current_state [23]}), .I2 ({Key_s1[47], Key_s0[47]}), .O ({new_AGEMA_signal_948, \TweakeyGeneration/StateRegInput [47]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[48].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_949, \TweakeyGeneration/StateReg/s_current_state [8]}), .I2 ({Key_s1[48], Key_s0[48]}), .O ({new_AGEMA_signal_951, \TweakeyGeneration/StateRegInput [48]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[49].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_952, \TweakeyGeneration/StateReg/s_current_state [9]}), .I2 ({Key_s1[49], Key_s0[49]}), .O ({new_AGEMA_signal_954, \TweakeyGeneration/StateRegInput [49]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[50].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_955, \TweakeyGeneration/StateReg/s_current_state [10]}), .I2 ({Key_s1[50], Key_s0[50]}), .O ({new_AGEMA_signal_957, \TweakeyGeneration/StateRegInput [50]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[51].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_958, \TweakeyGeneration/StateReg/s_current_state [11]}), .I2 ({Key_s1[51], Key_s0[51]}), .O ({new_AGEMA_signal_960, \TweakeyGeneration/StateRegInput [51]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[52].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_961, \TweakeyGeneration/StateReg/s_current_state [28]}), .I2 ({Key_s1[52], Key_s0[52]}), .O ({new_AGEMA_signal_963, \TweakeyGeneration/StateRegInput [52]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[53].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_964, \TweakeyGeneration/StateReg/s_current_state [29]}), .I2 ({Key_s1[53], Key_s0[53]}), .O ({new_AGEMA_signal_966, \TweakeyGeneration/StateRegInput [53]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[54].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_967, \TweakeyGeneration/StateReg/s_current_state [30]}), .I2 ({Key_s1[54], Key_s0[54]}), .O ({new_AGEMA_signal_969, \TweakeyGeneration/StateRegInput [54]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[55].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_970, \TweakeyGeneration/StateReg/s_current_state [31]}), .I2 ({Key_s1[55], Key_s0[55]}), .O ({new_AGEMA_signal_972, \TweakeyGeneration/StateRegInput [55]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[56].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_973, \TweakeyGeneration/StateReg/s_current_state [0]}), .I2 ({Key_s1[56], Key_s0[56]}), .O ({new_AGEMA_signal_975, \TweakeyGeneration/StateRegInput [56]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[57].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_976, \TweakeyGeneration/StateReg/s_current_state [1]}), .I2 ({Key_s1[57], Key_s0[57]}), .O ({new_AGEMA_signal_978, \TweakeyGeneration/StateRegInput [57]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[58].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_979, \TweakeyGeneration/StateReg/s_current_state [2]}), .I2 ({Key_s1[58], Key_s0[58]}), .O ({new_AGEMA_signal_981, \TweakeyGeneration/StateRegInput [58]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[59].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_982, \TweakeyGeneration/StateReg/s_current_state [3]}), .I2 ({Key_s1[59], Key_s0[59]}), .O ({new_AGEMA_signal_984, \TweakeyGeneration/StateRegInput [59]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[60].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_985, \TweakeyGeneration/StateReg/s_current_state [24]}), .I2 ({Key_s1[60], Key_s0[60]}), .O ({new_AGEMA_signal_987, \TweakeyGeneration/StateRegInput [60]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[61].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_988, \TweakeyGeneration/StateReg/s_current_state [25]}), .I2 ({Key_s1[61], Key_s0[61]}), .O ({new_AGEMA_signal_990, \TweakeyGeneration/StateRegInput [61]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[62].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_991, \TweakeyGeneration/StateReg/s_current_state [26]}), .I2 ({Key_s1[62], Key_s0[62]}), .O ({new_AGEMA_signal_993, \TweakeyGeneration/StateRegInput [62]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \TweakeyGeneration/KEYMUX/GEN[63].MUXInst/Mmux_Q11 ( .I0 ({1'b0, rst}), .I1 ({new_AGEMA_signal_994, \TweakeyGeneration/StateReg/s_current_state [27]}), .I2 ({Key_s1[63], Key_s0[63]}), .O ({new_AGEMA_signal_996, \TweakeyGeneration/StateRegInput [63]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b10 ), .INIT2 ( 4'hA ) ) \StateRegInput<60>_SW0 ( .I0 ({new_AGEMA_signal_889, \TweakeyGeneration/StateReg/s_current_state [60]}), .I1 ({1'b0, \FSMReg/s_current_state [0]}), .O ({new_AGEMA_signal_997, N01}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b10 ), .INIT2 ( 4'hA ) ) \StateRegInput<61>_SW0 ( .I0 ({new_AGEMA_signal_892, \TweakeyGeneration/StateReg/s_current_state [61]}), .I1 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_2_294 }), .O ({new_AGEMA_signal_998, N2}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b10 ), .INIT2 ( 4'hA ) ) \StateRegInput<62>_SW0 ( .I0 ({new_AGEMA_signal_895, \TweakeyGeneration/StateReg/s_current_state [62]}), .I1 ({1'b0, \FSMReg/s_current_state_sliced_3_293 }), .O ({new_AGEMA_signal_999, N4}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b10 ), .INIT2 ( 4'hA ) ) \StateRegInput<63>_SW0 ( .I0 ({new_AGEMA_signal_898, \TweakeyGeneration/StateReg/s_current_state [63]}), .I1 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_1_292 }), .O ({new_AGEMA_signal_1000, N6}) ) ;
    INV \FSM<0>_inv1_INV_0 ( .I (\FSMReg/s_current_state [0]), .O (\FSM<0>_inv ) ) ;
    INV \FSM<1>_inv1_INV_0 ( .I (\FSMReg/s_current_state_sliced_sliced_sliced_2_294 ), .O (\FSM<1>_inv ) ) ;
    INV \FSM<2>_inv1_INV_0 ( .I (\FSMReg/s_current_state_sliced_3_293 ), .O (\FSM<2>_inv ) ) ;
    INV \FSM<3>_inv1_INV_0 ( .I (\FSMReg/s_current_state_sliced_sliced_sliced_1_292 ), .O (\FSM<3>_inv ) ) ;
    INV \FSM<4>_inv1_INV_0 ( .I (\FSMReg/s_current_state_sliced_sliced_sliced_0_291 ), .O (\FSM<4>_inv ) ) ;
    INV \FSM<5>_inv1_INV_0 ( .I (\FSMReg/s_current_state_sliced_sliced_0_290 ), .O (\FSM<5>_inv ) ) ;
    LUT6 #( .INIT ( 64'h0000000000004000 ) ) \FSMSignalsInst/doneInst/Mram_output11 ( .I0 (\FSM<0>_inv ), .I1 (\FSM<1>_inv ), .I2 (\FSM<2>_inv ), .I3 (\FSM<3>_inv ), .I4 (\FSM<4>_inv ), .I5 (\FSM<5>_inv ), .O (done) ) ;
    LUT6 #( .INIT ( 64'h5555555557555555 ) ) \FSMUpdateInst/GEN[5].StateUpdateInst/Mram_output11 ( .I0 (\FSM<4>_inv ), .I1 (\FSM<1>_inv ), .I2 (\FSM<5>_inv ), .I3 (\FSM<3>_inv ), .I4 (\FSM<2>_inv ), .I5 (\FSM<0>_inv ), .O (\FSMUpdate [5]) ) ;
    LUT6 #( .INIT ( 64'h5555551555555555 ) ) \FSMUpdateInst/GEN[2].StateUpdateInst/Mram_output11 ( .I0 (\FSM<1>_inv ), .I1 (\FSM<4>_inv ), .I2 (\FSM<3>_inv ), .I3 (\FSM<5>_inv ), .I4 (\FSM<0>_inv ), .I5 (\FSM<2>_inv ), .O (\FSMUpdate [2]) ) ;
    LUT6 #( .INIT ( 64'h999D999999999999 ) ) \FSMUpdateInst/GEN[0].StateUpdateInst/Mram_output11 ( .I0 (\FSM<5>_inv ), .I1 (\FSM<4>_inv ), .I2 (\FSM<0>_inv ), .I3 (\FSM<1>_inv ), .I4 (\FSM<2>_inv ), .I5 (\FSM<3>_inv ), .O (\FSMUpdate [0]) ) ;
    ClockGatingController #(2) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[0].SboxInst/y_0 ( .I0 ({Ciphertext_s1[0], Ciphertext_s0[0]}), .I1 ({Ciphertext_s1[1], Ciphertext_s0[1]}), .I2 ({Ciphertext_s1[2], Ciphertext_s0[2]}), .I3 ({Ciphertext_s1[3], Ciphertext_s0[3]}), .clk (clk), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .O ({new_AGEMA_signal_681, SubCellOutput[0]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[0].SboxInst/y_1 ( .I0 ({Ciphertext_s1[0], Ciphertext_s0[0]}), .I1 ({Ciphertext_s1[1], Ciphertext_s0[1]}), .I2 ({Ciphertext_s1[2], Ciphertext_s0[2]}), .I3 ({Ciphertext_s1[3], Ciphertext_s0[3]}), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .O ({new_AGEMA_signal_682, SubCellOutput[1]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[0].SboxInst/y_2 ( .I0 ({Ciphertext_s1[0], Ciphertext_s0[0]}), .I1 ({Ciphertext_s1[1], Ciphertext_s0[1]}), .I2 ({Ciphertext_s1[2], Ciphertext_s0[2]}), .I3 ({Ciphertext_s1[3], Ciphertext_s0[3]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .O ({new_AGEMA_signal_683, SubCellOutput[2]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[0].SboxInst/y_3 ( .I0 ({Ciphertext_s1[0], Ciphertext_s0[0]}), .I1 ({Ciphertext_s1[1], Ciphertext_s0[1]}), .I2 ({Ciphertext_s1[2], Ciphertext_s0[2]}), .I3 ({Ciphertext_s1[3], Ciphertext_s0[3]}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .O ({new_AGEMA_signal_684, SubCellOutput[3]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[1].SboxInst/y_0 ( .I0 ({Ciphertext_s1[4], Ciphertext_s0[4]}), .I1 ({Ciphertext_s1[5], Ciphertext_s0[5]}), .I2 ({Ciphertext_s1[6], Ciphertext_s0[6]}), .I3 ({Ciphertext_s1[7], Ciphertext_s0[7]}), .clk (clk), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .O ({new_AGEMA_signal_689, SubCellOutput[4]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[1].SboxInst/y_1 ( .I0 ({Ciphertext_s1[4], Ciphertext_s0[4]}), .I1 ({Ciphertext_s1[5], Ciphertext_s0[5]}), .I2 ({Ciphertext_s1[6], Ciphertext_s0[6]}), .I3 ({Ciphertext_s1[7], Ciphertext_s0[7]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .O ({new_AGEMA_signal_690, SubCellOutput[5]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[1].SboxInst/y_2 ( .I0 ({Ciphertext_s1[4], Ciphertext_s0[4]}), .I1 ({Ciphertext_s1[5], Ciphertext_s0[5]}), .I2 ({Ciphertext_s1[6], Ciphertext_s0[6]}), .I3 ({Ciphertext_s1[7], Ciphertext_s0[7]}), .clk (clk), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .O ({new_AGEMA_signal_691, SubCellOutput[6]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[1].SboxInst/y_3 ( .I0 ({Ciphertext_s1[4], Ciphertext_s0[4]}), .I1 ({Ciphertext_s1[5], Ciphertext_s0[5]}), .I2 ({Ciphertext_s1[6], Ciphertext_s0[6]}), .I3 ({Ciphertext_s1[7], Ciphertext_s0[7]}), .clk (clk), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .O ({new_AGEMA_signal_692, SubCellOutput[7]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[2].SboxInst/y_0 ( .I0 ({Ciphertext_s1[8], Ciphertext_s0[8]}), .I1 ({Ciphertext_s1[9], Ciphertext_s0[9]}), .I2 ({Ciphertext_s1[10], Ciphertext_s0[10]}), .I3 ({Ciphertext_s1[11], Ciphertext_s0[11]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .O ({new_AGEMA_signal_697, SubCellOutput[8]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[2].SboxInst/y_1 ( .I0 ({Ciphertext_s1[8], Ciphertext_s0[8]}), .I1 ({Ciphertext_s1[9], Ciphertext_s0[9]}), .I2 ({Ciphertext_s1[10], Ciphertext_s0[10]}), .I3 ({Ciphertext_s1[11], Ciphertext_s0[11]}), .clk (clk), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .O ({new_AGEMA_signal_698, SubCellOutput[9]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[2].SboxInst/y_2 ( .I0 ({Ciphertext_s1[8], Ciphertext_s0[8]}), .I1 ({Ciphertext_s1[9], Ciphertext_s0[9]}), .I2 ({Ciphertext_s1[10], Ciphertext_s0[10]}), .I3 ({Ciphertext_s1[11], Ciphertext_s0[11]}), .clk (clk), .r ({Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .O ({new_AGEMA_signal_699, SubCellOutput[10]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[2].SboxInst/y_3 ( .I0 ({Ciphertext_s1[8], Ciphertext_s0[8]}), .I1 ({Ciphertext_s1[9], Ciphertext_s0[9]}), .I2 ({Ciphertext_s1[10], Ciphertext_s0[10]}), .I3 ({Ciphertext_s1[11], Ciphertext_s0[11]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176]}), .O ({new_AGEMA_signal_700, SubCellOutput[11]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[3].SboxInst/y_0 ( .I0 ({Ciphertext_s1[12], Ciphertext_s0[12]}), .I1 ({Ciphertext_s1[13], Ciphertext_s0[13]}), .I2 ({Ciphertext_s1[14], Ciphertext_s0[14]}), .I3 ({Ciphertext_s1[15], Ciphertext_s0[15]}), .clk (clk), .r ({Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .O ({new_AGEMA_signal_705, SubCellOutput[12]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[3].SboxInst/y_1 ( .I0 ({Ciphertext_s1[12], Ciphertext_s0[12]}), .I1 ({Ciphertext_s1[13], Ciphertext_s0[13]}), .I2 ({Ciphertext_s1[14], Ciphertext_s0[14]}), .I3 ({Ciphertext_s1[15], Ciphertext_s0[15]}), .clk (clk), .r ({Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208]}), .O ({new_AGEMA_signal_706, SubCellOutput[13]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[3].SboxInst/y_2 ( .I0 ({Ciphertext_s1[12], Ciphertext_s0[12]}), .I1 ({Ciphertext_s1[13], Ciphertext_s0[13]}), .I2 ({Ciphertext_s1[14], Ciphertext_s0[14]}), .I3 ({Ciphertext_s1[15], Ciphertext_s0[15]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224]}), .O ({new_AGEMA_signal_707, SubCellOutput[14]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[3].SboxInst/y_3 ( .I0 ({Ciphertext_s1[12], Ciphertext_s0[12]}), .I1 ({Ciphertext_s1[13], Ciphertext_s0[13]}), .I2 ({Ciphertext_s1[14], Ciphertext_s0[14]}), .I3 ({Ciphertext_s1[15], Ciphertext_s0[15]}), .clk (clk), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .O ({new_AGEMA_signal_708, SubCellOutput[15]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[4].SboxInst/y_0 ( .I0 ({Ciphertext_s1[16], Ciphertext_s0[16]}), .I1 ({Ciphertext_s1[17], Ciphertext_s0[17]}), .I2 ({Ciphertext_s1[18], Ciphertext_s0[18]}), .I3 ({Ciphertext_s1[19], Ciphertext_s0[19]}), .clk (clk), .r ({Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .O ({new_AGEMA_signal_713, SubCellOutput[16]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[4].SboxInst/y_1 ( .I0 ({Ciphertext_s1[16], Ciphertext_s0[16]}), .I1 ({Ciphertext_s1[17], Ciphertext_s0[17]}), .I2 ({Ciphertext_s1[18], Ciphertext_s0[18]}), .I3 ({Ciphertext_s1[19], Ciphertext_s0[19]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272]}), .O ({new_AGEMA_signal_714, SubCellOutput[17]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[4].SboxInst/y_2 ( .I0 ({Ciphertext_s1[16], Ciphertext_s0[16]}), .I1 ({Ciphertext_s1[17], Ciphertext_s0[17]}), .I2 ({Ciphertext_s1[18], Ciphertext_s0[18]}), .I3 ({Ciphertext_s1[19], Ciphertext_s0[19]}), .clk (clk), .r ({Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .O ({new_AGEMA_signal_715, SubCellOutput[18]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[4].SboxInst/y_3 ( .I0 ({Ciphertext_s1[16], Ciphertext_s0[16]}), .I1 ({Ciphertext_s1[17], Ciphertext_s0[17]}), .I2 ({Ciphertext_s1[18], Ciphertext_s0[18]}), .I3 ({Ciphertext_s1[19], Ciphertext_s0[19]}), .clk (clk), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304]}), .O ({new_AGEMA_signal_716, SubCellOutput[19]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[5].SboxInst/y_0 ( .I0 ({Ciphertext_s1[20], Ciphertext_s0[20]}), .I1 ({Ciphertext_s1[21], Ciphertext_s0[21]}), .I2 ({Ciphertext_s1[22], Ciphertext_s0[22]}), .I3 ({Ciphertext_s1[23], Ciphertext_s0[23]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .O ({new_AGEMA_signal_721, SubCellOutput[20]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[5].SboxInst/y_1 ( .I0 ({Ciphertext_s1[20], Ciphertext_s0[20]}), .I1 ({Ciphertext_s1[21], Ciphertext_s0[21]}), .I2 ({Ciphertext_s1[22], Ciphertext_s0[22]}), .I3 ({Ciphertext_s1[23], Ciphertext_s0[23]}), .clk (clk), .r ({Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .O ({new_AGEMA_signal_722, SubCellOutput[21]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[5].SboxInst/y_2 ( .I0 ({Ciphertext_s1[20], Ciphertext_s0[20]}), .I1 ({Ciphertext_s1[21], Ciphertext_s0[21]}), .I2 ({Ciphertext_s1[22], Ciphertext_s0[22]}), .I3 ({Ciphertext_s1[23], Ciphertext_s0[23]}), .clk (clk), .r ({Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352]}), .O ({new_AGEMA_signal_723, SubCellOutput[22]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[5].SboxInst/y_3 ( .I0 ({Ciphertext_s1[20], Ciphertext_s0[20]}), .I1 ({Ciphertext_s1[21], Ciphertext_s0[21]}), .I2 ({Ciphertext_s1[22], Ciphertext_s0[22]}), .I3 ({Ciphertext_s1[23], Ciphertext_s0[23]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368]}), .O ({new_AGEMA_signal_724, SubCellOutput[23]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[6].SboxInst/y_0 ( .I0 ({Ciphertext_s1[24], Ciphertext_s0[24]}), .I1 ({Ciphertext_s1[25], Ciphertext_s0[25]}), .I2 ({Ciphertext_s1[26], Ciphertext_s0[26]}), .I3 ({Ciphertext_s1[27], Ciphertext_s0[27]}), .clk (clk), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .O ({new_AGEMA_signal_729, SubCellOutput[24]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[6].SboxInst/y_1 ( .I0 ({Ciphertext_s1[24], Ciphertext_s0[24]}), .I1 ({Ciphertext_s1[25], Ciphertext_s0[25]}), .I2 ({Ciphertext_s1[26], Ciphertext_s0[26]}), .I3 ({Ciphertext_s1[27], Ciphertext_s0[27]}), .clk (clk), .r ({Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .O ({new_AGEMA_signal_730, SubCellOutput[25]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[6].SboxInst/y_2 ( .I0 ({Ciphertext_s1[24], Ciphertext_s0[24]}), .I1 ({Ciphertext_s1[25], Ciphertext_s0[25]}), .I2 ({Ciphertext_s1[26], Ciphertext_s0[26]}), .I3 ({Ciphertext_s1[27], Ciphertext_s0[27]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416]}), .O ({new_AGEMA_signal_731, SubCellOutput[26]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[6].SboxInst/y_3 ( .I0 ({Ciphertext_s1[24], Ciphertext_s0[24]}), .I1 ({Ciphertext_s1[25], Ciphertext_s0[25]}), .I2 ({Ciphertext_s1[26], Ciphertext_s0[26]}), .I3 ({Ciphertext_s1[27], Ciphertext_s0[27]}), .clk (clk), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .O ({new_AGEMA_signal_732, SubCellOutput[27]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[7].SboxInst/y_0 ( .I0 ({Ciphertext_s1[28], Ciphertext_s0[28]}), .I1 ({Ciphertext_s1[29], Ciphertext_s0[29]}), .I2 ({Ciphertext_s1[30], Ciphertext_s0[30]}), .I3 ({Ciphertext_s1[31], Ciphertext_s0[31]}), .clk (clk), .r ({Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .O ({new_AGEMA_signal_737, SubCellOutput[28]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[7].SboxInst/y_1 ( .I0 ({Ciphertext_s1[28], Ciphertext_s0[28]}), .I1 ({Ciphertext_s1[29], Ciphertext_s0[29]}), .I2 ({Ciphertext_s1[30], Ciphertext_s0[30]}), .I3 ({Ciphertext_s1[31], Ciphertext_s0[31]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464]}), .O ({new_AGEMA_signal_738, SubCellOutput[29]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[7].SboxInst/y_2 ( .I0 ({Ciphertext_s1[28], Ciphertext_s0[28]}), .I1 ({Ciphertext_s1[29], Ciphertext_s0[29]}), .I2 ({Ciphertext_s1[30], Ciphertext_s0[30]}), .I3 ({Ciphertext_s1[31], Ciphertext_s0[31]}), .clk (clk), .r ({Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .O ({new_AGEMA_signal_739, SubCellOutput[30]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[7].SboxInst/y_3 ( .I0 ({Ciphertext_s1[28], Ciphertext_s0[28]}), .I1 ({Ciphertext_s1[29], Ciphertext_s0[29]}), .I2 ({Ciphertext_s1[30], Ciphertext_s0[30]}), .I3 ({Ciphertext_s1[31], Ciphertext_s0[31]}), .clk (clk), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496]}), .O ({new_AGEMA_signal_740, SubCellOutput[31]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[8].SboxInst/y_0 ( .I0 ({Ciphertext_s1[32], Ciphertext_s0[32]}), .I1 ({Ciphertext_s1[33], Ciphertext_s0[33]}), .I2 ({Ciphertext_s1[34], Ciphertext_s0[34]}), .I3 ({Ciphertext_s1[35], Ciphertext_s0[35]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .O ({new_AGEMA_signal_745, SubCellOutput[32]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[8].SboxInst/y_1 ( .I0 ({Ciphertext_s1[32], Ciphertext_s0[32]}), .I1 ({Ciphertext_s1[33], Ciphertext_s0[33]}), .I2 ({Ciphertext_s1[34], Ciphertext_s0[34]}), .I3 ({Ciphertext_s1[35], Ciphertext_s0[35]}), .clk (clk), .r ({Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .O ({new_AGEMA_signal_746, SubCellOutput[33]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[8].SboxInst/y_2 ( .I0 ({Ciphertext_s1[32], Ciphertext_s0[32]}), .I1 ({Ciphertext_s1[33], Ciphertext_s0[33]}), .I2 ({Ciphertext_s1[34], Ciphertext_s0[34]}), .I3 ({Ciphertext_s1[35], Ciphertext_s0[35]}), .clk (clk), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544]}), .O ({new_AGEMA_signal_747, SubCellOutput[34]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[8].SboxInst/y_3 ( .I0 ({Ciphertext_s1[32], Ciphertext_s0[32]}), .I1 ({Ciphertext_s1[33], Ciphertext_s0[33]}), .I2 ({Ciphertext_s1[34], Ciphertext_s0[34]}), .I3 ({Ciphertext_s1[35], Ciphertext_s0[35]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .O ({new_AGEMA_signal_748, SubCellOutput[35]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[9].SboxInst/y_0 ( .I0 ({Ciphertext_s1[36], Ciphertext_s0[36]}), .I1 ({Ciphertext_s1[37], Ciphertext_s0[37]}), .I2 ({Ciphertext_s1[38], Ciphertext_s0[38]}), .I3 ({Ciphertext_s1[39], Ciphertext_s0[39]}), .clk (clk), .r ({Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .O ({new_AGEMA_signal_753, SubCellOutput[36]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[9].SboxInst/y_1 ( .I0 ({Ciphertext_s1[36], Ciphertext_s0[36]}), .I1 ({Ciphertext_s1[37], Ciphertext_s0[37]}), .I2 ({Ciphertext_s1[38], Ciphertext_s0[38]}), .I3 ({Ciphertext_s1[39], Ciphertext_s0[39]}), .clk (clk), .r ({Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592]}), .O ({new_AGEMA_signal_754, SubCellOutput[37]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[9].SboxInst/y_2 ( .I0 ({Ciphertext_s1[36], Ciphertext_s0[36]}), .I1 ({Ciphertext_s1[37], Ciphertext_s0[37]}), .I2 ({Ciphertext_s1[38], Ciphertext_s0[38]}), .I3 ({Ciphertext_s1[39], Ciphertext_s0[39]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608]}), .O ({new_AGEMA_signal_755, SubCellOutput[38]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[9].SboxInst/y_3 ( .I0 ({Ciphertext_s1[36], Ciphertext_s0[36]}), .I1 ({Ciphertext_s1[37], Ciphertext_s0[37]}), .I2 ({Ciphertext_s1[38], Ciphertext_s0[38]}), .I3 ({Ciphertext_s1[39], Ciphertext_s0[39]}), .clk (clk), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .O ({new_AGEMA_signal_756, SubCellOutput[39]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[10].SboxInst/y_0 ( .I0 ({Ciphertext_s1[40], Ciphertext_s0[40]}), .I1 ({Ciphertext_s1[41], Ciphertext_s0[41]}), .I2 ({Ciphertext_s1[42], Ciphertext_s0[42]}), .I3 ({Ciphertext_s1[43], Ciphertext_s0[43]}), .clk (clk), .r ({Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .O ({new_AGEMA_signal_761, SubCellOutput[40]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[10].SboxInst/y_1 ( .I0 ({Ciphertext_s1[40], Ciphertext_s0[40]}), .I1 ({Ciphertext_s1[41], Ciphertext_s0[41]}), .I2 ({Ciphertext_s1[42], Ciphertext_s0[42]}), .I3 ({Ciphertext_s1[43], Ciphertext_s0[43]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656]}), .O ({new_AGEMA_signal_762, SubCellOutput[41]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[10].SboxInst/y_2 ( .I0 ({Ciphertext_s1[40], Ciphertext_s0[40]}), .I1 ({Ciphertext_s1[41], Ciphertext_s0[41]}), .I2 ({Ciphertext_s1[42], Ciphertext_s0[42]}), .I3 ({Ciphertext_s1[43], Ciphertext_s0[43]}), .clk (clk), .r ({Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .O ({new_AGEMA_signal_763, SubCellOutput[42]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[10].SboxInst/y_3 ( .I0 ({Ciphertext_s1[40], Ciphertext_s0[40]}), .I1 ({Ciphertext_s1[41], Ciphertext_s0[41]}), .I2 ({Ciphertext_s1[42], Ciphertext_s0[42]}), .I3 ({Ciphertext_s1[43], Ciphertext_s0[43]}), .clk (clk), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688]}), .O ({new_AGEMA_signal_764, SubCellOutput[43]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[11].SboxInst/y_0 ( .I0 ({Ciphertext_s1[44], Ciphertext_s0[44]}), .I1 ({Ciphertext_s1[45], Ciphertext_s0[45]}), .I2 ({Ciphertext_s1[46], Ciphertext_s0[46]}), .I3 ({Ciphertext_s1[47], Ciphertext_s0[47]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .O ({new_AGEMA_signal_769, SubCellOutput[44]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[11].SboxInst/y_1 ( .I0 ({Ciphertext_s1[44], Ciphertext_s0[44]}), .I1 ({Ciphertext_s1[45], Ciphertext_s0[45]}), .I2 ({Ciphertext_s1[46], Ciphertext_s0[46]}), .I3 ({Ciphertext_s1[47], Ciphertext_s0[47]}), .clk (clk), .r ({Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .O ({new_AGEMA_signal_770, SubCellOutput[45]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[11].SboxInst/y_2 ( .I0 ({Ciphertext_s1[44], Ciphertext_s0[44]}), .I1 ({Ciphertext_s1[45], Ciphertext_s0[45]}), .I2 ({Ciphertext_s1[46], Ciphertext_s0[46]}), .I3 ({Ciphertext_s1[47], Ciphertext_s0[47]}), .clk (clk), .r ({Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736]}), .O ({new_AGEMA_signal_771, SubCellOutput[46]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[11].SboxInst/y_3 ( .I0 ({Ciphertext_s1[44], Ciphertext_s0[44]}), .I1 ({Ciphertext_s1[45], Ciphertext_s0[45]}), .I2 ({Ciphertext_s1[46], Ciphertext_s0[46]}), .I3 ({Ciphertext_s1[47], Ciphertext_s0[47]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752]}), .O ({new_AGEMA_signal_772, SubCellOutput[47]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[12].SboxInst/y_0 ( .I0 ({Ciphertext_s1[48], Ciphertext_s0[48]}), .I1 ({Ciphertext_s1[49], Ciphertext_s0[49]}), .I2 ({Ciphertext_s1[50], Ciphertext_s0[50]}), .I3 ({Ciphertext_s1[51], Ciphertext_s0[51]}), .clk (clk), .r ({Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .O ({new_AGEMA_signal_777, SubCellOutput[48]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[12].SboxInst/y_1 ( .I0 ({Ciphertext_s1[48], Ciphertext_s0[48]}), .I1 ({Ciphertext_s1[49], Ciphertext_s0[49]}), .I2 ({Ciphertext_s1[50], Ciphertext_s0[50]}), .I3 ({Ciphertext_s1[51], Ciphertext_s0[51]}), .clk (clk), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784]}), .O ({new_AGEMA_signal_778, SubCellOutput[49]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[12].SboxInst/y_2 ( .I0 ({Ciphertext_s1[48], Ciphertext_s0[48]}), .I1 ({Ciphertext_s1[49], Ciphertext_s0[49]}), .I2 ({Ciphertext_s1[50], Ciphertext_s0[50]}), .I3 ({Ciphertext_s1[51], Ciphertext_s0[51]}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .O ({new_AGEMA_signal_779, SubCellOutput[50]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[12].SboxInst/y_3 ( .I0 ({Ciphertext_s1[48], Ciphertext_s0[48]}), .I1 ({Ciphertext_s1[49], Ciphertext_s0[49]}), .I2 ({Ciphertext_s1[50], Ciphertext_s0[50]}), .I3 ({Ciphertext_s1[51], Ciphertext_s0[51]}), .clk (clk), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .O ({new_AGEMA_signal_780, SubCellOutput[51]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[13].SboxInst/y_0 ( .I0 ({Ciphertext_s1[52], Ciphertext_s0[52]}), .I1 ({Ciphertext_s1[53], Ciphertext_s0[53]}), .I2 ({Ciphertext_s1[54], Ciphertext_s0[54]}), .I3 ({Ciphertext_s1[55], Ciphertext_s0[55]}), .clk (clk), .r ({Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .O ({new_AGEMA_signal_785, SubCellOutput[52]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[13].SboxInst/y_1 ( .I0 ({Ciphertext_s1[52], Ciphertext_s0[52]}), .I1 ({Ciphertext_s1[53], Ciphertext_s0[53]}), .I2 ({Ciphertext_s1[54], Ciphertext_s0[54]}), .I3 ({Ciphertext_s1[55], Ciphertext_s0[55]}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848]}), .O ({new_AGEMA_signal_786, SubCellOutput[53]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[13].SboxInst/y_2 ( .I0 ({Ciphertext_s1[52], Ciphertext_s0[52]}), .I1 ({Ciphertext_s1[53], Ciphertext_s0[53]}), .I2 ({Ciphertext_s1[54], Ciphertext_s0[54]}), .I3 ({Ciphertext_s1[55], Ciphertext_s0[55]}), .clk (clk), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .O ({new_AGEMA_signal_787, SubCellOutput[54]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[13].SboxInst/y_3 ( .I0 ({Ciphertext_s1[52], Ciphertext_s0[52]}), .I1 ({Ciphertext_s1[53], Ciphertext_s0[53]}), .I2 ({Ciphertext_s1[54], Ciphertext_s0[54]}), .I3 ({Ciphertext_s1[55], Ciphertext_s0[55]}), .clk (clk), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .O ({new_AGEMA_signal_788, SubCellOutput[55]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[14].SboxInst/y_0 ( .I0 ({Ciphertext_s1[56], Ciphertext_s0[56]}), .I1 ({Ciphertext_s1[57], Ciphertext_s0[57]}), .I2 ({Ciphertext_s1[58], Ciphertext_s0[58]}), .I3 ({Ciphertext_s1[59], Ciphertext_s0[59]}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .O ({new_AGEMA_signal_793, SubCellOutput[56]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[14].SboxInst/y_1 ( .I0 ({Ciphertext_s1[56], Ciphertext_s0[56]}), .I1 ({Ciphertext_s1[57], Ciphertext_s0[57]}), .I2 ({Ciphertext_s1[58], Ciphertext_s0[58]}), .I3 ({Ciphertext_s1[59], Ciphertext_s0[59]}), .clk (clk), .r ({Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .O ({new_AGEMA_signal_794, SubCellOutput[57]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[14].SboxInst/y_2 ( .I0 ({Ciphertext_s1[56], Ciphertext_s0[56]}), .I1 ({Ciphertext_s1[57], Ciphertext_s0[57]}), .I2 ({Ciphertext_s1[58], Ciphertext_s0[58]}), .I3 ({Ciphertext_s1[59], Ciphertext_s0[59]}), .clk (clk), .r ({Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928]}), .O ({new_AGEMA_signal_795, SubCellOutput[58]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[14].SboxInst/y_3 ( .I0 ({Ciphertext_s1[56], Ciphertext_s0[56]}), .I1 ({Ciphertext_s1[57], Ciphertext_s0[57]}), .I2 ({Ciphertext_s1[58], Ciphertext_s0[58]}), .I3 ({Ciphertext_s1[59], Ciphertext_s0[59]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944]}), .O ({new_AGEMA_signal_796, SubCellOutput[59]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hCD94 ) ) \SubCellInst/GEN[15].SboxInst/y_0 ( .I0 ({Ciphertext_s1[60], Ciphertext_s0[60]}), .I1 ({Ciphertext_s1[61], Ciphertext_s0[61]}), .I2 ({Ciphertext_s1[62], Ciphertext_s0[62]}), .I3 ({Ciphertext_s1[63], Ciphertext_s0[63]}), .clk (clk), .r ({Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .O ({new_AGEMA_signal_801, SubCellOutput[60]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hE1E2 ) ) \SubCellInst/GEN[15].SboxInst/y_1 ( .I0 ({Ciphertext_s1[60], Ciphertext_s0[60]}), .I1 ({Ciphertext_s1[61], Ciphertext_s0[61]}), .I2 ({Ciphertext_s1[62], Ciphertext_s0[62]}), .I3 ({Ciphertext_s1[63], Ciphertext_s0[63]}), .clk (clk), .r ({Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976]}), .O ({new_AGEMA_signal_802, SubCellOutput[61]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hFC03 ) ) \SubCellInst/GEN[15].SboxInst/y_2 ( .I0 ({Ciphertext_s1[60], Ciphertext_s0[60]}), .I1 ({Ciphertext_s1[61], Ciphertext_s0[61]}), .I2 ({Ciphertext_s1[62], Ciphertext_s0[62]}), .I3 ({Ciphertext_s1[63], Ciphertext_s0[63]}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992]}), .O ({new_AGEMA_signal_803, SubCellOutput[62]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hAAA5 ) ) \SubCellInst/GEN[15].SboxInst/y_3 ( .I0 ({Ciphertext_s1[60], Ciphertext_s0[60]}), .I1 ({Ciphertext_s1[61], Ciphertext_s0[61]}), .I2 ({Ciphertext_s1[62], Ciphertext_s0[62]}), .I3 ({Ciphertext_s1[63], Ciphertext_s0[63]}), .clk (clk), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .O ({new_AGEMA_signal_804, SubCellOutput[63]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<48>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[48], Plaintext_s0[48]}), .I2 ({new_AGEMA_signal_853, \TweakeyGeneration/StateReg/s_current_state [48]}), .I3 ({new_AGEMA_signal_777, SubCellOutput[48]}), .I4 ({new_AGEMA_signal_729, SubCellOutput[24]}), .I5 ({new_AGEMA_signal_705, SubCellOutput[12]}), .O ({new_AGEMA_signal_1002, StateRegInput[48]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<32>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[32], Plaintext_s0[32]}), .I2 ({new_AGEMA_signal_853, \TweakeyGeneration/StateReg/s_current_state [48]}), .I3 ({new_AGEMA_signal_777, SubCellOutput[48]}), .O ({new_AGEMA_signal_1004, StateRegInput[32]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<0>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[0], Plaintext_s0[0]}), .I2 ({new_AGEMA_signal_853, \TweakeyGeneration/StateReg/s_current_state [48]}), .I3 ({new_AGEMA_signal_777, SubCellOutput[48]}), .I4 ({new_AGEMA_signal_729, SubCellOutput[24]}), .O ({new_AGEMA_signal_1006, StateRegInput[0]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<49>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[49], Plaintext_s0[49]}), .I2 ({new_AGEMA_signal_856, \TweakeyGeneration/StateReg/s_current_state [49]}), .I3 ({new_AGEMA_signal_778, SubCellOutput[49]}), .I4 ({new_AGEMA_signal_730, SubCellOutput[25]}), .I5 ({new_AGEMA_signal_706, SubCellOutput[13]}), .O ({new_AGEMA_signal_1008, StateRegInput[49]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<33>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[33], Plaintext_s0[33]}), .I2 ({new_AGEMA_signal_856, \TweakeyGeneration/StateReg/s_current_state [49]}), .I3 ({new_AGEMA_signal_778, SubCellOutput[49]}), .O ({new_AGEMA_signal_1010, StateRegInput[33]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<1>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[1], Plaintext_s0[1]}), .I2 ({new_AGEMA_signal_856, \TweakeyGeneration/StateReg/s_current_state [49]}), .I3 ({new_AGEMA_signal_778, SubCellOutput[49]}), .I4 ({new_AGEMA_signal_730, SubCellOutput[25]}), .O ({new_AGEMA_signal_1012, StateRegInput[1]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<50>1 ( .I0 ({Plaintext_s1[50], Plaintext_s0[50]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_859, \TweakeyGeneration/StateReg/s_current_state [50]}), .I3 ({new_AGEMA_signal_707, SubCellOutput[14]}), .I4 ({new_AGEMA_signal_731, SubCellOutput[26]}), .I5 ({new_AGEMA_signal_779, SubCellOutput[50]}), .O ({new_AGEMA_signal_1014, StateRegInput[50]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \StateRegInput<34>1 ( .I0 ({Plaintext_s1[34], Plaintext_s0[34]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_859, \TweakeyGeneration/StateReg/s_current_state [50]}), .I3 ({new_AGEMA_signal_779, SubCellOutput[50]}), .O ({new_AGEMA_signal_1016, StateRegInput[34]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<2>1 ( .I0 ({Plaintext_s1[2], Plaintext_s0[2]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_859, \TweakeyGeneration/StateReg/s_current_state [50]}), .I3 ({new_AGEMA_signal_731, SubCellOutput[26]}), .I4 ({new_AGEMA_signal_779, SubCellOutput[50]}), .O ({new_AGEMA_signal_1018, StateRegInput[2]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<51>1 ( .I0 ({Plaintext_s1[51], Plaintext_s0[51]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_862, \TweakeyGeneration/StateReg/s_current_state [51]}), .I3 ({new_AGEMA_signal_708, SubCellOutput[15]}), .I4 ({new_AGEMA_signal_732, SubCellOutput[27]}), .I5 ({new_AGEMA_signal_780, SubCellOutput[51]}), .O ({new_AGEMA_signal_1020, StateRegInput[51]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<3>1 ( .I0 ({Plaintext_s1[3], Plaintext_s0[3]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_862, \TweakeyGeneration/StateReg/s_current_state [51]}), .I3 ({new_AGEMA_signal_732, SubCellOutput[27]}), .I4 ({new_AGEMA_signal_780, SubCellOutput[51]}), .O ({new_AGEMA_signal_1022, StateRegInput[3]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \StateRegInput<35>1 ( .I0 ({Plaintext_s1[35], Plaintext_s0[35]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_862, \TweakeyGeneration/StateReg/s_current_state [51]}), .I3 ({new_AGEMA_signal_780, SubCellOutput[51]}), .O ({new_AGEMA_signal_1024, StateRegInput[35]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<52>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[52], Plaintext_s0[52]}), .I2 ({new_AGEMA_signal_865, \TweakeyGeneration/StateReg/s_current_state [52]}), .I3 ({new_AGEMA_signal_785, SubCellOutput[52]}), .I4 ({new_AGEMA_signal_737, SubCellOutput[28]}), .I5 ({new_AGEMA_signal_681, SubCellOutput[0]}), .O ({new_AGEMA_signal_1026, StateRegInput[52]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<4>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[4], Plaintext_s0[4]}), .I2 ({new_AGEMA_signal_865, \TweakeyGeneration/StateReg/s_current_state [52]}), .I3 ({new_AGEMA_signal_785, SubCellOutput[52]}), .I4 ({new_AGEMA_signal_737, SubCellOutput[28]}), .O ({new_AGEMA_signal_1028, StateRegInput[4]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<36>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[36], Plaintext_s0[36]}), .I2 ({new_AGEMA_signal_865, \TweakeyGeneration/StateReg/s_current_state [52]}), .I3 ({new_AGEMA_signal_785, SubCellOutput[52]}), .O ({new_AGEMA_signal_1030, StateRegInput[36]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hD88D8DD88DD8D88D ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<53>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[53], Plaintext_s0[53]}), .I2 ({new_AGEMA_signal_868, \TweakeyGeneration/StateReg/s_current_state [53]}), .I3 ({new_AGEMA_signal_786, SubCellOutput[53]}), .I4 ({new_AGEMA_signal_738, SubCellOutput[29]}), .I5 ({new_AGEMA_signal_682, SubCellOutput[1]}), .O ({new_AGEMA_signal_1032, StateRegInput[53]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h8DD8D88D ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<5>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[5], Plaintext_s0[5]}), .I2 ({new_AGEMA_signal_868, \TweakeyGeneration/StateReg/s_current_state [53]}), .I3 ({new_AGEMA_signal_786, SubCellOutput[53]}), .I4 ({new_AGEMA_signal_738, SubCellOutput[29]}), .O ({new_AGEMA_signal_1034, StateRegInput[5]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<37>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[37], Plaintext_s0[37]}), .I2 ({new_AGEMA_signal_868, \TweakeyGeneration/StateReg/s_current_state [53]}), .I3 ({new_AGEMA_signal_786, SubCellOutput[53]}), .O ({new_AGEMA_signal_1036, StateRegInput[37]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<54>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[54], Plaintext_s0[54]}), .I2 ({new_AGEMA_signal_871, \TweakeyGeneration/StateReg/s_current_state [54]}), .I3 ({new_AGEMA_signal_787, SubCellOutput[54]}), .I4 ({new_AGEMA_signal_739, SubCellOutput[30]}), .I5 ({new_AGEMA_signal_683, SubCellOutput[2]}), .O ({new_AGEMA_signal_1038, StateRegInput[54]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<6>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[6], Plaintext_s0[6]}), .I2 ({new_AGEMA_signal_871, \TweakeyGeneration/StateReg/s_current_state [54]}), .I3 ({new_AGEMA_signal_787, SubCellOutput[54]}), .I4 ({new_AGEMA_signal_739, SubCellOutput[30]}), .O ({new_AGEMA_signal_1040, StateRegInput[6]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<38>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[38], Plaintext_s0[38]}), .I2 ({new_AGEMA_signal_871, \TweakeyGeneration/StateReg/s_current_state [54]}), .I3 ({new_AGEMA_signal_787, SubCellOutput[54]}), .O ({new_AGEMA_signal_1042, StateRegInput[38]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<55>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[55], Plaintext_s0[55]}), .I2 ({new_AGEMA_signal_874, \TweakeyGeneration/StateReg/s_current_state [55]}), .I3 ({new_AGEMA_signal_788, SubCellOutput[55]}), .I4 ({new_AGEMA_signal_740, SubCellOutput[31]}), .I5 ({new_AGEMA_signal_684, SubCellOutput[3]}), .O ({new_AGEMA_signal_1044, StateRegInput[55]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<7>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[7], Plaintext_s0[7]}), .I2 ({new_AGEMA_signal_874, \TweakeyGeneration/StateReg/s_current_state [55]}), .I3 ({new_AGEMA_signal_788, SubCellOutput[55]}), .I4 ({new_AGEMA_signal_740, SubCellOutput[31]}), .O ({new_AGEMA_signal_1046, StateRegInput[7]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<39>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[39], Plaintext_s0[39]}), .I2 ({new_AGEMA_signal_874, \TweakeyGeneration/StateReg/s_current_state [55]}), .I3 ({new_AGEMA_signal_788, SubCellOutput[55]}), .O ({new_AGEMA_signal_1048, StateRegInput[39]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<56>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[56], Plaintext_s0[56]}), .I2 ({new_AGEMA_signal_877, \TweakeyGeneration/StateReg/s_current_state [56]}), .I3 ({new_AGEMA_signal_793, SubCellOutput[56]}), .I4 ({new_AGEMA_signal_713, SubCellOutput[16]}), .I5 ({new_AGEMA_signal_689, SubCellOutput[4]}), .O ({new_AGEMA_signal_1050, StateRegInput[56]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<8>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[8], Plaintext_s0[8]}), .I2 ({new_AGEMA_signal_877, \TweakeyGeneration/StateReg/s_current_state [56]}), .I3 ({new_AGEMA_signal_793, SubCellOutput[56]}), .I4 ({new_AGEMA_signal_713, SubCellOutput[16]}), .O ({new_AGEMA_signal_1052, StateRegInput[8]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<40>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[40], Plaintext_s0[40]}), .I2 ({new_AGEMA_signal_877, \TweakeyGeneration/StateReg/s_current_state [56]}), .I3 ({new_AGEMA_signal_793, SubCellOutput[56]}), .O ({new_AGEMA_signal_1054, StateRegInput[40]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<57>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[57], Plaintext_s0[57]}), .I2 ({new_AGEMA_signal_880, \TweakeyGeneration/StateReg/s_current_state [57]}), .I3 ({new_AGEMA_signal_794, SubCellOutput[57]}), .I4 ({new_AGEMA_signal_714, SubCellOutput[17]}), .I5 ({new_AGEMA_signal_690, SubCellOutput[5]}), .O ({new_AGEMA_signal_1056, StateRegInput[57]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<9>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[9], Plaintext_s0[9]}), .I2 ({new_AGEMA_signal_880, \TweakeyGeneration/StateReg/s_current_state [57]}), .I3 ({new_AGEMA_signal_794, SubCellOutput[57]}), .I4 ({new_AGEMA_signal_714, SubCellOutput[17]}), .O ({new_AGEMA_signal_1058, StateRegInput[9]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<41>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[41], Plaintext_s0[41]}), .I2 ({new_AGEMA_signal_880, \TweakeyGeneration/StateReg/s_current_state [57]}), .I3 ({new_AGEMA_signal_794, SubCellOutput[57]}), .O ({new_AGEMA_signal_1060, StateRegInput[41]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<58>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[58], Plaintext_s0[58]}), .I2 ({new_AGEMA_signal_883, \TweakeyGeneration/StateReg/s_current_state [58]}), .I3 ({new_AGEMA_signal_795, SubCellOutput[58]}), .I4 ({new_AGEMA_signal_715, SubCellOutput[18]}), .I5 ({new_AGEMA_signal_691, SubCellOutput[6]}), .O ({new_AGEMA_signal_1062, StateRegInput[58]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<42>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[42], Plaintext_s0[42]}), .I2 ({new_AGEMA_signal_883, \TweakeyGeneration/StateReg/s_current_state [58]}), .I3 ({new_AGEMA_signal_795, SubCellOutput[58]}), .O ({new_AGEMA_signal_1064, StateRegInput[42]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<10>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[10], Plaintext_s0[10]}), .I2 ({new_AGEMA_signal_883, \TweakeyGeneration/StateReg/s_current_state [58]}), .I3 ({new_AGEMA_signal_795, SubCellOutput[58]}), .I4 ({new_AGEMA_signal_715, SubCellOutput[18]}), .O ({new_AGEMA_signal_1066, StateRegInput[10]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \StateRegInput<59>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[59], Plaintext_s0[59]}), .I2 ({new_AGEMA_signal_886, \TweakeyGeneration/StateReg/s_current_state [59]}), .I3 ({new_AGEMA_signal_796, SubCellOutput[59]}), .I4 ({new_AGEMA_signal_716, SubCellOutput[19]}), .I5 ({new_AGEMA_signal_692, SubCellOutput[7]}), .O ({new_AGEMA_signal_1068, StateRegInput[59]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h8DD8 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'h8DD8 ) ) \StateRegInput<43>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[43], Plaintext_s0[43]}), .I2 ({new_AGEMA_signal_886, \TweakeyGeneration/StateReg/s_current_state [59]}), .I3 ({new_AGEMA_signal_796, SubCellOutput[59]}), .O ({new_AGEMA_signal_1070, StateRegInput[43]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \StateRegInput<11>1 ( .I0 ({1'b0, rst}), .I1 ({Plaintext_s1[11], Plaintext_s0[11]}), .I2 ({new_AGEMA_signal_886, \TweakeyGeneration/StateReg/s_current_state [59]}), .I3 ({new_AGEMA_signal_796, SubCellOutput[59]}), .I4 ({new_AGEMA_signal_716, SubCellOutput[19]}), .O ({new_AGEMA_signal_1072, StateRegInput[11]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b01010 ), .INIT2 ( 32'h8B8BB8B8 ) ) \StateRegInput<44>1 ( .I0 ({Plaintext_s1[44], Plaintext_s0[44]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_889, \TweakeyGeneration/StateReg/s_current_state [60]}), .I3 ({1'b0, \FSMReg/s_current_state [0]}), .I4 ({new_AGEMA_signal_801, SubCellOutput[60]}), .O ({new_AGEMA_signal_1074, StateRegInput[44]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b001010 ), .INIT2 ( 64'hB8B88B8B8B8BB8B8 ) ) \StateRegInput<12>1 ( .I0 ({Plaintext_s1[12], Plaintext_s0[12]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_889, \TweakeyGeneration/StateReg/s_current_state [60]}), .I3 ({1'b0, \FSMReg/s_current_state [0]}), .I4 ({new_AGEMA_signal_801, SubCellOutput[60]}), .I5 ({new_AGEMA_signal_721, SubCellOutput[20]}), .O ({new_AGEMA_signal_1076, StateRegInput[12]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00110 ), .INIT2 ( 32'h88BBBB88 ) ) \StateRegInput<45>1 ( .I0 ({Plaintext_s1[45], Plaintext_s0[45]}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_2_294 }), .I3 ({new_AGEMA_signal_892, \TweakeyGeneration/StateReg/s_current_state [61]}), .I4 ({new_AGEMA_signal_802, SubCellOutput[61]}), .O ({new_AGEMA_signal_1078, StateRegInput[45]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \StateRegInput<13>1 ( .I0 ({Plaintext_s1[13], Plaintext_s0[13]}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_2_294 }), .I3 ({new_AGEMA_signal_892, \TweakeyGeneration/StateReg/s_current_state [61]}), .I4 ({new_AGEMA_signal_802, SubCellOutput[61]}), .I5 ({new_AGEMA_signal_722, SubCellOutput[21]}), .O ({new_AGEMA_signal_1080, StateRegInput[13]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b01010 ), .INIT2 ( 32'h8B8BB8B8 ) ) \StateRegInput<46>1 ( .I0 ({Plaintext_s1[46], Plaintext_s0[46]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_895, \TweakeyGeneration/StateReg/s_current_state [62]}), .I3 ({1'b0, \FSMReg/s_current_state_sliced_3_293 }), .I4 ({new_AGEMA_signal_803, SubCellOutput[62]}), .O ({new_AGEMA_signal_1082, StateRegInput[46]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b001010 ), .INIT2 ( 64'hB8B88B8B8B8BB8B8 ) ) \StateRegInput<14>1 ( .I0 ({Plaintext_s1[14], Plaintext_s0[14]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_895, \TweakeyGeneration/StateReg/s_current_state [62]}), .I3 ({1'b0, \FSMReg/s_current_state_sliced_3_293 }), .I4 ({new_AGEMA_signal_803, SubCellOutput[62]}), .I5 ({new_AGEMA_signal_723, SubCellOutput[22]}), .O ({new_AGEMA_signal_1084, StateRegInput[14]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b01010 ), .INIT2 ( 32'h8B8BB8B8 ) ) \StateRegInput<47>1 ( .I0 ({Plaintext_s1[47], Plaintext_s0[47]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_898, \TweakeyGeneration/StateReg/s_current_state [63]}), .I3 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_1_292 }), .I4 ({new_AGEMA_signal_804, SubCellOutput[63]}), .O ({new_AGEMA_signal_1086, StateRegInput[47]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b001010 ), .INIT2 ( 64'hB8B88B8B8B8BB8B8 ) ) \StateRegInput<15>1 ( .I0 ({Plaintext_s1[15], Plaintext_s0[15]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_898, \TweakeyGeneration/StateReg/s_current_state [63]}), .I3 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_1_292 }), .I4 ({new_AGEMA_signal_804, SubCellOutput[63]}), .I5 ({new_AGEMA_signal_724, SubCellOutput[23]}), .O ({new_AGEMA_signal_1088, StateRegInput[15]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<28>1 ( .I0 ({Plaintext_s1[28], Plaintext_s0[28]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_805, \TweakeyGeneration/StateReg/s_current_state [32]}), .I3 ({new_AGEMA_signal_745, SubCellOutput[32]}), .I4 ({new_AGEMA_signal_721, SubCellOutput[20]}), .O ({new_AGEMA_signal_1090, StateRegInput[28]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<29>1 ( .I0 ({Plaintext_s1[29], Plaintext_s0[29]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_808, \TweakeyGeneration/StateReg/s_current_state [33]}), .I3 ({new_AGEMA_signal_746, SubCellOutput[33]}), .I4 ({new_AGEMA_signal_722, SubCellOutput[21]}), .O ({new_AGEMA_signal_1092, StateRegInput[29]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<30>1 ( .I0 ({Plaintext_s1[30], Plaintext_s0[30]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_811, \TweakeyGeneration/StateReg/s_current_state [34]}), .I3 ({new_AGEMA_signal_747, SubCellOutput[34]}), .I4 ({new_AGEMA_signal_723, SubCellOutput[22]}), .O ({new_AGEMA_signal_1094, StateRegInput[30]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<31>1 ( .I0 ({Plaintext_s1[31], Plaintext_s0[31]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_814, \TweakeyGeneration/StateReg/s_current_state [35]}), .I3 ({new_AGEMA_signal_748, SubCellOutput[35]}), .I4 ({new_AGEMA_signal_724, SubCellOutput[23]}), .O ({new_AGEMA_signal_1096, StateRegInput[31]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<16>1 ( .I0 ({Plaintext_s1[16], Plaintext_s0[16]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_817, \TweakeyGeneration/StateReg/s_current_state [36]}), .I3 ({new_AGEMA_signal_753, SubCellOutput[36]}), .I4 ({new_AGEMA_signal_729, SubCellOutput[24]}), .O ({new_AGEMA_signal_1098, StateRegInput[16]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<17>1 ( .I0 ({Plaintext_s1[17], Plaintext_s0[17]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_820, \TweakeyGeneration/StateReg/s_current_state [37]}), .I3 ({new_AGEMA_signal_754, SubCellOutput[37]}), .I4 ({new_AGEMA_signal_730, SubCellOutput[25]}), .O ({new_AGEMA_signal_1100, StateRegInput[17]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<18>1 ( .I0 ({Plaintext_s1[18], Plaintext_s0[18]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_823, \TweakeyGeneration/StateReg/s_current_state [38]}), .I3 ({new_AGEMA_signal_755, SubCellOutput[38]}), .I4 ({new_AGEMA_signal_731, SubCellOutput[26]}), .O ({new_AGEMA_signal_1102, StateRegInput[18]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<19>1 ( .I0 ({Plaintext_s1[19], Plaintext_s0[19]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_826, \TweakeyGeneration/StateReg/s_current_state [39]}), .I3 ({new_AGEMA_signal_756, SubCellOutput[39]}), .I4 ({new_AGEMA_signal_732, SubCellOutput[27]}), .O ({new_AGEMA_signal_1104, StateRegInput[19]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<20>1 ( .I0 ({Plaintext_s1[20], Plaintext_s0[20]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_829, \TweakeyGeneration/StateReg/s_current_state [40]}), .I3 ({new_AGEMA_signal_761, SubCellOutput[40]}), .I4 ({new_AGEMA_signal_737, SubCellOutput[28]}), .O ({new_AGEMA_signal_1106, StateRegInput[20]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h8BB8B88B ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<21>1 ( .I0 ({Plaintext_s1[21], Plaintext_s0[21]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_832, \TweakeyGeneration/StateReg/s_current_state [41]}), .I3 ({new_AGEMA_signal_762, SubCellOutput[41]}), .I4 ({new_AGEMA_signal_738, SubCellOutput[29]}), .O ({new_AGEMA_signal_1108, StateRegInput[21]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<22>1 ( .I0 ({Plaintext_s1[22], Plaintext_s0[22]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_835, \TweakeyGeneration/StateReg/s_current_state [42]}), .I3 ({new_AGEMA_signal_763, SubCellOutput[42]}), .I4 ({new_AGEMA_signal_739, SubCellOutput[30]}), .O ({new_AGEMA_signal_1110, StateRegInput[22]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<23>1 ( .I0 ({Plaintext_s1[23], Plaintext_s0[23]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_838, \TweakeyGeneration/StateReg/s_current_state [43]}), .I3 ({new_AGEMA_signal_764, SubCellOutput[43]}), .I4 ({new_AGEMA_signal_740, SubCellOutput[31]}), .O ({new_AGEMA_signal_1112, StateRegInput[23]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \StateRegInput<24>1 ( .I0 ({Plaintext_s1[24], Plaintext_s0[24]}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMReg/s_current_state_sliced_sliced_sliced_0_291 }), .I3 ({new_AGEMA_signal_841, \TweakeyGeneration/StateReg/s_current_state [44]}), .I4 ({new_AGEMA_signal_769, SubCellOutput[44]}), .I5 ({new_AGEMA_signal_713, SubCellOutput[16]}), .O ({new_AGEMA_signal_1114, StateRegInput[24]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \StateRegInput<25>1 ( .I0 ({Plaintext_s1[25], Plaintext_s0[25]}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMReg/s_current_state_sliced_sliced_0_290 }), .I3 ({new_AGEMA_signal_844, \TweakeyGeneration/StateReg/s_current_state [45]}), .I4 ({new_AGEMA_signal_770, SubCellOutput[45]}), .I5 ({new_AGEMA_signal_714, SubCellOutput[17]}), .O ({new_AGEMA_signal_1116, StateRegInput[25]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<26>1 ( .I0 ({Plaintext_s1[26], Plaintext_s0[26]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_847, \TweakeyGeneration/StateReg/s_current_state [46]}), .I3 ({new_AGEMA_signal_771, SubCellOutput[46]}), .I4 ({new_AGEMA_signal_715, SubCellOutput[18]}), .O ({new_AGEMA_signal_1118, StateRegInput[26]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \StateRegInput<27>1 ( .I0 ({Plaintext_s1[27], Plaintext_s0[27]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_850, \TweakeyGeneration/StateReg/s_current_state [47]}), .I3 ({new_AGEMA_signal_772, SubCellOutput[47]}), .I4 ({new_AGEMA_signal_716, SubCellOutput[19]}), .O ({new_AGEMA_signal_1120, StateRegInput[27]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<60> ( .I0 ({Plaintext_s1[60], Plaintext_s0[60]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_997, N01}), .I3 ({new_AGEMA_signal_697, SubCellOutput[8]}), .I4 ({new_AGEMA_signal_721, SubCellOutput[20]}), .I5 ({new_AGEMA_signal_801, SubCellOutput[60]}), .O ({new_AGEMA_signal_1122, StateRegInput[60]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<61> ( .I0 ({Plaintext_s1[61], Plaintext_s0[61]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_998, N2}), .I3 ({new_AGEMA_signal_698, SubCellOutput[9]}), .I4 ({new_AGEMA_signal_722, SubCellOutput[21]}), .I5 ({new_AGEMA_signal_802, SubCellOutput[61]}), .O ({new_AGEMA_signal_1124, StateRegInput[61]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<62> ( .I0 ({Plaintext_s1[62], Plaintext_s0[62]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_999, N4}), .I3 ({new_AGEMA_signal_699, SubCellOutput[10]}), .I4 ({new_AGEMA_signal_723, SubCellOutput[22]}), .I5 ({new_AGEMA_signal_803, SubCellOutput[62]}), .O ({new_AGEMA_signal_1126, StateRegInput[62]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h8BB8B88BB88B8BB8 ) ) \StateRegInput<63> ( .I0 ({Plaintext_s1[63], Plaintext_s0[63]}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_1000, N6}), .I3 ({new_AGEMA_signal_700, SubCellOutput[11]}), .I4 ({new_AGEMA_signal_724, SubCellOutput[23]}), .I5 ({new_AGEMA_signal_804, SubCellOutput[63]}), .O ({new_AGEMA_signal_1128, StateRegInput[63]}) ) ;

    /* register cells */
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_63 ( .D ({new_AGEMA_signal_996, \TweakeyGeneration/StateRegInput [63]}), .clk (clk_gated), .Q ({new_AGEMA_signal_898, \TweakeyGeneration/StateReg/s_current_state [63]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_62 ( .D ({new_AGEMA_signal_993, \TweakeyGeneration/StateRegInput [62]}), .clk (clk_gated), .Q ({new_AGEMA_signal_895, \TweakeyGeneration/StateReg/s_current_state [62]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_61 ( .D ({new_AGEMA_signal_990, \TweakeyGeneration/StateRegInput [61]}), .clk (clk_gated), .Q ({new_AGEMA_signal_892, \TweakeyGeneration/StateReg/s_current_state [61]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_60 ( .D ({new_AGEMA_signal_987, \TweakeyGeneration/StateRegInput [60]}), .clk (clk_gated), .Q ({new_AGEMA_signal_889, \TweakeyGeneration/StateReg/s_current_state [60]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_59 ( .D ({new_AGEMA_signal_984, \TweakeyGeneration/StateRegInput [59]}), .clk (clk_gated), .Q ({new_AGEMA_signal_886, \TweakeyGeneration/StateReg/s_current_state [59]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_58 ( .D ({new_AGEMA_signal_981, \TweakeyGeneration/StateRegInput [58]}), .clk (clk_gated), .Q ({new_AGEMA_signal_883, \TweakeyGeneration/StateReg/s_current_state [58]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_57 ( .D ({new_AGEMA_signal_978, \TweakeyGeneration/StateRegInput [57]}), .clk (clk_gated), .Q ({new_AGEMA_signal_880, \TweakeyGeneration/StateReg/s_current_state [57]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_56 ( .D ({new_AGEMA_signal_975, \TweakeyGeneration/StateRegInput [56]}), .clk (clk_gated), .Q ({new_AGEMA_signal_877, \TweakeyGeneration/StateReg/s_current_state [56]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_55 ( .D ({new_AGEMA_signal_972, \TweakeyGeneration/StateRegInput [55]}), .clk (clk_gated), .Q ({new_AGEMA_signal_874, \TweakeyGeneration/StateReg/s_current_state [55]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_54 ( .D ({new_AGEMA_signal_969, \TweakeyGeneration/StateRegInput [54]}), .clk (clk_gated), .Q ({new_AGEMA_signal_871, \TweakeyGeneration/StateReg/s_current_state [54]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_53 ( .D ({new_AGEMA_signal_966, \TweakeyGeneration/StateRegInput [53]}), .clk (clk_gated), .Q ({new_AGEMA_signal_868, \TweakeyGeneration/StateReg/s_current_state [53]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_52 ( .D ({new_AGEMA_signal_963, \TweakeyGeneration/StateRegInput [52]}), .clk (clk_gated), .Q ({new_AGEMA_signal_865, \TweakeyGeneration/StateReg/s_current_state [52]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_51 ( .D ({new_AGEMA_signal_960, \TweakeyGeneration/StateRegInput [51]}), .clk (clk_gated), .Q ({new_AGEMA_signal_862, \TweakeyGeneration/StateReg/s_current_state [51]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_50 ( .D ({new_AGEMA_signal_957, \TweakeyGeneration/StateRegInput [50]}), .clk (clk_gated), .Q ({new_AGEMA_signal_859, \TweakeyGeneration/StateReg/s_current_state [50]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_49 ( .D ({new_AGEMA_signal_954, \TweakeyGeneration/StateRegInput [49]}), .clk (clk_gated), .Q ({new_AGEMA_signal_856, \TweakeyGeneration/StateReg/s_current_state [49]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_48 ( .D ({new_AGEMA_signal_951, \TweakeyGeneration/StateRegInput [48]}), .clk (clk_gated), .Q ({new_AGEMA_signal_853, \TweakeyGeneration/StateReg/s_current_state [48]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_47 ( .D ({new_AGEMA_signal_948, \TweakeyGeneration/StateRegInput [47]}), .clk (clk_gated), .Q ({new_AGEMA_signal_850, \TweakeyGeneration/StateReg/s_current_state [47]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_46 ( .D ({new_AGEMA_signal_945, \TweakeyGeneration/StateRegInput [46]}), .clk (clk_gated), .Q ({new_AGEMA_signal_847, \TweakeyGeneration/StateReg/s_current_state [46]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_45 ( .D ({new_AGEMA_signal_942, \TweakeyGeneration/StateRegInput [45]}), .clk (clk_gated), .Q ({new_AGEMA_signal_844, \TweakeyGeneration/StateReg/s_current_state [45]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_44 ( .D ({new_AGEMA_signal_939, \TweakeyGeneration/StateRegInput [44]}), .clk (clk_gated), .Q ({new_AGEMA_signal_841, \TweakeyGeneration/StateReg/s_current_state [44]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_43 ( .D ({new_AGEMA_signal_936, \TweakeyGeneration/StateRegInput [43]}), .clk (clk_gated), .Q ({new_AGEMA_signal_838, \TweakeyGeneration/StateReg/s_current_state [43]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_42 ( .D ({new_AGEMA_signal_933, \TweakeyGeneration/StateRegInput [42]}), .clk (clk_gated), .Q ({new_AGEMA_signal_835, \TweakeyGeneration/StateReg/s_current_state [42]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_41 ( .D ({new_AGEMA_signal_930, \TweakeyGeneration/StateRegInput [41]}), .clk (clk_gated), .Q ({new_AGEMA_signal_832, \TweakeyGeneration/StateReg/s_current_state [41]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_40 ( .D ({new_AGEMA_signal_927, \TweakeyGeneration/StateRegInput [40]}), .clk (clk_gated), .Q ({new_AGEMA_signal_829, \TweakeyGeneration/StateReg/s_current_state [40]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_39 ( .D ({new_AGEMA_signal_924, \TweakeyGeneration/StateRegInput [39]}), .clk (clk_gated), .Q ({new_AGEMA_signal_826, \TweakeyGeneration/StateReg/s_current_state [39]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_38 ( .D ({new_AGEMA_signal_921, \TweakeyGeneration/StateRegInput [38]}), .clk (clk_gated), .Q ({new_AGEMA_signal_823, \TweakeyGeneration/StateReg/s_current_state [38]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_37 ( .D ({new_AGEMA_signal_918, \TweakeyGeneration/StateRegInput [37]}), .clk (clk_gated), .Q ({new_AGEMA_signal_820, \TweakeyGeneration/StateReg/s_current_state [37]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_36 ( .D ({new_AGEMA_signal_915, \TweakeyGeneration/StateRegInput [36]}), .clk (clk_gated), .Q ({new_AGEMA_signal_817, \TweakeyGeneration/StateReg/s_current_state [36]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_35 ( .D ({new_AGEMA_signal_912, \TweakeyGeneration/StateRegInput [35]}), .clk (clk_gated), .Q ({new_AGEMA_signal_814, \TweakeyGeneration/StateReg/s_current_state [35]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_34 ( .D ({new_AGEMA_signal_909, \TweakeyGeneration/StateRegInput [34]}), .clk (clk_gated), .Q ({new_AGEMA_signal_811, \TweakeyGeneration/StateReg/s_current_state [34]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_33 ( .D ({new_AGEMA_signal_906, \TweakeyGeneration/StateRegInput [33]}), .clk (clk_gated), .Q ({new_AGEMA_signal_808, \TweakeyGeneration/StateReg/s_current_state [33]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_32 ( .D ({new_AGEMA_signal_903, \TweakeyGeneration/StateRegInput [32]}), .clk (clk_gated), .Q ({new_AGEMA_signal_805, \TweakeyGeneration/StateReg/s_current_state [32]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_31 ( .D ({new_AGEMA_signal_900, \TweakeyGeneration/StateRegInput [31]}), .clk (clk_gated), .Q ({new_AGEMA_signal_970, \TweakeyGeneration/StateReg/s_current_state [31]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_30 ( .D ({new_AGEMA_signal_897, \TweakeyGeneration/StateRegInput [30]}), .clk (clk_gated), .Q ({new_AGEMA_signal_967, \TweakeyGeneration/StateReg/s_current_state [30]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_29 ( .D ({new_AGEMA_signal_894, \TweakeyGeneration/StateRegInput [29]}), .clk (clk_gated), .Q ({new_AGEMA_signal_964, \TweakeyGeneration/StateReg/s_current_state [29]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_28 ( .D ({new_AGEMA_signal_891, \TweakeyGeneration/StateRegInput [28]}), .clk (clk_gated), .Q ({new_AGEMA_signal_961, \TweakeyGeneration/StateReg/s_current_state [28]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_27 ( .D ({new_AGEMA_signal_888, \TweakeyGeneration/StateRegInput [27]}), .clk (clk_gated), .Q ({new_AGEMA_signal_994, \TweakeyGeneration/StateReg/s_current_state [27]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_26 ( .D ({new_AGEMA_signal_885, \TweakeyGeneration/StateRegInput [26]}), .clk (clk_gated), .Q ({new_AGEMA_signal_991, \TweakeyGeneration/StateReg/s_current_state [26]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_25 ( .D ({new_AGEMA_signal_882, \TweakeyGeneration/StateRegInput [25]}), .clk (clk_gated), .Q ({new_AGEMA_signal_988, \TweakeyGeneration/StateReg/s_current_state [25]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_24 ( .D ({new_AGEMA_signal_879, \TweakeyGeneration/StateRegInput [24]}), .clk (clk_gated), .Q ({new_AGEMA_signal_985, \TweakeyGeneration/StateReg/s_current_state [24]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_23 ( .D ({new_AGEMA_signal_876, \TweakeyGeneration/StateRegInput [23]}), .clk (clk_gated), .Q ({new_AGEMA_signal_946, \TweakeyGeneration/StateReg/s_current_state [23]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_22 ( .D ({new_AGEMA_signal_873, \TweakeyGeneration/StateRegInput [22]}), .clk (clk_gated), .Q ({new_AGEMA_signal_943, \TweakeyGeneration/StateReg/s_current_state [22]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_21 ( .D ({new_AGEMA_signal_870, \TweakeyGeneration/StateRegInput [21]}), .clk (clk_gated), .Q ({new_AGEMA_signal_940, \TweakeyGeneration/StateReg/s_current_state [21]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_20 ( .D ({new_AGEMA_signal_867, \TweakeyGeneration/StateRegInput [20]}), .clk (clk_gated), .Q ({new_AGEMA_signal_937, \TweakeyGeneration/StateReg/s_current_state [20]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_19 ( .D ({new_AGEMA_signal_864, \TweakeyGeneration/StateRegInput [19]}), .clk (clk_gated), .Q ({new_AGEMA_signal_910, \TweakeyGeneration/StateReg/s_current_state [19]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_18 ( .D ({new_AGEMA_signal_861, \TweakeyGeneration/StateRegInput [18]}), .clk (clk_gated), .Q ({new_AGEMA_signal_907, \TweakeyGeneration/StateReg/s_current_state [18]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_17 ( .D ({new_AGEMA_signal_858, \TweakeyGeneration/StateRegInput [17]}), .clk (clk_gated), .Q ({new_AGEMA_signal_904, \TweakeyGeneration/StateReg/s_current_state [17]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_16 ( .D ({new_AGEMA_signal_855, \TweakeyGeneration/StateRegInput [16]}), .clk (clk_gated), .Q ({new_AGEMA_signal_901, \TweakeyGeneration/StateReg/s_current_state [16]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_15 ( .D ({new_AGEMA_signal_852, \TweakeyGeneration/StateRegInput [15]}), .clk (clk_gated), .Q ({new_AGEMA_signal_922, \TweakeyGeneration/StateReg/s_current_state [15]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_14 ( .D ({new_AGEMA_signal_849, \TweakeyGeneration/StateRegInput [14]}), .clk (clk_gated), .Q ({new_AGEMA_signal_919, \TweakeyGeneration/StateReg/s_current_state [14]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_13 ( .D ({new_AGEMA_signal_846, \TweakeyGeneration/StateRegInput [13]}), .clk (clk_gated), .Q ({new_AGEMA_signal_916, \TweakeyGeneration/StateReg/s_current_state [13]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_12 ( .D ({new_AGEMA_signal_843, \TweakeyGeneration/StateRegInput [12]}), .clk (clk_gated), .Q ({new_AGEMA_signal_913, \TweakeyGeneration/StateReg/s_current_state [12]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_11 ( .D ({new_AGEMA_signal_840, \TweakeyGeneration/StateRegInput [11]}), .clk (clk_gated), .Q ({new_AGEMA_signal_958, \TweakeyGeneration/StateReg/s_current_state [11]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_10 ( .D ({new_AGEMA_signal_837, \TweakeyGeneration/StateRegInput [10]}), .clk (clk_gated), .Q ({new_AGEMA_signal_955, \TweakeyGeneration/StateReg/s_current_state [10]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_9 ( .D ({new_AGEMA_signal_834, \TweakeyGeneration/StateRegInput [9]}), .clk (clk_gated), .Q ({new_AGEMA_signal_952, \TweakeyGeneration/StateReg/s_current_state [9]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_8 ( .D ({new_AGEMA_signal_831, \TweakeyGeneration/StateRegInput [8]}), .clk (clk_gated), .Q ({new_AGEMA_signal_949, \TweakeyGeneration/StateReg/s_current_state [8]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_7 ( .D ({new_AGEMA_signal_828, \TweakeyGeneration/StateRegInput [7]}), .clk (clk_gated), .Q ({new_AGEMA_signal_934, \TweakeyGeneration/StateReg/s_current_state [7]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_6 ( .D ({new_AGEMA_signal_825, \TweakeyGeneration/StateRegInput [6]}), .clk (clk_gated), .Q ({new_AGEMA_signal_931, \TweakeyGeneration/StateReg/s_current_state [6]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_5 ( .D ({new_AGEMA_signal_822, \TweakeyGeneration/StateRegInput [5]}), .clk (clk_gated), .Q ({new_AGEMA_signal_928, \TweakeyGeneration/StateReg/s_current_state [5]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_4 ( .D ({new_AGEMA_signal_819, \TweakeyGeneration/StateRegInput [4]}), .clk (clk_gated), .Q ({new_AGEMA_signal_925, \TweakeyGeneration/StateReg/s_current_state [4]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_3 ( .D ({new_AGEMA_signal_816, \TweakeyGeneration/StateRegInput [3]}), .clk (clk_gated), .Q ({new_AGEMA_signal_982, \TweakeyGeneration/StateReg/s_current_state [3]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_2 ( .D ({new_AGEMA_signal_813, \TweakeyGeneration/StateRegInput [2]}), .clk (clk_gated), .Q ({new_AGEMA_signal_979, \TweakeyGeneration/StateReg/s_current_state [2]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_1 ( .D ({new_AGEMA_signal_810, \TweakeyGeneration/StateRegInput [1]}), .clk (clk_gated), .Q ({new_AGEMA_signal_976, \TweakeyGeneration/StateReg/s_current_state [1]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \TweakeyGeneration/StateReg/s_current_state_0 ( .D ({new_AGEMA_signal_807, \TweakeyGeneration/StateRegInput [0]}), .clk (clk_gated), .Q ({new_AGEMA_signal_973, \TweakeyGeneration/StateReg/s_current_state [0]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_63 ( .D ({new_AGEMA_signal_1128, StateRegInput[63]}), .clk (clk_gated), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_62 ( .D ({new_AGEMA_signal_1126, StateRegInput[62]}), .clk (clk_gated), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_61 ( .D ({new_AGEMA_signal_1124, StateRegInput[61]}), .clk (clk_gated), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_60 ( .D ({new_AGEMA_signal_1122, StateRegInput[60]}), .clk (clk_gated), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_59 ( .D ({new_AGEMA_signal_1068, StateRegInput[59]}), .clk (clk_gated), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_58 ( .D ({new_AGEMA_signal_1062, StateRegInput[58]}), .clk (clk_gated), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_57 ( .D ({new_AGEMA_signal_1056, StateRegInput[57]}), .clk (clk_gated), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_56 ( .D ({new_AGEMA_signal_1050, StateRegInput[56]}), .clk (clk_gated), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_55 ( .D ({new_AGEMA_signal_1044, StateRegInput[55]}), .clk (clk_gated), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_54 ( .D ({new_AGEMA_signal_1038, StateRegInput[54]}), .clk (clk_gated), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_53 ( .D ({new_AGEMA_signal_1032, StateRegInput[53]}), .clk (clk_gated), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_52 ( .D ({new_AGEMA_signal_1026, StateRegInput[52]}), .clk (clk_gated), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_51 ( .D ({new_AGEMA_signal_1020, StateRegInput[51]}), .clk (clk_gated), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_50 ( .D ({new_AGEMA_signal_1014, StateRegInput[50]}), .clk (clk_gated), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_49 ( .D ({new_AGEMA_signal_1008, StateRegInput[49]}), .clk (clk_gated), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_48 ( .D ({new_AGEMA_signal_1002, StateRegInput[48]}), .clk (clk_gated), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_47 ( .D ({new_AGEMA_signal_1086, StateRegInput[47]}), .clk (clk_gated), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_46 ( .D ({new_AGEMA_signal_1082, StateRegInput[46]}), .clk (clk_gated), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_45 ( .D ({new_AGEMA_signal_1078, StateRegInput[45]}), .clk (clk_gated), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_44 ( .D ({new_AGEMA_signal_1074, StateRegInput[44]}), .clk (clk_gated), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_43 ( .D ({new_AGEMA_signal_1070, StateRegInput[43]}), .clk (clk_gated), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_42 ( .D ({new_AGEMA_signal_1064, StateRegInput[42]}), .clk (clk_gated), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_41 ( .D ({new_AGEMA_signal_1060, StateRegInput[41]}), .clk (clk_gated), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_40 ( .D ({new_AGEMA_signal_1054, StateRegInput[40]}), .clk (clk_gated), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_39 ( .D ({new_AGEMA_signal_1048, StateRegInput[39]}), .clk (clk_gated), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_38 ( .D ({new_AGEMA_signal_1042, StateRegInput[38]}), .clk (clk_gated), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_37 ( .D ({new_AGEMA_signal_1036, StateRegInput[37]}), .clk (clk_gated), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_36 ( .D ({new_AGEMA_signal_1030, StateRegInput[36]}), .clk (clk_gated), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_35 ( .D ({new_AGEMA_signal_1024, StateRegInput[35]}), .clk (clk_gated), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_34 ( .D ({new_AGEMA_signal_1016, StateRegInput[34]}), .clk (clk_gated), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_33 ( .D ({new_AGEMA_signal_1010, StateRegInput[33]}), .clk (clk_gated), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_32 ( .D ({new_AGEMA_signal_1004, StateRegInput[32]}), .clk (clk_gated), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_31 ( .D ({new_AGEMA_signal_1096, StateRegInput[31]}), .clk (clk_gated), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_30 ( .D ({new_AGEMA_signal_1094, StateRegInput[30]}), .clk (clk_gated), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_29 ( .D ({new_AGEMA_signal_1092, StateRegInput[29]}), .clk (clk_gated), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_28 ( .D ({new_AGEMA_signal_1090, StateRegInput[28]}), .clk (clk_gated), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_27 ( .D ({new_AGEMA_signal_1120, StateRegInput[27]}), .clk (clk_gated), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_26 ( .D ({new_AGEMA_signal_1118, StateRegInput[26]}), .clk (clk_gated), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_25 ( .D ({new_AGEMA_signal_1116, StateRegInput[25]}), .clk (clk_gated), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_24 ( .D ({new_AGEMA_signal_1114, StateRegInput[24]}), .clk (clk_gated), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_23 ( .D ({new_AGEMA_signal_1112, StateRegInput[23]}), .clk (clk_gated), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_22 ( .D ({new_AGEMA_signal_1110, StateRegInput[22]}), .clk (clk_gated), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_21 ( .D ({new_AGEMA_signal_1108, StateRegInput[21]}), .clk (clk_gated), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_20 ( .D ({new_AGEMA_signal_1106, StateRegInput[20]}), .clk (clk_gated), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_19 ( .D ({new_AGEMA_signal_1104, StateRegInput[19]}), .clk (clk_gated), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_18 ( .D ({new_AGEMA_signal_1102, StateRegInput[18]}), .clk (clk_gated), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_17 ( .D ({new_AGEMA_signal_1100, StateRegInput[17]}), .clk (clk_gated), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_16 ( .D ({new_AGEMA_signal_1098, StateRegInput[16]}), .clk (clk_gated), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_15 ( .D ({new_AGEMA_signal_1088, StateRegInput[15]}), .clk (clk_gated), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_14 ( .D ({new_AGEMA_signal_1084, StateRegInput[14]}), .clk (clk_gated), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_13 ( .D ({new_AGEMA_signal_1080, StateRegInput[13]}), .clk (clk_gated), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_12 ( .D ({new_AGEMA_signal_1076, StateRegInput[12]}), .clk (clk_gated), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_11 ( .D ({new_AGEMA_signal_1072, StateRegInput[11]}), .clk (clk_gated), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_10 ( .D ({new_AGEMA_signal_1066, StateRegInput[10]}), .clk (clk_gated), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_9 ( .D ({new_AGEMA_signal_1058, StateRegInput[9]}), .clk (clk_gated), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_8 ( .D ({new_AGEMA_signal_1052, StateRegInput[8]}), .clk (clk_gated), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_7 ( .D ({new_AGEMA_signal_1046, StateRegInput[7]}), .clk (clk_gated), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_6 ( .D ({new_AGEMA_signal_1040, StateRegInput[6]}), .clk (clk_gated), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_5 ( .D ({new_AGEMA_signal_1034, StateRegInput[5]}), .clk (clk_gated), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_4 ( .D ({new_AGEMA_signal_1028, StateRegInput[4]}), .clk (clk_gated), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_3 ( .D ({new_AGEMA_signal_1022, StateRegInput[3]}), .clk (clk_gated), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_2 ( .D ({new_AGEMA_signal_1018, StateRegInput[2]}), .clk (clk_gated), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_1 ( .D ({new_AGEMA_signal_1012, StateRegInput[1]}), .clk (clk_gated), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_0 ( .D ({new_AGEMA_signal_1006, StateRegInput[0]}), .clk (clk_gated), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_sliced_sliced_sliced_0 ( .D (FSMSelected[4]), .C (clk_gated), .Q (\FSMReg/s_current_state_sliced_sliced_sliced_0_291 ) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_sliced_sliced_sliced_1 ( .D (FSMSelected[3]), .C (clk_gated), .Q (\FSMReg/s_current_state_sliced_sliced_sliced_1_292 ) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_sliced_sliced_sliced_2 ( .D (FSMSelected[1]), .C (clk_gated), .Q (\FSMReg/s_current_state_sliced_sliced_sliced_2_294 ) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_sliced_sliced_0 ( .D (FSMSelected[5]), .C (clk_gated), .Q (\FSMReg/s_current_state_sliced_sliced_0_290 ) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_sliced_3 ( .D (FSMSelected[2]), .C (clk_gated), .Q (\FSMReg/s_current_state_sliced_3_293 ) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMReg/s_current_state_0 ( .D (FSMSelected[0]), .C (clk_gated), .Q (\FSMReg/s_current_state [0]) ) ;
endmodule
