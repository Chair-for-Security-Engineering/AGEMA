////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module SkinnyTop in file /AGEMA/Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module SkinnyTop_HPC3_Pipeline_d2 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Key_s2, Plaintext_s1, Plaintext_s2, Fresh, Ciphertext_s0, done, Ciphertext_s1, Ciphertext_s2);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Key_s2 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Plaintext_s2 ;
    input [383:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output [63:0] Ciphertext_s2 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_YY_0_ ;
    wire SubCellInst_SboxInst_0_YY_1_ ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_0_XX_1_ ;
    wire SubCellInst_SboxInst_0_XX_2_ ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_YY_0_ ;
    wire SubCellInst_SboxInst_1_YY_1_ ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_1_XX_1_ ;
    wire SubCellInst_SboxInst_1_XX_2_ ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_YY_0_ ;
    wire SubCellInst_SboxInst_2_YY_1_ ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_2_XX_1_ ;
    wire SubCellInst_SboxInst_2_XX_2_ ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_YY_0_ ;
    wire SubCellInst_SboxInst_3_YY_1_ ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_3_XX_1_ ;
    wire SubCellInst_SboxInst_3_XX_2_ ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_YY_0_ ;
    wire SubCellInst_SboxInst_4_YY_1_ ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_4_XX_1_ ;
    wire SubCellInst_SboxInst_4_XX_2_ ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_YY_0_ ;
    wire SubCellInst_SboxInst_5_YY_1_ ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_5_XX_1_ ;
    wire SubCellInst_SboxInst_5_XX_2_ ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_YY_0_ ;
    wire SubCellInst_SboxInst_6_YY_1_ ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_6_XX_1_ ;
    wire SubCellInst_SboxInst_6_XX_2_ ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_YY_0_ ;
    wire SubCellInst_SboxInst_7_YY_1_ ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_7_XX_1_ ;
    wire SubCellInst_SboxInst_7_XX_2_ ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_YY_0_ ;
    wire SubCellInst_SboxInst_8_YY_1_ ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_8_XX_1_ ;
    wire SubCellInst_SboxInst_8_XX_2_ ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_YY_0_ ;
    wire SubCellInst_SboxInst_9_YY_1_ ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_9_XX_1_ ;
    wire SubCellInst_SboxInst_9_XX_2_ ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_YY_0_ ;
    wire SubCellInst_SboxInst_10_YY_1_ ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_10_XX_1_ ;
    wire SubCellInst_SboxInst_10_XX_2_ ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_YY_0_ ;
    wire SubCellInst_SboxInst_11_YY_1_ ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_11_XX_1_ ;
    wire SubCellInst_SboxInst_11_XX_2_ ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_YY_0_ ;
    wire SubCellInst_SboxInst_12_YY_1_ ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_12_XX_1_ ;
    wire SubCellInst_SboxInst_12_XX_2_ ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_YY_0_ ;
    wire SubCellInst_SboxInst_13_YY_1_ ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_13_XX_1_ ;
    wire SubCellInst_SboxInst_13_XX_2_ ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_YY_0_ ;
    wire SubCellInst_SboxInst_14_YY_1_ ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_14_XX_1_ ;
    wire SubCellInst_SboxInst_14_XX_2_ ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_YY_0_ ;
    wire SubCellInst_SboxInst_15_YY_1_ ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire SubCellInst_SboxInst_15_XX_1_ ;
    wire SubCellInst_SboxInst_15_XX_2_ ;
    wire AddConstXOR_AddConstXOR_XORInst_0_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_3_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_3_n1 ;
    wire MCInst_MCR0_XORInst_0_0_n2 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n2 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n2 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n2 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n2 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n2 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n2 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n2 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n2 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n2 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n2 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n2 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n2 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n2 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n2 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n2 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire MCInst_MCR2_XORInst_0_0_n1 ;
    wire MCInst_MCR2_XORInst_0_1_n1 ;
    wire MCInst_MCR2_XORInst_0_2_n1 ;
    wire MCInst_MCR2_XORInst_0_3_n1 ;
    wire MCInst_MCR2_XORInst_1_0_n1 ;
    wire MCInst_MCR2_XORInst_1_1_n1 ;
    wire MCInst_MCR2_XORInst_1_2_n1 ;
    wire MCInst_MCR2_XORInst_1_3_n1 ;
    wire MCInst_MCR2_XORInst_2_0_n1 ;
    wire MCInst_MCR2_XORInst_2_1_n1 ;
    wire MCInst_MCR2_XORInst_2_2_n1 ;
    wire MCInst_MCR2_XORInst_2_3_n1 ;
    wire MCInst_MCR2_XORInst_3_0_n1 ;
    wire MCInst_MCR2_XORInst_3_1_n1 ;
    wire MCInst_MCR2_XORInst_3_2_n1 ;
    wire MCInst_MCR2_XORInst_3_3_n1 ;
    wire MCInst_MCR3_XORInst_0_0_n1 ;
    wire MCInst_MCR3_XORInst_0_1_n1 ;
    wire MCInst_MCR3_XORInst_0_2_n1 ;
    wire MCInst_MCR3_XORInst_0_3_n1 ;
    wire MCInst_MCR3_XORInst_1_0_n1 ;
    wire MCInst_MCR3_XORInst_1_1_n1 ;
    wire MCInst_MCR3_XORInst_1_2_n1 ;
    wire MCInst_MCR3_XORInst_1_3_n1 ;
    wire MCInst_MCR3_XORInst_2_0_n1 ;
    wire MCInst_MCR3_XORInst_2_1_n1 ;
    wire MCInst_MCR3_XORInst_2_2_n1 ;
    wire MCInst_MCR3_XORInst_2_3_n1 ;
    wire MCInst_MCR3_XORInst_3_0_n1 ;
    wire MCInst_MCR3_XORInst_3_1_n1 ;
    wire MCInst_MCR3_XORInst_3_2_n1 ;
    wire MCInst_MCR3_XORInst_3_3_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire FSMSignalsInst_doneInst_n1 ;
    wire [63:0] MCOutput ;
    wire [63:0] StateRegInput ;
    wire [63:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [5:0] FSMSelected ;
    wire [63:0] TweakeyGeneration_StateRegInput ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U1 ( .a ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .a ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .a ({Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR0_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, SubCellInst_SboxInst_0_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR1_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR3_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR5_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, SubCellInst_SboxInst_0_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR6_U1 ( .a ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}), .b ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, SubCellInst_SboxInst_0_Q6}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, SubCellInst_SboxInst_0_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR8_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, SubCellInst_SboxInst_0_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U1 ( .a ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .a ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, SubCellInst_SboxInst_1_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .a ({Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR0_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, SubCellInst_SboxInst_1_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR1_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, SubCellInst_SboxInst_1_XX_1_}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR3_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, SubCellInst_SboxInst_1_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR5_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR6_U1 ( .a ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, SubCellInst_SboxInst_1_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR8_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, SubCellInst_SboxInst_1_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U1 ( .a ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .a ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .a ({Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR0_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, SubCellInst_SboxInst_2_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR1_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR3_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR5_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, SubCellInst_SboxInst_2_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR6_U1 ( .a ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}), .b ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, SubCellInst_SboxInst_2_Q6}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, SubCellInst_SboxInst_2_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR8_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, SubCellInst_SboxInst_2_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U1 ( .a ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .a ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, SubCellInst_SboxInst_3_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .a ({Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR0_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, SubCellInst_SboxInst_3_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR1_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, SubCellInst_SboxInst_3_XX_1_}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR3_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, SubCellInst_SboxInst_3_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR5_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR6_U1 ( .a ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, SubCellInst_SboxInst_3_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR8_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, SubCellInst_SboxInst_3_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U1 ( .a ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .a ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .a ({Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR0_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, SubCellInst_SboxInst_4_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR1_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR3_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR5_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, SubCellInst_SboxInst_4_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR6_U1 ( .a ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}), .b ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, SubCellInst_SboxInst_4_Q6}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, SubCellInst_SboxInst_4_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR8_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, SubCellInst_SboxInst_4_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U1 ( .a ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .a ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, SubCellInst_SboxInst_5_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .a ({Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR0_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, SubCellInst_SboxInst_5_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR1_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, SubCellInst_SboxInst_5_XX_1_}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR3_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, SubCellInst_SboxInst_5_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR5_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR6_U1 ( .a ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, SubCellInst_SboxInst_5_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR8_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, SubCellInst_SboxInst_5_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U1 ( .a ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .a ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .a ({Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR0_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, SubCellInst_SboxInst_6_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR1_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR3_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR5_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, SubCellInst_SboxInst_6_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR6_U1 ( .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}), .b ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, SubCellInst_SboxInst_6_Q6}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, SubCellInst_SboxInst_6_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR8_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, SubCellInst_SboxInst_6_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U1 ( .a ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .a ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, SubCellInst_SboxInst_7_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .a ({Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR0_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, SubCellInst_SboxInst_7_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR1_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, SubCellInst_SboxInst_7_XX_1_}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR3_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, SubCellInst_SboxInst_7_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR5_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR6_U1 ( .a ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, SubCellInst_SboxInst_7_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR8_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, SubCellInst_SboxInst_7_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U1 ( .a ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .a ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .a ({Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR0_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, SubCellInst_SboxInst_8_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR1_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR3_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR5_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_8_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR6_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}), .b ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_8_Q6}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, SubCellInst_SboxInst_8_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR8_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, SubCellInst_SboxInst_8_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U1 ( .a ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .a ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, SubCellInst_SboxInst_9_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .a ({Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR0_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, SubCellInst_SboxInst_9_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR1_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, SubCellInst_SboxInst_9_XX_1_}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR3_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, SubCellInst_SboxInst_9_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR5_U1 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR6_U1 ( .a ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}), .b ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, SubCellInst_SboxInst_9_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR8_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, SubCellInst_SboxInst_9_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U1 ( .a ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .a ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .a ({Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR0_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, SubCellInst_SboxInst_10_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR1_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR3_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR5_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_10_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR6_U1 ( .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_10_Q6}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, SubCellInst_SboxInst_10_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR8_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, SubCellInst_SboxInst_10_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U1 ( .a ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .a ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, SubCellInst_SboxInst_11_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .a ({Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR0_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, SubCellInst_SboxInst_11_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR1_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, SubCellInst_SboxInst_11_XX_1_}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR3_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, SubCellInst_SboxInst_11_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR5_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR6_U1 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, SubCellInst_SboxInst_11_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR8_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, SubCellInst_SboxInst_11_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U1 ( .a ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .a ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .a ({Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR0_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, SubCellInst_SboxInst_12_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR1_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR3_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR5_U1 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_12_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR6_U1 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_12_Q6}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, SubCellInst_SboxInst_12_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR8_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, SubCellInst_SboxInst_12_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U1 ( .a ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .a ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, SubCellInst_SboxInst_13_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .a ({Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR0_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, SubCellInst_SboxInst_13_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR1_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, SubCellInst_SboxInst_13_XX_1_}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR3_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, SubCellInst_SboxInst_13_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR5_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR6_U1 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, SubCellInst_SboxInst_13_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR8_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, SubCellInst_SboxInst_13_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U1 ( .a ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .a ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .a ({Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR0_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, SubCellInst_SboxInst_14_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR1_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR3_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR5_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_14_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR6_U1 ( .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_14_Q6}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, SubCellInst_SboxInst_14_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR8_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, SubCellInst_SboxInst_14_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U1 ( .a ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .a ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, SubCellInst_SboxInst_15_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .a ({Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR0_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, SubCellInst_SboxInst_15_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR1_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, SubCellInst_SboxInst_15_XX_1_}), .c ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR3_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, SubCellInst_SboxInst_15_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR5_U1 ( .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR6_U1 ( .a ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, SubCellInst_SboxInst_15_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR8_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, SubCellInst_SboxInst_15_L2}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[0]}), .a ({Key_s2[0], Key_s1[0], Key_s0[0]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, TweakeyGeneration_StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[1]}), .a ({Key_s2[1], Key_s1[1], Key_s0[1]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, TweakeyGeneration_StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[2]}), .a ({Key_s2[2], Key_s1[2], Key_s0[2]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, TweakeyGeneration_StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[3]}), .a ({Key_s2[3], Key_s1[3], Key_s0[3]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, TweakeyGeneration_StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[4]}), .a ({Key_s2[4], Key_s1[4], Key_s0[4]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, TweakeyGeneration_StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[5]}), .a ({Key_s2[5], Key_s1[5], Key_s0[5]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, TweakeyGeneration_StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[6]}), .a ({Key_s2[6], Key_s1[6], Key_s0[6]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, TweakeyGeneration_StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[7]}), .a ({Key_s2[7], Key_s1[7], Key_s0[7]}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, TweakeyGeneration_StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[8]}), .a ({Key_s2[8], Key_s1[8], Key_s0[8]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, TweakeyGeneration_StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[9]}), .a ({Key_s2[9], Key_s1[9], Key_s0[9]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, TweakeyGeneration_StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[10]}), .a ({Key_s2[10], Key_s1[10], Key_s0[10]}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, TweakeyGeneration_StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[11]}), .a ({Key_s2[11], Key_s1[11], Key_s0[11]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, TweakeyGeneration_StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[12]}), .a ({Key_s2[12], Key_s1[12], Key_s0[12]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, TweakeyGeneration_StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[13]}), .a ({Key_s2[13], Key_s1[13], Key_s0[13]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, TweakeyGeneration_StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[14]}), .a ({Key_s2[14], Key_s1[14], Key_s0[14]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, TweakeyGeneration_StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[15]}), .a ({Key_s2[15], Key_s1[15], Key_s0[15]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, TweakeyGeneration_StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[16]}), .a ({Key_s2[16], Key_s1[16], Key_s0[16]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, TweakeyGeneration_StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_key_Feedback[17]}), .a ({Key_s2[17], Key_s1[17], Key_s0[17]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, TweakeyGeneration_StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, TweakeyGeneration_key_Feedback[18]}), .a ({Key_s2[18], Key_s1[18], Key_s0[18]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, TweakeyGeneration_StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[19]}), .a ({Key_s2[19], Key_s1[19], Key_s0[19]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, TweakeyGeneration_StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_key_Feedback[20]}), .a ({Key_s2[20], Key_s1[20], Key_s0[20]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, TweakeyGeneration_StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, TweakeyGeneration_key_Feedback[21]}), .a ({Key_s2[21], Key_s1[21], Key_s0[21]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, TweakeyGeneration_StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[22]}), .a ({Key_s2[22], Key_s1[22], Key_s0[22]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, TweakeyGeneration_StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_key_Feedback[23]}), .a ({Key_s2[23], Key_s1[23], Key_s0[23]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, TweakeyGeneration_StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, TweakeyGeneration_key_Feedback[24]}), .a ({Key_s2[24], Key_s1[24], Key_s0[24]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, TweakeyGeneration_StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[25]}), .a ({Key_s2[25], Key_s1[25], Key_s0[25]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, TweakeyGeneration_StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_key_Feedback[26]}), .a ({Key_s2[26], Key_s1[26], Key_s0[26]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, TweakeyGeneration_StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, TweakeyGeneration_key_Feedback[27]}), .a ({Key_s2[27], Key_s1[27], Key_s0[27]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, TweakeyGeneration_StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[28]}), .a ({Key_s2[28], Key_s1[28], Key_s0[28]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, TweakeyGeneration_StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_key_Feedback[29]}), .a ({Key_s2[29], Key_s1[29], Key_s0[29]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, TweakeyGeneration_StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, TweakeyGeneration_key_Feedback[30]}), .a ({Key_s2[30], Key_s1[30], Key_s0[30]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, TweakeyGeneration_StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[31]}), .a ({Key_s2[31], Key_s1[31], Key_s0[31]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, TweakeyGeneration_StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_key_Feedback[32]}), .a ({Key_s2[32], Key_s1[32], Key_s0[32]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, TweakeyGeneration_StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, TweakeyGeneration_key_Feedback[33]}), .a ({Key_s2[33], Key_s1[33], Key_s0[33]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, TweakeyGeneration_StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[34]}), .a ({Key_s2[34], Key_s1[34], Key_s0[34]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, TweakeyGeneration_StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_key_Feedback[35]}), .a ({Key_s2[35], Key_s1[35], Key_s0[35]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, TweakeyGeneration_StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, TweakeyGeneration_key_Feedback[36]}), .a ({Key_s2[36], Key_s1[36], Key_s0[36]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, TweakeyGeneration_StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[37]}), .a ({Key_s2[37], Key_s1[37], Key_s0[37]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, TweakeyGeneration_StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_key_Feedback[38]}), .a ({Key_s2[38], Key_s1[38], Key_s0[38]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, TweakeyGeneration_StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, TweakeyGeneration_key_Feedback[39]}), .a ({Key_s2[39], Key_s1[39], Key_s0[39]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, TweakeyGeneration_StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[40]}), .a ({Key_s2[40], Key_s1[40], Key_s0[40]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, TweakeyGeneration_StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_key_Feedback[41]}), .a ({Key_s2[41], Key_s1[41], Key_s0[41]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, TweakeyGeneration_StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, TweakeyGeneration_key_Feedback[42]}), .a ({Key_s2[42], Key_s1[42], Key_s0[42]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, TweakeyGeneration_StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[43]}), .a ({Key_s2[43], Key_s1[43], Key_s0[43]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, TweakeyGeneration_StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_key_Feedback[44]}), .a ({Key_s2[44], Key_s1[44], Key_s0[44]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, TweakeyGeneration_StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, TweakeyGeneration_key_Feedback[45]}), .a ({Key_s2[45], Key_s1[45], Key_s0[45]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, TweakeyGeneration_StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[46]}), .a ({Key_s2[46], Key_s1[46], Key_s0[46]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, TweakeyGeneration_StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_key_Feedback[47]}), .a ({Key_s2[47], Key_s1[47], Key_s0[47]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, TweakeyGeneration_StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, TweakeyGeneration_key_Feedback[48]}), .a ({Key_s2[48], Key_s1[48], Key_s0[48]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, TweakeyGeneration_StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[49]}), .a ({Key_s2[49], Key_s1[49], Key_s0[49]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, TweakeyGeneration_StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_key_Feedback[50]}), .a ({Key_s2[50], Key_s1[50], Key_s0[50]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, TweakeyGeneration_StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, TweakeyGeneration_key_Feedback[51]}), .a ({Key_s2[51], Key_s1[51], Key_s0[51]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, TweakeyGeneration_StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[52]}), .a ({Key_s2[52], Key_s1[52], Key_s0[52]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, TweakeyGeneration_StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_key_Feedback[53]}), .a ({Key_s2[53], Key_s1[53], Key_s0[53]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, TweakeyGeneration_StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, TweakeyGeneration_key_Feedback[54]}), .a ({Key_s2[54], Key_s1[54], Key_s0[54]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, TweakeyGeneration_StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[55]}), .a ({Key_s2[55], Key_s1[55], Key_s0[55]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, TweakeyGeneration_StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_key_Feedback[56]}), .a ({Key_s2[56], Key_s1[56], Key_s0[56]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, TweakeyGeneration_StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, TweakeyGeneration_key_Feedback[57]}), .a ({Key_s2[57], Key_s1[57], Key_s0[57]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, TweakeyGeneration_StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[58]}), .a ({Key_s2[58], Key_s1[58], Key_s0[58]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, TweakeyGeneration_StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_key_Feedback[59]}), .a ({Key_s2[59], Key_s1[59], Key_s0[59]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, TweakeyGeneration_StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, TweakeyGeneration_key_Feedback[60]}), .a ({Key_s2[60], Key_s1[60], Key_s0[60]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, TweakeyGeneration_StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[61]}), .a ({Key_s2[61], Key_s1[61], Key_s0[61]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, TweakeyGeneration_StateRegInput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_key_Feedback[62]}), .a ({Key_s2[62], Key_s1[62], Key_s0[62]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, TweakeyGeneration_StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, TweakeyGeneration_key_Feedback[63]}), .a ({Key_s2[63], Key_s1[63], Key_s0[63]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, TweakeyGeneration_StateRegInput[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMUpdate[0]), .B (1'b1), .Z (FSMSelected[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMUpdate[1]), .B (1'b0), .Z (FSMSelected[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMUpdate[2]), .B (1'b0), .Z (FSMSelected[2]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMUpdate[3]), .B (1'b0), .Z (FSMSelected[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMUpdate[4]), .B (1'b0), .Z (FSMSelected[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMUpdate[5]), .B (1'b0), .Z (FSMSelected[5]) ) ;
    MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .S (FSM[4]), .A (FSMUpdateInst_StateUpdateInst_0_n4), .B (FSM[5]), .Z (FSMUpdate[0]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_0_n3), .ZN (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1 (FSMUpdateInst_StateUpdateInst_0_n2), .A2 (FSMUpdateInst_StateUpdateInst_0_n1), .ZN (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n4), .A2 (FSM[1]), .ZN (FSMUpdate[2]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n3), .A2 (FSM[5]), .ZN (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_2_n2), .ZN (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1 (FSMUpdate[1]), .A2 (FSMUpdateInst_StateUpdateInst_2_n1), .ZN (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n4), .ZN (FSMUpdate[5]) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1 (FSMUpdate[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n3), .ZN (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_5_n2), .ZN (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdateInst_StateUpdateInst_5_n1), .ZN (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1 (FSMSignalsInst_doneInst_n5), .A2 (FSMSignalsInst_doneInst_n4), .ZN (done) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1 (FSM[4]), .A2 (FSM[5]), .ZN (FSMSignalsInst_doneInst_n4) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1 (FSMSignalsInst_doneInst_n3), .A2 (FSMSignalsInst_doneInst_n2), .ZN (FSMSignalsInst_doneInst_n5) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1 (FSMUpdate[4]), .A2 (FSMSignalsInst_doneInst_n1), .ZN (FSMSignalsInst_doneInst_n2) ) ;
    INV_X1 FSMSignalsInst_doneInst_U2 ( .A (FSMUpdate[1]), .ZN (FSMSignalsInst_doneInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1 (FSM[1]), .A2 (FSMUpdate[3]), .ZN (FSMSignalsInst_doneInst_n3) ) ;

    /* cells in depth 1 */
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_2_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, MCOutput[2]}), .a ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_3_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[3]}), .a ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_6_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, MCOutput[6]}), .a ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_7_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, MCOutput[7]}), .a ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_10_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, MCOutput[10]}), .a ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_11_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, MCOutput[11]}), .a ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_14_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, MCOutput[14]}), .a ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, new_AGEMA_signal_3489}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_15_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCOutput[15]}), .a ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_18_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, MCOutput[18]}), .a ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_19_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, MCOutput[19]}), .a ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_22_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, MCOutput[22]}), .a ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_23_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, MCOutput[23]}), .a ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_26_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[26]}), .a ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_27_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCOutput[27]}), .a ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_30_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, MCOutput[30]}), .a ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_31_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, MCOutput[31]}), .a ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_34_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .a ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_35_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .a ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_38_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .a ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_39_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .a ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_42_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_43_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .a ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_46_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .a ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_47_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .a ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_50_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, MCOutput[50]}), .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_51_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[51]}), .a ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_54_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, MCOutput[54]}), .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_55_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[55]}), .a ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_58_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, MCOutput[58]}), .a ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_59_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, MCOutput[59]}), .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_62_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[62]}), .a ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_63_U1 ( .s (new_AGEMA_signal_3470), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCOutput[63]}), .a ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564}), .c ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, StateRegInput[63]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, ShiftRowsOutput[7]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_U2 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_YY_0_}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, ShiftRowsOutput[6]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_AND1_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR2_U1 ( .a ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_AND3_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR7_U1 ( .a ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR11_U1 ( .a ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, SubCellInst_SboxInst_0_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR12_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, SubCellInst_SboxInst_0_L3}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, SubCellInst_SboxInst_0_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR13_U1 ( .a ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, ShiftRowsOutput[11]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_U2 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_1_YY_0_}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, ShiftRowsOutput[10]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_AND1_U1 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR2_U1 ( .a ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_1_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_AND3_U1 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, SubCellInst_SboxInst_1_Q4}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR7_U1 ( .a ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, SubCellInst_SboxInst_1_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR11_U1 ( .a ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR12_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, SubCellInst_SboxInst_1_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR13_U1 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_1_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, ShiftRowsOutput[15]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_U2 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, SubCellInst_SboxInst_2_YY_0_}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, ShiftRowsOutput[14]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_AND1_U1 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR2_U1 ( .a ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_AND3_U1 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR7_U1 ( .a ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR11_U1 ( .a ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_2_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR12_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_2_L3}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_2_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR13_U1 ( .a ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, SubCellInst_SboxInst_2_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, ShiftRowsOutput[3]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_U2 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_3_YY_0_}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, ShiftRowsOutput[2]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_AND1_U1 ( .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR2_U1 ( .a ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_3_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_AND3_U1 ( .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, SubCellInst_SboxInst_3_Q4}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR7_U1 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_3_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR11_U1 ( .a ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR12_U1 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, SubCellInst_SboxInst_3_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR13_U1 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_3_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_U2 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_4_YY_0_}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_AND1_U1 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR2_U1 ( .a ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_AND3_U1 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR7_U1 ( .a ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR11_U1 ( .a ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, SubCellInst_SboxInst_4_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR12_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, SubCellInst_SboxInst_4_L3}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, SubCellInst_SboxInst_4_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR13_U1 ( .a ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_4_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_U2 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, SubCellInst_SboxInst_5_YY_0_}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_AND1_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR2_U1 ( .a ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, SubCellInst_SboxInst_5_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_AND3_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, SubCellInst_SboxInst_5_Q4}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR7_U1 ( .a ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_5_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR11_U1 ( .a ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR12_U1 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_5_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR13_U1 ( .a ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, SubCellInst_SboxInst_5_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_U2 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, SubCellInst_SboxInst_6_YY_0_}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_AND1_U1 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR2_U1 ( .a ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_AND3_U1 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR7_U1 ( .a ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR11_U1 ( .a ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, SubCellInst_SboxInst_6_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR12_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, SubCellInst_SboxInst_6_L3}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, SubCellInst_SboxInst_6_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR13_U1 ( .a ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, SubCellInst_SboxInst_6_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_U2 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, SubCellInst_SboxInst_7_YY_0_}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_AND1_U1 ( .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR2_U1 ( .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, SubCellInst_SboxInst_7_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_AND3_U1 ( .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, SubCellInst_SboxInst_7_Q4}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR7_U1 ( .a ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, SubCellInst_SboxInst_7_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR11_U1 ( .a ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR12_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, SubCellInst_SboxInst_7_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR13_U1 ( .a ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, SubCellInst_SboxInst_7_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, AddRoundConstantOutput[35]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_U2 ( .a ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, SubCellInst_SboxInst_8_YY_0_}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, AddRoundConstantOutput[34]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_AND1_U1 ( .a ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR2_U1 ( .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_AND3_U1 ( .a ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR7_U1 ( .a ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR11_U1 ( .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, SubCellInst_SboxInst_8_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR12_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, SubCellInst_SboxInst_8_L3}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, SubCellInst_SboxInst_8_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR13_U1 ( .a ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, SubCellInst_SboxInst_8_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, AddRoundConstantOutput[39]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_U2 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_9_YY_0_}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, AddRoundConstantOutput[38]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_AND1_U1 ( .a ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR2_U1 ( .a ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, SubCellInst_SboxInst_9_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_AND3_U1 ( .a ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, SubCellInst_SboxInst_9_Q4}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR7_U1 ( .a ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, SubCellInst_SboxInst_9_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR11_U1 ( .a ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR12_U1 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, SubCellInst_SboxInst_9_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR13_U1 ( .a ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_9_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, AddRoundConstantOutput[43]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_U2 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, SubCellInst_SboxInst_10_YY_0_}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, AddRoundConstantOutput[42]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_AND1_U1 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR2_U1 ( .a ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_AND3_U1 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR7_U1 ( .a ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR11_U1 ( .a ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_10_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR12_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_10_L3}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, SubCellInst_SboxInst_10_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR13_U1 ( .a ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, SubCellInst_SboxInst_10_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellOutput[47]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_U2 ( .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, SubCellInst_SboxInst_11_YY_0_}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, SubCellOutput[46]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_AND1_U1 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR2_U1 ( .a ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_AND3_U1 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, SubCellInst_SboxInst_11_Q4}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR7_U1 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR11_U1 ( .a ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, SubCellInst_SboxInst_11_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR12_U1 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, SubCellInst_SboxInst_11_L3}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_11_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR13_U1 ( .a ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, SubCellInst_SboxInst_11_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, AddRoundConstantOutput[51]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_U2 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_12_YY_0_}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, AddRoundConstantOutput[50]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_AND1_U1 ( .a ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR2_U1 ( .a ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_12_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_AND3_U1 ( .a ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR7_U1 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, SubCellInst_SboxInst_12_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR11_U1 ( .a ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR12_U1 ( .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, SubCellInst_SboxInst_12_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR13_U1 ( .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_12_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, AddRoundConstantOutput[55]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_U2 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, SubCellInst_SboxInst_13_YY_0_}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, AddRoundConstantOutput[54]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_AND1_U1 ( .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR2_U1 ( .a ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_AND3_U1 ( .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, SubCellInst_SboxInst_13_Q4}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR7_U1 ( .a ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR11_U1 ( .a ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, new_AGEMA_signal_3729}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, SubCellInst_SboxInst_13_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR12_U1 ( .a ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, SubCellInst_SboxInst_13_L3}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, SubCellInst_SboxInst_13_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR13_U1 ( .a ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, new_AGEMA_signal_3732}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, SubCellInst_SboxInst_13_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, AddRoundConstantOutput[59]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_U2 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, SubCellInst_SboxInst_14_YY_0_}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, AddRoundConstantOutput[58]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_AND1_U1 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR2_U1 ( .a ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, SubCellInst_SboxInst_14_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_AND3_U1 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR7_U1 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_14_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR11_U1 ( .a ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, new_AGEMA_signal_3741}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR12_U1 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_14_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR13_U1 ( .a ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, new_AGEMA_signal_3744}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, SubCellInst_SboxInst_14_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, SubCellOutput[63]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_U2 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, SubCellInst_SboxInst_15_YY_0_}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, SubCellOutput[62]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_AND1_U1 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR2_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_AND3_U1 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, SubCellInst_SboxInst_15_Q4}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR7_U1 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR11_U1 ( .a ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, new_AGEMA_signal_3753}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, SubCellInst_SboxInst_15_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR12_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, SubCellInst_SboxInst_15_L3}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, SubCellInst_SboxInst_15_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR13_U1 ( .a ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, new_AGEMA_signal_3756}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, SubCellInst_SboxInst_15_YY_0_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, AddConstXOR_AddConstXOR_XORInst_0_2_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_3759}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, AddRoundConstantOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, SubCellOutput[62]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, AddConstXOR_AddConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, AddConstXOR_AddConstXOR_XORInst_0_3_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_3760}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, AddRoundConstantOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, SubCellOutput[63]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, AddConstXOR_AddConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, AddConstXOR_AddConstXOR_XORInst_1_2_n1}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, AddRoundConstantOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, SubCellOutput[46]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, AddConstXOR_AddConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, AddConstXOR_AddConstXOR_XORInst_1_3_n1}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, AddRoundConstantOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellOutput[47]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, AddConstXOR_AddConstXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, AddRoundTweakeyXOR_XORInst_0_2_n1}), .b ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, new_AGEMA_signal_3761}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, AddRoundConstantOutput[34]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, AddRoundTweakeyXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, AddRoundTweakeyXOR_XORInst_0_3_n1}), .b ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, new_AGEMA_signal_3764}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, ShiftRowsOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, AddRoundConstantOutput[35]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, AddRoundTweakeyXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, AddRoundTweakeyXOR_XORInst_1_2_n1}), .b ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, new_AGEMA_signal_3767}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, ShiftRowsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, AddRoundConstantOutput[38]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, AddRoundTweakeyXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, AddRoundTweakeyXOR_XORInst_1_3_n1}), .b ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, AddRoundConstantOutput[39]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, AddRoundTweakeyXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, AddRoundTweakeyXOR_XORInst_2_2_n1}), .b ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, new_AGEMA_signal_3773}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, AddRoundConstantOutput[42]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, AddRoundTweakeyXOR_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, AddRoundTweakeyXOR_XORInst_2_3_n1}), .b ({new_AGEMA_signal_3778, new_AGEMA_signal_3777, new_AGEMA_signal_3776}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, ShiftRowsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, AddRoundConstantOutput[43]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, AddRoundTweakeyXOR_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, AddRoundTweakeyXOR_XORInst_3_2_n1}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, ShiftRowsOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, AddRoundConstantOutput[46]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, AddRoundTweakeyXOR_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, AddRoundTweakeyXOR_XORInst_3_3_n1}), .b ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, new_AGEMA_signal_3782}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, ShiftRowsOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, AddRoundConstantOutput[47]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, AddRoundTweakeyXOR_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1}), .b ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, new_AGEMA_signal_3785}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, AddRoundConstantOutput[50]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, AddRoundTweakeyXOR_XORInst_4_3_n1}), .b ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, new_AGEMA_signal_3788}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, AddRoundConstantOutput[51]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, AddRoundTweakeyXOR_XORInst_4_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_3791}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, AddRoundConstantOutput[54]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, AddRoundTweakeyXOR_XORInst_5_3_n1}), .b ({new_AGEMA_signal_3796, new_AGEMA_signal_3795, new_AGEMA_signal_3794}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, AddRoundConstantOutput[55]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, AddRoundTweakeyXOR_XORInst_5_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, new_AGEMA_signal_3797}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, AddRoundConstantOutput[58]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, AddRoundTweakeyXOR_XORInst_6_3_n1}), .b ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, new_AGEMA_signal_3800}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, AddRoundConstantOutput[59]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, AddRoundTweakeyXOR_XORInst_6_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1}), .b ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, new_AGEMA_signal_3803}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, AddRoundConstantOutput[62]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, AddRoundTweakeyXOR_XORInst_7_3_n1}), .b ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, AddRoundConstantOutput[63]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, AddRoundTweakeyXOR_XORInst_7_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, MCInst_MCR0_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, MCOutput[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, MCInst_MCR0_XORInst_0_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, MCInst_MCR0_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[51]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, MCInst_MCR0_XORInst_0_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, MCInst_MCR0_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, MCOutput[54]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, MCInst_MCR0_XORInst_1_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, MCInst_MCR0_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[55]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .b ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, MCInst_MCR0_XORInst_1_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U3 ( .a ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, MCInst_MCR0_XORInst_2_2_n2}), .b ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, MCOutput[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, MCInst_MCR0_XORInst_2_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U3 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, MCInst_MCR0_XORInst_2_3_n2}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, MCOutput[59]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, MCInst_MCR0_XORInst_2_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U3 ( .a ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCInst_MCR0_XORInst_3_2_n2}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCInst_MCR0_XORInst_3_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U3 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, MCInst_MCR0_XORInst_3_3_n2}), .b ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, MCInst_MCR0_XORInst_3_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, MCOutput[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, MCInst_MCR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, MCOutput[19]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, MCInst_MCR2_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, MCOutput[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, MCInst_MCR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, MCOutput[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, MCInst_MCR2_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, MCInst_MCR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCOutput[27]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, MCInst_MCR2_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, MCOutput[30]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, MCInst_MCR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, MCOutput[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, MCInst_MCR2_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, MCOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, MCInst_MCR3_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, MCInst_MCR3_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, MCOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, MCInst_MCR3_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, MCOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, MCInst_MCR3_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, MCOutput[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, MCInst_MCR3_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, MCOutput[11]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, MCInst_MCR3_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, MCOutput[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, MCInst_MCR3_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCOutput[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, MCInst_MCR3_XORInst_3_3_n1}) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (rst), .Q (new_AGEMA_signal_3470) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (Plaintext_s0[2]), .Q (new_AGEMA_signal_3471) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (Plaintext_s1[2]), .Q (new_AGEMA_signal_3472) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (Plaintext_s2[2]), .Q (new_AGEMA_signal_3473) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (Plaintext_s0[3]), .Q (new_AGEMA_signal_3474) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (Plaintext_s1[3]), .Q (new_AGEMA_signal_3475) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (Plaintext_s2[3]), .Q (new_AGEMA_signal_3476) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (Plaintext_s0[6]), .Q (new_AGEMA_signal_3477) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (Plaintext_s1[6]), .Q (new_AGEMA_signal_3478) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (Plaintext_s2[6]), .Q (new_AGEMA_signal_3479) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (Plaintext_s0[7]), .Q (new_AGEMA_signal_3480) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (Plaintext_s1[7]), .Q (new_AGEMA_signal_3481) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (Plaintext_s2[7]), .Q (new_AGEMA_signal_3482) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (Plaintext_s0[10]), .Q (new_AGEMA_signal_3483) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (Plaintext_s1[10]), .Q (new_AGEMA_signal_3484) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (Plaintext_s2[10]), .Q (new_AGEMA_signal_3485) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (Plaintext_s0[11]), .Q (new_AGEMA_signal_3486) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (Plaintext_s1[11]), .Q (new_AGEMA_signal_3487) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (Plaintext_s2[11]), .Q (new_AGEMA_signal_3488) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (Plaintext_s0[14]), .Q (new_AGEMA_signal_3489) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (Plaintext_s1[14]), .Q (new_AGEMA_signal_3490) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (Plaintext_s2[14]), .Q (new_AGEMA_signal_3491) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (Plaintext_s0[15]), .Q (new_AGEMA_signal_3492) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (Plaintext_s1[15]), .Q (new_AGEMA_signal_3493) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (Plaintext_s2[15]), .Q (new_AGEMA_signal_3494) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (Plaintext_s0[18]), .Q (new_AGEMA_signal_3495) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (Plaintext_s1[18]), .Q (new_AGEMA_signal_3496) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (Plaintext_s2[18]), .Q (new_AGEMA_signal_3497) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (Plaintext_s0[19]), .Q (new_AGEMA_signal_3498) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (Plaintext_s1[19]), .Q (new_AGEMA_signal_3499) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (Plaintext_s2[19]), .Q (new_AGEMA_signal_3500) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (Plaintext_s0[22]), .Q (new_AGEMA_signal_3501) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (Plaintext_s1[22]), .Q (new_AGEMA_signal_3502) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (Plaintext_s2[22]), .Q (new_AGEMA_signal_3503) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (Plaintext_s0[23]), .Q (new_AGEMA_signal_3504) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (Plaintext_s1[23]), .Q (new_AGEMA_signal_3505) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (Plaintext_s2[23]), .Q (new_AGEMA_signal_3506) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (Plaintext_s0[26]), .Q (new_AGEMA_signal_3507) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (Plaintext_s1[26]), .Q (new_AGEMA_signal_3508) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (Plaintext_s2[26]), .Q (new_AGEMA_signal_3509) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (Plaintext_s0[27]), .Q (new_AGEMA_signal_3510) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (Plaintext_s1[27]), .Q (new_AGEMA_signal_3511) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (Plaintext_s2[27]), .Q (new_AGEMA_signal_3512) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (Plaintext_s0[30]), .Q (new_AGEMA_signal_3513) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (Plaintext_s1[30]), .Q (new_AGEMA_signal_3514) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (Plaintext_s2[30]), .Q (new_AGEMA_signal_3515) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (Plaintext_s0[31]), .Q (new_AGEMA_signal_3516) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (Plaintext_s1[31]), .Q (new_AGEMA_signal_3517) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (Plaintext_s2[31]), .Q (new_AGEMA_signal_3518) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (Plaintext_s0[34]), .Q (new_AGEMA_signal_3519) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (Plaintext_s1[34]), .Q (new_AGEMA_signal_3520) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (Plaintext_s2[34]), .Q (new_AGEMA_signal_3521) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (Plaintext_s0[35]), .Q (new_AGEMA_signal_3522) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (Plaintext_s1[35]), .Q (new_AGEMA_signal_3523) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (Plaintext_s2[35]), .Q (new_AGEMA_signal_3524) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (Plaintext_s0[38]), .Q (new_AGEMA_signal_3525) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (Plaintext_s1[38]), .Q (new_AGEMA_signal_3526) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (Plaintext_s2[38]), .Q (new_AGEMA_signal_3527) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (Plaintext_s0[39]), .Q (new_AGEMA_signal_3528) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (Plaintext_s1[39]), .Q (new_AGEMA_signal_3529) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (Plaintext_s2[39]), .Q (new_AGEMA_signal_3530) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (Plaintext_s0[42]), .Q (new_AGEMA_signal_3531) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (Plaintext_s1[42]), .Q (new_AGEMA_signal_3532) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (Plaintext_s2[42]), .Q (new_AGEMA_signal_3533) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (Plaintext_s0[43]), .Q (new_AGEMA_signal_3534) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (Plaintext_s1[43]), .Q (new_AGEMA_signal_3535) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (Plaintext_s2[43]), .Q (new_AGEMA_signal_3536) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (Plaintext_s0[46]), .Q (new_AGEMA_signal_3537) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (Plaintext_s1[46]), .Q (new_AGEMA_signal_3538) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (Plaintext_s2[46]), .Q (new_AGEMA_signal_3539) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (Plaintext_s0[47]), .Q (new_AGEMA_signal_3540) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (Plaintext_s1[47]), .Q (new_AGEMA_signal_3541) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (Plaintext_s2[47]), .Q (new_AGEMA_signal_3542) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (Plaintext_s0[50]), .Q (new_AGEMA_signal_3543) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (Plaintext_s1[50]), .Q (new_AGEMA_signal_3544) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (Plaintext_s2[50]), .Q (new_AGEMA_signal_3545) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (Plaintext_s0[51]), .Q (new_AGEMA_signal_3546) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (Plaintext_s1[51]), .Q (new_AGEMA_signal_3547) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (Plaintext_s2[51]), .Q (new_AGEMA_signal_3548) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (Plaintext_s0[54]), .Q (new_AGEMA_signal_3549) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (Plaintext_s1[54]), .Q (new_AGEMA_signal_3550) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (Plaintext_s2[54]), .Q (new_AGEMA_signal_3551) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (Plaintext_s0[55]), .Q (new_AGEMA_signal_3552) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (Plaintext_s1[55]), .Q (new_AGEMA_signal_3553) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (Plaintext_s2[55]), .Q (new_AGEMA_signal_3554) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (Plaintext_s0[58]), .Q (new_AGEMA_signal_3555) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (Plaintext_s1[58]), .Q (new_AGEMA_signal_3556) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (Plaintext_s2[58]), .Q (new_AGEMA_signal_3557) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (Plaintext_s0[59]), .Q (new_AGEMA_signal_3558) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (Plaintext_s1[59]), .Q (new_AGEMA_signal_3559) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (Plaintext_s2[59]), .Q (new_AGEMA_signal_3560) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (Plaintext_s0[62]), .Q (new_AGEMA_signal_3561) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (Plaintext_s1[62]), .Q (new_AGEMA_signal_3562) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (Plaintext_s2[62]), .Q (new_AGEMA_signal_3563) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (Plaintext_s0[63]), .Q (new_AGEMA_signal_3564) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (Plaintext_s1[63]), .Q (new_AGEMA_signal_3565) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (Plaintext_s2[63]), .Q (new_AGEMA_signal_3566) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (SubCellInst_SboxInst_0_Q0), .Q (new_AGEMA_signal_3567) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (new_AGEMA_signal_1742), .Q (new_AGEMA_signal_3568) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (new_AGEMA_signal_1743), .Q (new_AGEMA_signal_3569) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (SubCellInst_SboxInst_0_L1), .Q (new_AGEMA_signal_3570) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (new_AGEMA_signal_1936), .Q (new_AGEMA_signal_3571) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (new_AGEMA_signal_1937), .Q (new_AGEMA_signal_3572) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (SubCellInst_SboxInst_0_XX_2_), .Q (new_AGEMA_signal_3573) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (new_AGEMA_signal_1174), .Q (new_AGEMA_signal_3574) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (new_AGEMA_signal_1175), .Q (new_AGEMA_signal_3575) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (SubCellInst_SboxInst_0_XX_1_), .Q (new_AGEMA_signal_3576) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (new_AGEMA_signal_1170), .Q (new_AGEMA_signal_3577) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (new_AGEMA_signal_1171), .Q (new_AGEMA_signal_3578) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (SubCellInst_SboxInst_1_Q0), .Q (new_AGEMA_signal_3579) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (new_AGEMA_signal_1754), .Q (new_AGEMA_signal_3580) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (new_AGEMA_signal_1755), .Q (new_AGEMA_signal_3581) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (SubCellInst_SboxInst_1_L1), .Q (new_AGEMA_signal_3582) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (new_AGEMA_signal_1942), .Q (new_AGEMA_signal_3583) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (new_AGEMA_signal_1943), .Q (new_AGEMA_signal_3584) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (SubCellInst_SboxInst_1_XX_2_), .Q (new_AGEMA_signal_3585) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (new_AGEMA_signal_1186), .Q (new_AGEMA_signal_3586) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (new_AGEMA_signal_1187), .Q (new_AGEMA_signal_3587) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (SubCellInst_SboxInst_1_XX_1_), .Q (new_AGEMA_signal_3588) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (new_AGEMA_signal_1182), .Q (new_AGEMA_signal_3589) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (new_AGEMA_signal_1183), .Q (new_AGEMA_signal_3590) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (SubCellInst_SboxInst_2_Q0), .Q (new_AGEMA_signal_3591) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_3592) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (new_AGEMA_signal_1767), .Q (new_AGEMA_signal_3593) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (SubCellInst_SboxInst_2_L1), .Q (new_AGEMA_signal_3594) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (new_AGEMA_signal_1948), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (new_AGEMA_signal_1949), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (SubCellInst_SboxInst_2_XX_2_), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (new_AGEMA_signal_1198), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (new_AGEMA_signal_1199), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (SubCellInst_SboxInst_2_XX_1_), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (new_AGEMA_signal_1195), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (SubCellInst_SboxInst_3_Q0), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (new_AGEMA_signal_1779), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (SubCellInst_SboxInst_3_L1), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (new_AGEMA_signal_1954), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (new_AGEMA_signal_1955), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (SubCellInst_SboxInst_3_XX_2_), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (new_AGEMA_signal_1210), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (new_AGEMA_signal_1211), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (SubCellInst_SboxInst_3_XX_1_), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (new_AGEMA_signal_1207), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (SubCellInst_SboxInst_4_Q0), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (new_AGEMA_signal_1791), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (SubCellInst_SboxInst_4_L1), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (new_AGEMA_signal_1960), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (new_AGEMA_signal_1961), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (SubCellInst_SboxInst_4_XX_2_), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (new_AGEMA_signal_1222), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (new_AGEMA_signal_1223), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (SubCellInst_SboxInst_4_XX_1_), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (new_AGEMA_signal_1218), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (new_AGEMA_signal_1219), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (SubCellInst_SboxInst_5_Q0), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (new_AGEMA_signal_1803), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (SubCellInst_SboxInst_5_L1), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (new_AGEMA_signal_1966), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (new_AGEMA_signal_1967), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (SubCellInst_SboxInst_5_XX_2_), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (new_AGEMA_signal_1234), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (new_AGEMA_signal_1235), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (SubCellInst_SboxInst_5_XX_1_), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (new_AGEMA_signal_1230), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (new_AGEMA_signal_1231), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (SubCellInst_SboxInst_6_Q0), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (new_AGEMA_signal_1815), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (SubCellInst_SboxInst_6_L1), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (new_AGEMA_signal_1973), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (SubCellInst_SboxInst_6_XX_2_), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (new_AGEMA_signal_1246), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (new_AGEMA_signal_1247), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (SubCellInst_SboxInst_6_XX_1_), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (new_AGEMA_signal_1243), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (SubCellInst_SboxInst_7_Q0), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (new_AGEMA_signal_1827), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (SubCellInst_SboxInst_7_L1), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (new_AGEMA_signal_1978), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (new_AGEMA_signal_1979), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (SubCellInst_SboxInst_7_XX_2_), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (new_AGEMA_signal_1258), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (new_AGEMA_signal_1259), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (SubCellInst_SboxInst_7_XX_1_), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (new_AGEMA_signal_1255), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (SubCellInst_SboxInst_8_Q0), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (new_AGEMA_signal_1839), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (SubCellInst_SboxInst_8_L1), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (new_AGEMA_signal_1984), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (new_AGEMA_signal_1985), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (SubCellInst_SboxInst_8_XX_2_), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (new_AGEMA_signal_1270), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (new_AGEMA_signal_1271), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (SubCellInst_SboxInst_8_XX_1_), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (new_AGEMA_signal_1266), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (new_AGEMA_signal_1267), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (SubCellInst_SboxInst_9_Q0), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (new_AGEMA_signal_1850), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (new_AGEMA_signal_1851), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (SubCellInst_SboxInst_9_L1), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (new_AGEMA_signal_1991), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (SubCellInst_SboxInst_9_XX_2_), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (new_AGEMA_signal_1282), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (new_AGEMA_signal_1283), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (SubCellInst_SboxInst_9_XX_1_), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (new_AGEMA_signal_1279), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (SubCellInst_SboxInst_10_Q0), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (new_AGEMA_signal_1863), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (SubCellInst_SboxInst_10_L1), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (new_AGEMA_signal_1996), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (new_AGEMA_signal_1997), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (SubCellInst_SboxInst_10_XX_2_), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (new_AGEMA_signal_1294), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (new_AGEMA_signal_1295), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (SubCellInst_SboxInst_10_XX_1_), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (new_AGEMA_signal_1291), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (SubCellInst_SboxInst_11_Q0), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (new_AGEMA_signal_1875), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (SubCellInst_SboxInst_11_L1), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (new_AGEMA_signal_2002), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (new_AGEMA_signal_2003), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (SubCellInst_SboxInst_11_XX_2_), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (new_AGEMA_signal_1306), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (new_AGEMA_signal_1307), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (SubCellInst_SboxInst_11_XX_1_), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (new_AGEMA_signal_1302), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (new_AGEMA_signal_1303), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (SubCellInst_SboxInst_12_Q0), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (new_AGEMA_signal_1886), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (new_AGEMA_signal_1887), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (SubCellInst_SboxInst_12_L1), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (new_AGEMA_signal_2009), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (SubCellInst_SboxInst_12_XX_2_), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (new_AGEMA_signal_1318), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (new_AGEMA_signal_1319), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (SubCellInst_SboxInst_12_XX_1_), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (new_AGEMA_signal_1314), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (new_AGEMA_signal_1315), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (SubCellInst_SboxInst_13_Q0), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_1899), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (SubCellInst_SboxInst_13_L1), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_2014), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_2015), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (SubCellInst_SboxInst_13_XX_2_), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_1330), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_1331), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (SubCellInst_SboxInst_13_XX_1_), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_1326), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_1327), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (SubCellInst_SboxInst_14_Q0), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_1911), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (SubCellInst_SboxInst_14_L1), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_2021), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (SubCellInst_SboxInst_14_XX_2_), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_1342), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_1343), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (SubCellInst_SboxInst_14_XX_1_), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_1338), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_1339), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (SubCellInst_SboxInst_15_Q0), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_1923), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (SubCellInst_SboxInst_15_L1), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (SubCellInst_SboxInst_15_XX_2_), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_1354), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_1355), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (SubCellInst_SboxInst_15_XX_1_), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_1350), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_1351), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (FSMUpdate[3]), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (FSMUpdate[4]), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (TweakeyGeneration_key_Feedback[2]), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_1368), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_1369), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (TweakeyGeneration_key_Feedback[3]), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_1374), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_1375), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (TweakeyGeneration_key_Feedback[6]), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_1392), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_1393), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (TweakeyGeneration_key_Feedback[7]), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_1398), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_1399), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (TweakeyGeneration_key_Feedback[10]), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_1416), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_1417), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (TweakeyGeneration_key_Feedback[11]), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_1422), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_1423), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (TweakeyGeneration_key_Feedback[14]), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_1441), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (TweakeyGeneration_key_Feedback[15]), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_1447), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (TweakeyGeneration_key_Feedback[18]), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_1464), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_1465), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (TweakeyGeneration_key_Feedback[19]), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_1471), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (TweakeyGeneration_key_Feedback[22]), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_1489), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (TweakeyGeneration_key_Feedback[23]), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_1495), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (TweakeyGeneration_key_Feedback[26]), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_1513), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (TweakeyGeneration_key_Feedback[27]), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_1519), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (TweakeyGeneration_key_Feedback[30]), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_1536), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_1537), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (TweakeyGeneration_key_Feedback[31]), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_1542), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_1543), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (Plaintext_s0[0]), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (Plaintext_s1[0]), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (Plaintext_s2[0]), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (Plaintext_s0[1]), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (Plaintext_s1[1]), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (Plaintext_s2[1]), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (Plaintext_s0[4]), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (Plaintext_s1[4]), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (Plaintext_s2[4]), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (Plaintext_s0[5]), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (Plaintext_s1[5]), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (Plaintext_s2[5]), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (Plaintext_s0[8]), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (Plaintext_s1[8]), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (Plaintext_s2[8]), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (Plaintext_s0[9]), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (Plaintext_s1[9]), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (Plaintext_s2[9]), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (Plaintext_s0[12]), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (Plaintext_s1[12]), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (Plaintext_s2[12]), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (Plaintext_s0[13]), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (Plaintext_s1[13]), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (Plaintext_s2[13]), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (Plaintext_s0[16]), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (Plaintext_s1[16]), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (Plaintext_s2[16]), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (Plaintext_s0[17]), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (Plaintext_s1[17]), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (Plaintext_s2[17]), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (Plaintext_s0[20]), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (Plaintext_s1[20]), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (Plaintext_s2[20]), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (Plaintext_s0[21]), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (Plaintext_s1[21]), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (Plaintext_s2[21]), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (Plaintext_s0[24]), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (Plaintext_s1[24]), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (Plaintext_s2[24]), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (Plaintext_s0[25]), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (Plaintext_s1[25]), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (Plaintext_s2[25]), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (Plaintext_s0[28]), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (Plaintext_s1[28]), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (Plaintext_s2[28]), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (Plaintext_s0[29]), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (Plaintext_s1[29]), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (Plaintext_s2[29]), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (Plaintext_s0[32]), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (Plaintext_s1[32]), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (Plaintext_s2[32]), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (Plaintext_s0[33]), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (Plaintext_s1[33]), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (Plaintext_s2[33]), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (Plaintext_s0[36]), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (Plaintext_s1[36]), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (Plaintext_s2[36]), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (Plaintext_s0[37]), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (Plaintext_s1[37]), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (Plaintext_s2[37]), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (Plaintext_s0[40]), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (Plaintext_s1[40]), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (Plaintext_s2[40]), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (Plaintext_s0[41]), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (Plaintext_s1[41]), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (Plaintext_s2[41]), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (Plaintext_s0[44]), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (Plaintext_s1[44]), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (Plaintext_s2[44]), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (Plaintext_s0[45]), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (Plaintext_s1[45]), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (Plaintext_s2[45]), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (Plaintext_s0[48]), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (Plaintext_s1[48]), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (Plaintext_s2[48]), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (Plaintext_s0[49]), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (Plaintext_s1[49]), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (Plaintext_s2[49]), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (Plaintext_s0[52]), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (Plaintext_s1[52]), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (Plaintext_s2[52]), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (Plaintext_s0[53]), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (Plaintext_s1[53]), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (Plaintext_s2[53]), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (Plaintext_s0[56]), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (Plaintext_s1[56]), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (Plaintext_s2[56]), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (Plaintext_s0[57]), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (Plaintext_s1[57]), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (Plaintext_s2[57]), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (Plaintext_s0[60]), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (Plaintext_s1[60]), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (Plaintext_s2[60]), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (Plaintext_s0[61]), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (Plaintext_s1[61]), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (Plaintext_s2[61]), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (Ciphertext_s0[1]), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (Ciphertext_s1[1]), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (Ciphertext_s2[1]), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (SubCellInst_SboxInst_0_Q6), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_1749), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (SubCellInst_SboxInst_0_L2), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_1750), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_1751), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (Ciphertext_s0[5]), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (Ciphertext_s1[5]), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (Ciphertext_s2[5]), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (SubCellInst_SboxInst_1_Q6), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_1760), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_1761), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (SubCellInst_SboxInst_1_L2), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_1762), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (new_AGEMA_signal_1763), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (Ciphertext_s0[9]), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (Ciphertext_s1[9]), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (Ciphertext_s2[9]), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (SubCellInst_SboxInst_2_Q6), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (SubCellInst_SboxInst_2_L2), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_1774), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_1775), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (Ciphertext_s0[13]), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (Ciphertext_s1[13]), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (Ciphertext_s2[13]), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (SubCellInst_SboxInst_3_Q6), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_1785), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (SubCellInst_SboxInst_3_L2), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_1786), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (new_AGEMA_signal_1787), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (Ciphertext_s0[17]), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (Ciphertext_s1[17]), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (Ciphertext_s2[17]), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (SubCellInst_SboxInst_4_Q6), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_1797), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (SubCellInst_SboxInst_4_L2), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_1798), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_1799), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (Ciphertext_s0[21]), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (Ciphertext_s1[21]), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (Ciphertext_s2[21]), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (SubCellInst_SboxInst_5_Q6), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_1808), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_1809), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (SubCellInst_SboxInst_5_L2), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_1810), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (new_AGEMA_signal_1811), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (Ciphertext_s0[25]), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (Ciphertext_s1[25]), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (Ciphertext_s2[25]), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (SubCellInst_SboxInst_6_Q6), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_1821), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (SubCellInst_SboxInst_6_L2), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_1822), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_1823), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (Ciphertext_s0[29]), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (Ciphertext_s1[29]), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (Ciphertext_s2[29]), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (SubCellInst_SboxInst_7_Q6), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_1833), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (SubCellInst_SboxInst_7_L2), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (new_AGEMA_signal_1835), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (Ciphertext_s0[33]), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (Ciphertext_s1[33]), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (Ciphertext_s2[33]), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (SubCellInst_SboxInst_8_Q6), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_1845), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (SubCellInst_SboxInst_8_L2), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_1847), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (Ciphertext_s0[37]), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (Ciphertext_s1[37]), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (Ciphertext_s2[37]), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (SubCellInst_SboxInst_9_Q6), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_1857), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (SubCellInst_SboxInst_9_L2), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (new_AGEMA_signal_1859), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (Ciphertext_s0[41]), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (Ciphertext_s1[41]), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (Ciphertext_s2[41]), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (SubCellInst_SboxInst_10_Q6), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (new_AGEMA_signal_1868), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_1869), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (SubCellInst_SboxInst_10_L2), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_1870), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_1871), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (Ciphertext_s0[45]), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (Ciphertext_s1[45]), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (Ciphertext_s2[45]), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (SubCellInst_SboxInst_11_Q6), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_1881), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (SubCellInst_SboxInst_11_L2), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (new_AGEMA_signal_1883), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (Ciphertext_s0[49]), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (Ciphertext_s1[49]), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (Ciphertext_s2[49]), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (SubCellInst_SboxInst_12_Q6), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_1893), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (SubCellInst_SboxInst_12_L2), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_1894), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_1895), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (Ciphertext_s0[53]), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (Ciphertext_s1[53]), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (Ciphertext_s2[53]), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (SubCellInst_SboxInst_13_Q6), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_1905), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (SubCellInst_SboxInst_13_L2), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_1907), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (Ciphertext_s0[57]), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (Ciphertext_s1[57]), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (Ciphertext_s2[57]), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (SubCellInst_SboxInst_14_Q6), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_1917), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (SubCellInst_SboxInst_14_L2), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_1919), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (Ciphertext_s0[61]), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (Ciphertext_s1[61]), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (Ciphertext_s2[61]), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (SubCellInst_SboxInst_15_Q6), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_1929), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (SubCellInst_SboxInst_15_L2), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_1930), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_1931), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (FSMUpdate[1]), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (FSM[1]), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (FSM[4]), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (FSM[5]), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (TweakeyGeneration_key_Feedback[0]), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_1356), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_1357), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (TweakeyGeneration_key_Feedback[1]), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_1362), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_1363), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (TweakeyGeneration_key_Feedback[4]), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_1380), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_1381), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (TweakeyGeneration_key_Feedback[5]), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_1386), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_1387), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (TweakeyGeneration_key_Feedback[8]), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_1404), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_1405), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (TweakeyGeneration_key_Feedback[9]), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_1410), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_1411), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (TweakeyGeneration_key_Feedback[12]), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_1428), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_1429), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (TweakeyGeneration_key_Feedback[13]), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_1434), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_1435), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (TweakeyGeneration_key_Feedback[16]), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_1452), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_1453), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (TweakeyGeneration_key_Feedback[17]), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_1459), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (TweakeyGeneration_key_Feedback[20]), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_1477), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (TweakeyGeneration_key_Feedback[21]), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_1482), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_1483), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (TweakeyGeneration_key_Feedback[24]), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_1500), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_1501), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (TweakeyGeneration_key_Feedback[25]), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_1507), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (TweakeyGeneration_key_Feedback[28]), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_1524), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_1525), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (TweakeyGeneration_key_Feedback[29]), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_1530), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_1531), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (TweakeyGeneration_StateRegInput[63]), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_1738), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_1739), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (TweakeyGeneration_StateRegInput[62]), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_1732), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_1733), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (TweakeyGeneration_StateRegInput[61]), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_1726), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_1727), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (TweakeyGeneration_StateRegInput[60]), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_1720), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_1721), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (TweakeyGeneration_StateRegInput[59]), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_1715), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (TweakeyGeneration_StateRegInput[58]), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (TweakeyGeneration_StateRegInput[57]), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_1702), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_1703), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (TweakeyGeneration_StateRegInput[56]), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_1696), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_1697), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (TweakeyGeneration_StateRegInput[55]), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_1690), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_1691), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (TweakeyGeneration_StateRegInput[54]), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_1684), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_1685), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (TweakeyGeneration_StateRegInput[53]), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_1678), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_1679), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (TweakeyGeneration_StateRegInput[52]), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_1672), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_1673), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (TweakeyGeneration_StateRegInput[51]), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_1666), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_1667), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (TweakeyGeneration_StateRegInput[50]), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_1660), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_1661), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (TweakeyGeneration_StateRegInput[49]), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_1654), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_1655), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (TweakeyGeneration_StateRegInput[48]), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_1648), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_1649), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (TweakeyGeneration_StateRegInput[47]), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_1642), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_1643), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (TweakeyGeneration_StateRegInput[46]), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_1636), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_1637), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (TweakeyGeneration_StateRegInput[45]), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_1630), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_1631), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (TweakeyGeneration_StateRegInput[44]), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_1624), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_1625), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (TweakeyGeneration_StateRegInput[43]), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_1618), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_1619), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (TweakeyGeneration_StateRegInput[42]), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_1612), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_1613), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (TweakeyGeneration_StateRegInput[41]), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_1606), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_1607), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (TweakeyGeneration_StateRegInput[40]), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_1600), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_1601), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (TweakeyGeneration_StateRegInput[39]), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_1594), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_1595), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (TweakeyGeneration_StateRegInput[38]), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_1588), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_1589), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (TweakeyGeneration_StateRegInput[37]), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_1582), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_1583), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (TweakeyGeneration_StateRegInput[36]), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_1576), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_1577), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (TweakeyGeneration_StateRegInput[35]), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_1570), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_1571), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (TweakeyGeneration_StateRegInput[34]), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_1564), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_1565), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (TweakeyGeneration_StateRegInput[33]), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_1558), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_1559), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (TweakeyGeneration_StateRegInput[32]), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_1552), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_1553), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (TweakeyGeneration_StateRegInput[31]), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_1546), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_1547), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (TweakeyGeneration_StateRegInput[30]), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_1540), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_1541), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (TweakeyGeneration_StateRegInput[29]), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_1534), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_1535), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (TweakeyGeneration_StateRegInput[28]), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_1528), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_1529), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (TweakeyGeneration_StateRegInput[27]), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_1522), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_1523), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (TweakeyGeneration_StateRegInput[26]), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_1516), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_1517), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (TweakeyGeneration_StateRegInput[25]), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_1510), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_1511), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (TweakeyGeneration_StateRegInput[24]), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_1504), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_1505), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (TweakeyGeneration_StateRegInput[23]), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_1498), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_1499), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (TweakeyGeneration_StateRegInput[22]), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_1492), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_1493), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (TweakeyGeneration_StateRegInput[21]), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_1486), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_1487), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (TweakeyGeneration_StateRegInput[20]), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_1480), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_1481), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (TweakeyGeneration_StateRegInput[19]), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_1474), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_1475), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (TweakeyGeneration_StateRegInput[18]), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_1468), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_1469), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (TweakeyGeneration_StateRegInput[17]), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_1462), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_1463), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (TweakeyGeneration_StateRegInput[16]), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_1456), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_1457), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (TweakeyGeneration_StateRegInput[15]), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_1450), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_1451), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (TweakeyGeneration_StateRegInput[14]), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_1444), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (TweakeyGeneration_StateRegInput[13]), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_1438), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_1439), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (TweakeyGeneration_StateRegInput[12]), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_1432), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (TweakeyGeneration_StateRegInput[11]), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_1426), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_1427), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (TweakeyGeneration_StateRegInput[10]), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_1420), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_1421), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (TweakeyGeneration_StateRegInput[9]), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_1414), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_1415), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (TweakeyGeneration_StateRegInput[8]), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_1408), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (TweakeyGeneration_StateRegInput[7]), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_1402), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_1403), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (TweakeyGeneration_StateRegInput[6]), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_1396), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (TweakeyGeneration_StateRegInput[5]), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_1390), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_1391), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (TweakeyGeneration_StateRegInput[4]), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_1384), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_1385), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (TweakeyGeneration_StateRegInput[3]), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_1378), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_1379), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (TweakeyGeneration_StateRegInput[2]), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_1372), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (TweakeyGeneration_StateRegInput[1]), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_1366), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_1367), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (TweakeyGeneration_StateRegInput[0]), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_1360), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (FSMSelected[5]), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (FSMSelected[4]), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (FSMSelected[3]), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (FSMSelected[2]), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (FSMSelected[1]), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (FSMSelected[0]), .Q (new_AGEMA_signal_4884) ) ;

    /* cells in depth 2 */
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_0_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, MCOutput[0]}), .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3813, new_AGEMA_signal_3811}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_1_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, MCOutput[1]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3819, new_AGEMA_signal_3817}), .c ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_4_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCOutput[4]}), .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3825, new_AGEMA_signal_3823}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_5_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCOutput[5]}), .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3831, new_AGEMA_signal_3829}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_8_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, MCOutput[8]}), .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3837, new_AGEMA_signal_3835}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_9_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, MCOutput[9]}), .a ({new_AGEMA_signal_3845, new_AGEMA_signal_3843, new_AGEMA_signal_3841}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_12_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, MCOutput[12]}), .a ({new_AGEMA_signal_3851, new_AGEMA_signal_3849, new_AGEMA_signal_3847}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_13_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, MCOutput[13]}), .a ({new_AGEMA_signal_3857, new_AGEMA_signal_3855, new_AGEMA_signal_3853}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_16_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, MCOutput[16]}), .a ({new_AGEMA_signal_3863, new_AGEMA_signal_3861, new_AGEMA_signal_3859}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_17_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCOutput[17]}), .a ({new_AGEMA_signal_3869, new_AGEMA_signal_3867, new_AGEMA_signal_3865}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_20_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, MCOutput[20]}), .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3873, new_AGEMA_signal_3871}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_21_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, MCOutput[21]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3879, new_AGEMA_signal_3877}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_24_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, MCOutput[24]}), .a ({new_AGEMA_signal_3887, new_AGEMA_signal_3885, new_AGEMA_signal_3883}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_25_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, MCOutput[25]}), .a ({new_AGEMA_signal_3893, new_AGEMA_signal_3891, new_AGEMA_signal_3889}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_28_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, MCOutput[28]}), .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3897, new_AGEMA_signal_3895}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_29_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, MCOutput[29]}), .a ({new_AGEMA_signal_3905, new_AGEMA_signal_3903, new_AGEMA_signal_3901}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_32_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .a ({new_AGEMA_signal_3911, new_AGEMA_signal_3909, new_AGEMA_signal_3907}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_33_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .a ({new_AGEMA_signal_3917, new_AGEMA_signal_3915, new_AGEMA_signal_3913}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_36_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .a ({new_AGEMA_signal_3923, new_AGEMA_signal_3921, new_AGEMA_signal_3919}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_37_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .a ({new_AGEMA_signal_3929, new_AGEMA_signal_3927, new_AGEMA_signal_3925}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_40_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .a ({new_AGEMA_signal_3935, new_AGEMA_signal_3933, new_AGEMA_signal_3931}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_41_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .a ({new_AGEMA_signal_3941, new_AGEMA_signal_3939, new_AGEMA_signal_3937}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_44_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .a ({new_AGEMA_signal_3947, new_AGEMA_signal_3945, new_AGEMA_signal_3943}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_45_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .a ({new_AGEMA_signal_3953, new_AGEMA_signal_3951, new_AGEMA_signal_3949}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_48_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[48]}), .a ({new_AGEMA_signal_3959, new_AGEMA_signal_3957, new_AGEMA_signal_3955}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_49_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, MCOutput[49]}), .a ({new_AGEMA_signal_3965, new_AGEMA_signal_3963, new_AGEMA_signal_3961}), .c ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_52_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, MCOutput[52]}), .a ({new_AGEMA_signal_3971, new_AGEMA_signal_3969, new_AGEMA_signal_3967}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_53_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCOutput[53]}), .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3975, new_AGEMA_signal_3973}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_56_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, MCOutput[56]}), .a ({new_AGEMA_signal_3983, new_AGEMA_signal_3981, new_AGEMA_signal_3979}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_57_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCOutput[57]}), .a ({new_AGEMA_signal_3989, new_AGEMA_signal_3987, new_AGEMA_signal_3985}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_60_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCOutput[60]}), .a ({new_AGEMA_signal_3995, new_AGEMA_signal_3993, new_AGEMA_signal_3991}), .c ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) PlaintextMUX_MUXInst_61_U1 ( .s (new_AGEMA_signal_3809), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCOutput[61]}), .a ({new_AGEMA_signal_4001, new_AGEMA_signal_3999, new_AGEMA_signal_3997}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, StateRegInput[61]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_AND2_U1 ( .a ({new_AGEMA_signal_4004, new_AGEMA_signal_4003, new_AGEMA_signal_4002}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, SubCellInst_SboxInst_0_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR4_U1 ( .a ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, SubCellInst_SboxInst_0_T1}), .b ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, new_AGEMA_signal_4005}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_AND4_U1 ( .a ({new_AGEMA_signal_4010, new_AGEMA_signal_4009, new_AGEMA_signal_4008}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_0_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR9_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_4016, new_AGEMA_signal_4014, new_AGEMA_signal_4012}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, SubCellInst_SboxInst_0_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR10_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_0_T3}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, ShiftRowsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .a ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, new_AGEMA_signal_4017}), .b ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, SubCellInst_SboxInst_0_YY_3}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, ShiftRowsOutput[5]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_AND2_U1 ( .a ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_1_Q2}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_1_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR4_U1 ( .a ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_1_T1}), .b ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_AND4_U1 ( .a ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, SubCellInst_SboxInst_1_Q7}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, SubCellInst_SboxInst_1_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR9_U1 ( .a ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_4034, new_AGEMA_signal_4032, new_AGEMA_signal_4030}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR10_U1 ( .a ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, SubCellInst_SboxInst_1_T3}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .a ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, new_AGEMA_signal_4035}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, ShiftRowsOutput[9]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_AND2_U1 ( .a ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, SubCellInst_SboxInst_2_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR4_U1 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, SubCellInst_SboxInst_2_T1}), .b ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, new_AGEMA_signal_4041}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_AND4_U1 ( .a ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, new_AGEMA_signal_4044}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, SubCellInst_SboxInst_2_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR9_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_4052, new_AGEMA_signal_4050, new_AGEMA_signal_4048}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR10_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, SubCellInst_SboxInst_2_T3}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, ShiftRowsOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .a ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, new_AGEMA_signal_4053}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[13]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_AND2_U1 ( .a ({new_AGEMA_signal_4058, new_AGEMA_signal_4057, new_AGEMA_signal_4056}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_3_Q2}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, SubCellInst_SboxInst_3_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR4_U1 ( .a ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, SubCellInst_SboxInst_3_T1}), .b ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, new_AGEMA_signal_4059}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_AND4_U1 ( .a ({new_AGEMA_signal_4064, new_AGEMA_signal_4063, new_AGEMA_signal_4062}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_3_Q7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_3_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR9_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_4070, new_AGEMA_signal_4068, new_AGEMA_signal_4066}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR10_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_3_T3}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, ShiftRowsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .a ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, new_AGEMA_signal_4071}), .b ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, ShiftRowsOutput[1]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_AND2_U1 ( .a ({new_AGEMA_signal_4076, new_AGEMA_signal_4075, new_AGEMA_signal_4074}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, SubCellInst_SboxInst_4_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR4_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, SubCellInst_SboxInst_4_T1}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, new_AGEMA_signal_4077}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_AND4_U1 ( .a ({new_AGEMA_signal_4082, new_AGEMA_signal_4081, new_AGEMA_signal_4080}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, SubCellInst_SboxInst_4_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR9_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_4088, new_AGEMA_signal_4086, new_AGEMA_signal_4084}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR10_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, SubCellInst_SboxInst_4_T3}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .a ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, new_AGEMA_signal_4089}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_AND2_U1 ( .a ({new_AGEMA_signal_4094, new_AGEMA_signal_4093, new_AGEMA_signal_4092}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, SubCellInst_SboxInst_5_Q2}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, SubCellInst_SboxInst_5_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR4_U1 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, SubCellInst_SboxInst_5_T1}), .b ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, new_AGEMA_signal_4095}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_AND4_U1 ( .a ({new_AGEMA_signal_4100, new_AGEMA_signal_4099, new_AGEMA_signal_4098}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_5_Q7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, SubCellInst_SboxInst_5_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR9_U1 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_4106, new_AGEMA_signal_4104, new_AGEMA_signal_4102}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR10_U1 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, SubCellInst_SboxInst_5_T3}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, new_AGEMA_signal_4107}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_AND2_U1 ( .a ({new_AGEMA_signal_4112, new_AGEMA_signal_4111, new_AGEMA_signal_4110}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, SubCellInst_SboxInst_6_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR4_U1 ( .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, SubCellInst_SboxInst_6_T1}), .b ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, new_AGEMA_signal_4113}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_AND4_U1 ( .a ({new_AGEMA_signal_4118, new_AGEMA_signal_4117, new_AGEMA_signal_4116}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, SubCellInst_SboxInst_6_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR9_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_4124, new_AGEMA_signal_4122, new_AGEMA_signal_4120}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR10_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, SubCellInst_SboxInst_6_T3}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, new_AGEMA_signal_4125}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_AND2_U1 ( .a ({new_AGEMA_signal_4130, new_AGEMA_signal_4129, new_AGEMA_signal_4128}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, SubCellInst_SboxInst_7_Q2}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_7_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR4_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_7_T1}), .b ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, new_AGEMA_signal_4131}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_AND4_U1 ( .a ({new_AGEMA_signal_4136, new_AGEMA_signal_4135, new_AGEMA_signal_4134}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, SubCellInst_SboxInst_7_Q7}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, SubCellInst_SboxInst_7_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR9_U1 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_4142, new_AGEMA_signal_4140, new_AGEMA_signal_4138}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR10_U1 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, SubCellInst_SboxInst_7_T3}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .a ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, new_AGEMA_signal_4143}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellOutput[29]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_AND2_U1 ( .a ({new_AGEMA_signal_4148, new_AGEMA_signal_4147, new_AGEMA_signal_4146}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR4_U1 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1}), .b ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, new_AGEMA_signal_4149}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_AND4_U1 ( .a ({new_AGEMA_signal_4154, new_AGEMA_signal_4153, new_AGEMA_signal_4152}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR9_U1 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_4160, new_AGEMA_signal_4158, new_AGEMA_signal_4156}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, SubCellInst_SboxInst_8_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR10_U1 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, AddRoundConstantOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, new_AGEMA_signal_4161}), .b ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, SubCellInst_SboxInst_8_YY_3}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, AddRoundConstantOutput[33]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_AND2_U1 ( .a ({new_AGEMA_signal_4166, new_AGEMA_signal_4165, new_AGEMA_signal_4164}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, SubCellInst_SboxInst_9_Q2}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, SubCellInst_SboxInst_9_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR4_U1 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, SubCellInst_SboxInst_9_T1}), .b ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, new_AGEMA_signal_4167}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_AND4_U1 ( .a ({new_AGEMA_signal_4172, new_AGEMA_signal_4171, new_AGEMA_signal_4170}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, SubCellInst_SboxInst_9_Q7}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_9_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR9_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_4178, new_AGEMA_signal_4176, new_AGEMA_signal_4174}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR10_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_9_T3}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, AddRoundConstantOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .a ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, new_AGEMA_signal_4179}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, AddRoundConstantOutput[37]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_AND2_U1 ( .a ({new_AGEMA_signal_4184, new_AGEMA_signal_4183, new_AGEMA_signal_4182}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_10_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR4_U1 ( .a ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_10_T1}), .b ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, new_AGEMA_signal_4185}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_AND4_U1 ( .a ({new_AGEMA_signal_4190, new_AGEMA_signal_4189, new_AGEMA_signal_4188}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, SubCellInst_SboxInst_10_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR9_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_4196, new_AGEMA_signal_4194, new_AGEMA_signal_4192}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR10_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, SubCellInst_SboxInst_10_T3}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, AddRoundConstantOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .a ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, new_AGEMA_signal_4197}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, AddRoundConstantOutput[41]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_AND2_U1 ( .a ({new_AGEMA_signal_4202, new_AGEMA_signal_4201, new_AGEMA_signal_4200}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, SubCellInst_SboxInst_11_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR4_U1 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, SubCellInst_SboxInst_11_T1}), .b ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, new_AGEMA_signal_4203}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_AND4_U1 ( .a ({new_AGEMA_signal_4208, new_AGEMA_signal_4207, new_AGEMA_signal_4206}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, SubCellInst_SboxInst_11_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR9_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_4214, new_AGEMA_signal_4212, new_AGEMA_signal_4210}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR10_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, SubCellInst_SboxInst_11_T3}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .a ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, new_AGEMA_signal_4215}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, SubCellOutput[45]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_AND2_U1 ( .a ({new_AGEMA_signal_4220, new_AGEMA_signal_4219, new_AGEMA_signal_4218}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_12_Q2}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, SubCellInst_SboxInst_12_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR4_U1 ( .a ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, SubCellInst_SboxInst_12_T1}), .b ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, new_AGEMA_signal_4221}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_AND4_U1 ( .a ({new_AGEMA_signal_4226, new_AGEMA_signal_4225, new_AGEMA_signal_4224}), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, SubCellInst_SboxInst_12_Q7}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR9_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_4232, new_AGEMA_signal_4230, new_AGEMA_signal_4228}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR10_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_T3}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, AddRoundConstantOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .a ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, new_AGEMA_signal_4233}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, AddRoundConstantOutput[49]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_AND2_U1 ( .a ({new_AGEMA_signal_4238, new_AGEMA_signal_4237, new_AGEMA_signal_4236}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, SubCellInst_SboxInst_13_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR4_U1 ( .a ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, SubCellInst_SboxInst_13_T1}), .b ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, new_AGEMA_signal_4239}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_AND4_U1 ( .a ({new_AGEMA_signal_4244, new_AGEMA_signal_4243, new_AGEMA_signal_4242}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, SubCellInst_SboxInst_13_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR9_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_4250, new_AGEMA_signal_4248, new_AGEMA_signal_4246}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR10_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, SubCellInst_SboxInst_13_T3}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, AddRoundConstantOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, new_AGEMA_signal_4251}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, AddRoundConstantOutput[53]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_AND2_U1 ( .a ({new_AGEMA_signal_4256, new_AGEMA_signal_4255, new_AGEMA_signal_4254}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, SubCellInst_SboxInst_14_Q2}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, SubCellInst_SboxInst_14_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR4_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, SubCellInst_SboxInst_14_T1}), .b ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, new_AGEMA_signal_4257}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_AND4_U1 ( .a ({new_AGEMA_signal_4262, new_AGEMA_signal_4261, new_AGEMA_signal_4260}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_14_Q7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, SubCellInst_SboxInst_14_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR9_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_4268, new_AGEMA_signal_4266, new_AGEMA_signal_4264}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR10_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, SubCellInst_SboxInst_14_T3}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, AddRoundConstantOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, new_AGEMA_signal_4269}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, AddRoundConstantOutput[57]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_AND2_U1 ( .a ({new_AGEMA_signal_4274, new_AGEMA_signal_4273, new_AGEMA_signal_4272}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, SubCellInst_SboxInst_15_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR4_U1 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, SubCellInst_SboxInst_15_T1}), .b ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, new_AGEMA_signal_4275}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_AND4_U1 ( .a ({new_AGEMA_signal_4280, new_AGEMA_signal_4279, new_AGEMA_signal_4278}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, SubCellInst_SboxInst_15_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR9_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_4286, new_AGEMA_signal_4284, new_AGEMA_signal_4282}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR10_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, SubCellInst_SboxInst_15_T3}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, SubCellOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .a ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, new_AGEMA_signal_4287}), .b ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, SubCellOutput[61]}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) AddConstXOR_U2 ( .a ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellOutput[29]}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, AddConstXOR_AddConstXOR_XORInst_0_0_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_4291}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, AddRoundConstantOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, SubCellOutput[60]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, AddConstXOR_AddConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_4293}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, AddRoundConstantOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, SubCellOutput[61]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, AddConstXOR_AddConstXOR_XORInst_1_0_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_4295}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, AddRoundConstantOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellOutput[44]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, AddConstXOR_AddConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1}), .b ({1'b0, 1'b0, new_AGEMA_signal_4297}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, AddRoundConstantOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, SubCellOutput[45]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1}), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4301, new_AGEMA_signal_4299}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, ShiftRowsOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, AddRoundConstantOutput[32]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1}), .b ({new_AGEMA_signal_4309, new_AGEMA_signal_4307, new_AGEMA_signal_4305}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, ShiftRowsOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, AddRoundConstantOutput[33]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1}), .b ({new_AGEMA_signal_4315, new_AGEMA_signal_4313, new_AGEMA_signal_4311}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, ShiftRowsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, AddRoundConstantOutput[36]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1}), .b ({new_AGEMA_signal_4321, new_AGEMA_signal_4319, new_AGEMA_signal_4317}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, AddRoundConstantOutput[37]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1}), .b ({new_AGEMA_signal_4327, new_AGEMA_signal_4325, new_AGEMA_signal_4323}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, AddRoundConstantOutput[40]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1}), .b ({new_AGEMA_signal_4333, new_AGEMA_signal_4331, new_AGEMA_signal_4329}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, AddRoundConstantOutput[41]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1}), .b ({new_AGEMA_signal_4339, new_AGEMA_signal_4337, new_AGEMA_signal_4335}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, AddRoundConstantOutput[44]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1}), .b ({new_AGEMA_signal_4345, new_AGEMA_signal_4343, new_AGEMA_signal_4341}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, ShiftRowsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, AddRoundConstantOutput[45]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, AddRoundTweakeyXOR_XORInst_4_0_n1}), .b ({new_AGEMA_signal_4351, new_AGEMA_signal_4349, new_AGEMA_signal_4347}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, AddRoundConstantOutput[48]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, AddRoundTweakeyXOR_XORInst_4_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1}), .b ({new_AGEMA_signal_4357, new_AGEMA_signal_4355, new_AGEMA_signal_4353}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, AddRoundConstantOutput[49]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, AddRoundTweakeyXOR_XORInst_5_0_n1}), .b ({new_AGEMA_signal_4363, new_AGEMA_signal_4361, new_AGEMA_signal_4359}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, AddRoundConstantOutput[52]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, AddRoundTweakeyXOR_XORInst_5_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1}), .b ({new_AGEMA_signal_4369, new_AGEMA_signal_4367, new_AGEMA_signal_4365}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, AddRoundConstantOutput[53]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, AddRoundTweakeyXOR_XORInst_6_0_n1}), .b ({new_AGEMA_signal_4375, new_AGEMA_signal_4373, new_AGEMA_signal_4371}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, AddRoundConstantOutput[56]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, AddRoundTweakeyXOR_XORInst_6_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1}), .b ({new_AGEMA_signal_4381, new_AGEMA_signal_4379, new_AGEMA_signal_4377}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, AddRoundConstantOutput[57]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, AddRoundTweakeyXOR_XORInst_7_0_n1}), .b ({new_AGEMA_signal_4387, new_AGEMA_signal_4385, new_AGEMA_signal_4383}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, AddRoundConstantOutput[60]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, AddRoundTweakeyXOR_XORInst_7_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1}), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4391, new_AGEMA_signal_4389}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, AddRoundConstantOutput[61]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, MCInst_MCR0_XORInst_0_0_n1}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, MCInst_MCR0_XORInst_0_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, MCInst_MCR0_XORInst_0_1_n1}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, MCOutput[49]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, MCInst_MCR0_XORInst_0_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, MCInst_MCR0_XORInst_1_0_n1}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, MCOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, MCInst_MCR0_XORInst_1_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, MCInst_MCR0_XORInst_1_1_n1}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCOutput[53]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, MCInst_MCR0_XORInst_1_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U3 ( .a ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2}), .b ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, MCInst_MCR0_XORInst_2_0_n1}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, MCOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, MCInst_MCR0_XORInst_2_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U3 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, MCInst_MCR0_XORInst_2_1_n1}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, MCInst_MCR0_XORInst_2_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U3 ( .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, MCInst_MCR0_XORInst_3_0_n1}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, MCInst_MCR0_XORInst_3_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U3 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, MCInst_MCR0_XORInst_3_1_n1}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, MCInst_MCR0_XORInst_3_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR0_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, MCInst_MCR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, MCOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, MCInst_MCR2_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCOutput[17]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCInst_MCR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, MCOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCInst_MCR2_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, MCOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, MCInst_MCR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, MCOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, MCInst_MCR2_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, MCOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCInst_MCR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, MCOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCInst_MCR2_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, MCOutput[29]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, MCInst_MCR3_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, MCOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, MCInst_MCR3_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, MCOutput[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, MCInst_MCR3_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, MCInst_MCR3_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCInst_MCR3_XORInst_2_0_n1}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, MCOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCInst_MCR3_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, MCOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, MCInst_MCR3_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, MCOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .c ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, MCInst_MCR3_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, MCOutput[13]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MCInst_MCR3_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1}) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_3470), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_3810), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_3818), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_3820), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_3822), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_3824), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_3826), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_3834), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_3842), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_3850), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_3858), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_3866), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_3874), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_3882), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_3906), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_3930), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (SubCellInst_SboxInst_0_T2), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_1934), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_1935), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (SubCellInst_SboxInst_0_YY_1_), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_2162), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_2163), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (SubCellInst_SboxInst_1_T2), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_1941), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (SubCellInst_SboxInst_1_YY_1_), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_2170), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_2171), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (SubCellInst_SboxInst_2_T2), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_1947), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (SubCellInst_SboxInst_2_YY_1_), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_2178), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_2179), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (SubCellInst_SboxInst_3_T2), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_1952), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_1953), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (SubCellInst_SboxInst_3_YY_1_), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_2186), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_2187), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (SubCellInst_SboxInst_4_T2), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_1958), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_1959), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (SubCellInst_SboxInst_4_YY_1_), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_2194), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_2195), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (SubCellInst_SboxInst_5_T2), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_1964), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_1965), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_4101), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (SubCellInst_SboxInst_5_YY_1_), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_2202), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_2203), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (SubCellInst_SboxInst_6_T2), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_1970), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_1971), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (SubCellInst_SboxInst_6_YY_1_), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_2210), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_2211), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (SubCellInst_SboxInst_7_T2), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_1977), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_4137), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (SubCellInst_SboxInst_7_YY_1_), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_2218), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_2219), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (SubCellInst_SboxInst_8_T2), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_1983), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_4157), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (SubCellInst_SboxInst_8_YY_1_), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_2226), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_2227), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (SubCellInst_SboxInst_9_T2), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (SubCellInst_SboxInst_9_YY_1_), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_2234), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_2235), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (SubCellInst_SboxInst_10_T2), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_1995), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_4193), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (SubCellInst_SboxInst_10_YY_1_), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_2242), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_2243), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (SubCellInst_SboxInst_11_T2), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_2001), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_4211), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (SubCellInst_SboxInst_11_YY_1_), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_2250), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_2251), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (SubCellInst_SboxInst_12_T2), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_2006), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_2007), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_4227), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (SubCellInst_SboxInst_12_YY_1_), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_2258), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_2259), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (SubCellInst_SboxInst_13_T2), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_2012), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_2013), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_4245), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_4247), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (SubCellInst_SboxInst_13_YY_1_), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_2266), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_2267), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (SubCellInst_SboxInst_14_T2), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_2019), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_4263), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (SubCellInst_SboxInst_14_YY_1_), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_2274), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_2275), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (SubCellInst_SboxInst_15_T2), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_2025), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_4281), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_4283), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (SubCellInst_SboxInst_15_YY_1_), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_2282), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_2283), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_4290), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_4296), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_4302), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_4314), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_4338), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_4362), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_4374), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_4378), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (new_AGEMA_signal_4380), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_4386), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_4392), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (StateRegInput[63]), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (StateRegInput[62]), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_2956), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_2957), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (StateRegInput[59]), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_2848), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_2849), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (StateRegInput[58]), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_2728), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (StateRegInput[55]), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_2844), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (StateRegInput[54]), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_2724), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_2725), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (StateRegInput[51]), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_2840), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_2841), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (StateRegInput[50]), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_2721), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (StateRegInput[47]), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_2836), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (StateRegInput[46]), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_2716), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (StateRegInput[43]), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (StateRegInput[42]), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_2486), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_2487), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (StateRegInput[39]), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_2589), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (StateRegInput[38]), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_2482), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_2483), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (StateRegInput[35]), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (StateRegInput[34]), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_2479), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (StateRegInput[31]), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_2820), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (StateRegInput[30]), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_2700), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (StateRegInput[27]), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_3019), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (StateRegInput[26]), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_2932), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_2933), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (StateRegInput[23]), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_2816), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_2817), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (StateRegInput[22]), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_2697), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (StateRegInput[19]), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (StateRegInput[18]), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (StateRegInput[15]), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (StateRegInput[14]), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_2920), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_2921), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (StateRegInput[11]), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_2808), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (StateRegInput[10]), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_2688), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (StateRegInput[7]), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_2804), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (StateRegInput[6]), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (StateRegInput[3]), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_2800), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (StateRegInput[2]), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_2680), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_4494), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_4498), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_4500), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_4502), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_4506), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_4512), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_4518), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_4522), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (new_AGEMA_signal_4524), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_4526), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_4530), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_4534), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_4536), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_4538), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_4542), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_4548), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_4554), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (new_AGEMA_signal_4560), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_4566), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_4578), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_4584), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_4596), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_4602), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_4620), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_4650), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_4656), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_4668), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_4674), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_4692), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_4704), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4396, new_AGEMA_signal_4395, new_AGEMA_signal_4394}), .Q ({Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, new_AGEMA_signal_4397}), .Q ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, StateRegInput[61]}), .Q ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, StateRegInput[60]}), .Q ({Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4402, new_AGEMA_signal_4401, new_AGEMA_signal_4400}), .Q ({Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, new_AGEMA_signal_4403}), .Q ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, StateRegInput[57]}), .Q ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, StateRegInput[56]}), .Q ({Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4408, new_AGEMA_signal_4407, new_AGEMA_signal_4406}), .Q ({Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, new_AGEMA_signal_4409}), .Q ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, StateRegInput[53]}), .Q ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, StateRegInput[52]}), .Q ({Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4414, new_AGEMA_signal_4413, new_AGEMA_signal_4412}), .Q ({Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, new_AGEMA_signal_4415}), .Q ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, StateRegInput[49]}), .Q ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, StateRegInput[48]}), .Q ({Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, new_AGEMA_signal_4418}), .Q ({Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, new_AGEMA_signal_4421}), .Q ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, StateRegInput[45]}), .Q ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, StateRegInput[44]}), .Q ({Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, new_AGEMA_signal_4424}), .Q ({Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, new_AGEMA_signal_4427}), .Q ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, StateRegInput[41]}), .Q ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, StateRegInput[40]}), .Q ({Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, new_AGEMA_signal_4430}), .Q ({Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, new_AGEMA_signal_4433}), .Q ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, StateRegInput[37]}), .Q ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, StateRegInput[36]}), .Q ({Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, new_AGEMA_signal_4436}), .Q ({Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, new_AGEMA_signal_4439}), .Q ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, StateRegInput[33]}), .Q ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, StateRegInput[32]}), .Q ({Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, new_AGEMA_signal_4442}), .Q ({Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, new_AGEMA_signal_4445}), .Q ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, StateRegInput[29]}), .Q ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, StateRegInput[28]}), .Q ({Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, new_AGEMA_signal_4448}), .Q ({Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, new_AGEMA_signal_4451}), .Q ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, StateRegInput[25]}), .Q ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, StateRegInput[24]}), .Q ({Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4456, new_AGEMA_signal_4455, new_AGEMA_signal_4454}), .Q ({Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, new_AGEMA_signal_4457}), .Q ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, StateRegInput[21]}), .Q ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, StateRegInput[20]}), .Q ({Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4462, new_AGEMA_signal_4461, new_AGEMA_signal_4460}), .Q ({Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, new_AGEMA_signal_4463}), .Q ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, StateRegInput[17]}), .Q ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, StateRegInput[16]}), .Q ({Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4468, new_AGEMA_signal_4467, new_AGEMA_signal_4466}), .Q ({Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, new_AGEMA_signal_4469}), .Q ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, StateRegInput[13]}), .Q ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, StateRegInput[12]}), .Q ({Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4474, new_AGEMA_signal_4473, new_AGEMA_signal_4472}), .Q ({Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, new_AGEMA_signal_4475}), .Q ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, StateRegInput[9]}), .Q ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, StateRegInput[8]}), .Q ({Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4480, new_AGEMA_signal_4479, new_AGEMA_signal_4478}), .Q ({Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, new_AGEMA_signal_4481}), .Q ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, StateRegInput[5]}), .Q ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, StateRegInput[4]}), .Q ({Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4486, new_AGEMA_signal_4485, new_AGEMA_signal_4484}), .Q ({Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, new_AGEMA_signal_4487}), .Q ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, StateRegInput[1]}), .Q ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, StateRegInput[0]}), .Q ({Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4495, new_AGEMA_signal_4493, new_AGEMA_signal_4491}), .Q ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4501, new_AGEMA_signal_4499, new_AGEMA_signal_4497}), .Q ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, TweakeyGeneration_key_Feedback[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4507, new_AGEMA_signal_4505, new_AGEMA_signal_4503}), .Q ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_key_Feedback[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4513, new_AGEMA_signal_4511, new_AGEMA_signal_4509}), .Q ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4519, new_AGEMA_signal_4517, new_AGEMA_signal_4515}), .Q ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, TweakeyGeneration_key_Feedback[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4525, new_AGEMA_signal_4523, new_AGEMA_signal_4521}), .Q ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_key_Feedback[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4531, new_AGEMA_signal_4529, new_AGEMA_signal_4527}), .Q ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4537, new_AGEMA_signal_4535, new_AGEMA_signal_4533}), .Q ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, TweakeyGeneration_key_Feedback[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4543, new_AGEMA_signal_4541, new_AGEMA_signal_4539}), .Q ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_key_Feedback[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4549, new_AGEMA_signal_4547, new_AGEMA_signal_4545}), .Q ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4555, new_AGEMA_signal_4553, new_AGEMA_signal_4551}), .Q ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, TweakeyGeneration_key_Feedback[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4561, new_AGEMA_signal_4559, new_AGEMA_signal_4557}), .Q ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_key_Feedback[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4567, new_AGEMA_signal_4565, new_AGEMA_signal_4563}), .Q ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4573, new_AGEMA_signal_4571, new_AGEMA_signal_4569}), .Q ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, TweakeyGeneration_key_Feedback[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4579, new_AGEMA_signal_4577, new_AGEMA_signal_4575}), .Q ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_key_Feedback[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4585, new_AGEMA_signal_4583, new_AGEMA_signal_4581}), .Q ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4591, new_AGEMA_signal_4589, new_AGEMA_signal_4587}), .Q ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4597, new_AGEMA_signal_4595, new_AGEMA_signal_4593}), .Q ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4603, new_AGEMA_signal_4601, new_AGEMA_signal_4599}), .Q ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4609, new_AGEMA_signal_4607, new_AGEMA_signal_4605}), .Q ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4615, new_AGEMA_signal_4613, new_AGEMA_signal_4611}), .Q ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4621, new_AGEMA_signal_4619, new_AGEMA_signal_4617}), .Q ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4627, new_AGEMA_signal_4625, new_AGEMA_signal_4623}), .Q ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4633, new_AGEMA_signal_4631, new_AGEMA_signal_4629}), .Q ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4639, new_AGEMA_signal_4637, new_AGEMA_signal_4635}), .Q ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4645, new_AGEMA_signal_4643, new_AGEMA_signal_4641}), .Q ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4651, new_AGEMA_signal_4649, new_AGEMA_signal_4647}), .Q ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4657, new_AGEMA_signal_4655, new_AGEMA_signal_4653}), .Q ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4663, new_AGEMA_signal_4661, new_AGEMA_signal_4659}), .Q ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4669, new_AGEMA_signal_4667, new_AGEMA_signal_4665}), .Q ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4675, new_AGEMA_signal_4673, new_AGEMA_signal_4671}), .Q ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4681, new_AGEMA_signal_4679, new_AGEMA_signal_4677}), .Q ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4687, new_AGEMA_signal_4685, new_AGEMA_signal_4683}), .Q ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4693, new_AGEMA_signal_4691, new_AGEMA_signal_4689}), .Q ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, TweakeyGeneration_key_Feedback[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4699, new_AGEMA_signal_4697, new_AGEMA_signal_4695}), .Q ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_key_Feedback[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4705, new_AGEMA_signal_4703, new_AGEMA_signal_4701}), .Q ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4711, new_AGEMA_signal_4709, new_AGEMA_signal_4707}), .Q ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, TweakeyGeneration_key_Feedback[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4717, new_AGEMA_signal_4715, new_AGEMA_signal_4713}), .Q ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_key_Feedback[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4723, new_AGEMA_signal_4721, new_AGEMA_signal_4719}), .Q ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4729, new_AGEMA_signal_4727, new_AGEMA_signal_4725}), .Q ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, TweakeyGeneration_key_Feedback[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4735, new_AGEMA_signal_4733, new_AGEMA_signal_4731}), .Q ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_key_Feedback[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4741, new_AGEMA_signal_4739, new_AGEMA_signal_4737}), .Q ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4747, new_AGEMA_signal_4745, new_AGEMA_signal_4743}), .Q ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, TweakeyGeneration_key_Feedback[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4753, new_AGEMA_signal_4751, new_AGEMA_signal_4749}), .Q ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_key_Feedback[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4759, new_AGEMA_signal_4757, new_AGEMA_signal_4755}), .Q ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_key_Feedback[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4765, new_AGEMA_signal_4763, new_AGEMA_signal_4761}), .Q ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4771, new_AGEMA_signal_4769, new_AGEMA_signal_4767}), .Q ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, TweakeyGeneration_key_Feedback[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4777, new_AGEMA_signal_4775, new_AGEMA_signal_4773}), .Q ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_key_Feedback[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4783, new_AGEMA_signal_4781, new_AGEMA_signal_4779}), .Q ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, TweakeyGeneration_key_Feedback[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4789, new_AGEMA_signal_4787, new_AGEMA_signal_4785}), .Q ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_key_Feedback[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4795, new_AGEMA_signal_4793, new_AGEMA_signal_4791}), .Q ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4801, new_AGEMA_signal_4799, new_AGEMA_signal_4797}), .Q ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, TweakeyGeneration_key_Feedback[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4807, new_AGEMA_signal_4805, new_AGEMA_signal_4803}), .Q ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, TweakeyGeneration_key_Feedback[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4813, new_AGEMA_signal_4811, new_AGEMA_signal_4809}), .Q ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_key_Feedback[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4819, new_AGEMA_signal_4817, new_AGEMA_signal_4815}), .Q ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4825, new_AGEMA_signal_4823, new_AGEMA_signal_4821}), .Q ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, TweakeyGeneration_key_Feedback[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4831, new_AGEMA_signal_4829, new_AGEMA_signal_4827}), .Q ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4837, new_AGEMA_signal_4835, new_AGEMA_signal_4833}), .Q ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, TweakeyGeneration_key_Feedback[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4843, new_AGEMA_signal_4841, new_AGEMA_signal_4839}), .Q ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_key_Feedback[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4849, new_AGEMA_signal_4847, new_AGEMA_signal_4845}), .Q ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4855, new_AGEMA_signal_4853, new_AGEMA_signal_4851}), .Q ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_key_Feedback[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4861, new_AGEMA_signal_4859, new_AGEMA_signal_4857}), .Q ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4867, new_AGEMA_signal_4865, new_AGEMA_signal_4863}), .Q ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, TweakeyGeneration_key_Feedback[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4873, new_AGEMA_signal_4871, new_AGEMA_signal_4869}), .Q ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_key_Feedback[56]}) ) ;
    DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4875), .Q (FSM[5]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4877), .Q (FSM[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4879), .Q (FSMUpdate[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4881), .Q (FSMUpdate[3]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4883), .Q (FSM[1]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4885), .Q (FSMUpdate[1]), .QN () ) ;
endmodule
