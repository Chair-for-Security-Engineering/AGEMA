////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module SkinnyTop in file /AGEMA/Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module SkinnyTop_HPC3_ClockGating_d2 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Key_s2, Plaintext_s1, Plaintext_s2, Fresh, Ciphertext_s0, done, Ciphertext_s1, Ciphertext_s2, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Key_s2 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Plaintext_s2 ;
    input [383:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output [63:0] Ciphertext_s2 ;
    output Synch ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_YY_0_ ;
    wire SubCellInst_SboxInst_0_YY_1_ ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_0_XX_1_ ;
    wire SubCellInst_SboxInst_0_XX_2_ ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_YY_0_ ;
    wire SubCellInst_SboxInst_1_YY_1_ ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_1_XX_1_ ;
    wire SubCellInst_SboxInst_1_XX_2_ ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_YY_0_ ;
    wire SubCellInst_SboxInst_2_YY_1_ ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_2_XX_1_ ;
    wire SubCellInst_SboxInst_2_XX_2_ ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_YY_0_ ;
    wire SubCellInst_SboxInst_3_YY_1_ ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_3_XX_1_ ;
    wire SubCellInst_SboxInst_3_XX_2_ ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_YY_0_ ;
    wire SubCellInst_SboxInst_4_YY_1_ ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_4_XX_1_ ;
    wire SubCellInst_SboxInst_4_XX_2_ ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_YY_0_ ;
    wire SubCellInst_SboxInst_5_YY_1_ ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_5_XX_1_ ;
    wire SubCellInst_SboxInst_5_XX_2_ ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_YY_0_ ;
    wire SubCellInst_SboxInst_6_YY_1_ ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_6_XX_1_ ;
    wire SubCellInst_SboxInst_6_XX_2_ ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_YY_0_ ;
    wire SubCellInst_SboxInst_7_YY_1_ ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_7_XX_1_ ;
    wire SubCellInst_SboxInst_7_XX_2_ ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_YY_0_ ;
    wire SubCellInst_SboxInst_8_YY_1_ ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_8_XX_1_ ;
    wire SubCellInst_SboxInst_8_XX_2_ ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_YY_0_ ;
    wire SubCellInst_SboxInst_9_YY_1_ ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_9_XX_1_ ;
    wire SubCellInst_SboxInst_9_XX_2_ ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_YY_0_ ;
    wire SubCellInst_SboxInst_10_YY_1_ ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_10_XX_1_ ;
    wire SubCellInst_SboxInst_10_XX_2_ ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_YY_0_ ;
    wire SubCellInst_SboxInst_11_YY_1_ ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_11_XX_1_ ;
    wire SubCellInst_SboxInst_11_XX_2_ ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_YY_0_ ;
    wire SubCellInst_SboxInst_12_YY_1_ ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_12_XX_1_ ;
    wire SubCellInst_SboxInst_12_XX_2_ ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_YY_0_ ;
    wire SubCellInst_SboxInst_13_YY_1_ ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_13_XX_1_ ;
    wire SubCellInst_SboxInst_13_XX_2_ ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_YY_0_ ;
    wire SubCellInst_SboxInst_14_YY_1_ ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_14_XX_1_ ;
    wire SubCellInst_SboxInst_14_XX_2_ ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_YY_0_ ;
    wire SubCellInst_SboxInst_15_YY_1_ ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire SubCellInst_SboxInst_15_XX_1_ ;
    wire SubCellInst_SboxInst_15_XX_2_ ;
    wire AddConstXOR_AddConstXOR_XORInst_0_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_3_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_3_n1 ;
    wire MCInst_MCR0_XORInst_0_0_n2 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n2 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n2 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n2 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n2 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n2 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n2 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n2 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n2 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n2 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n2 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n2 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n2 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n2 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n2 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n2 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire MCInst_MCR2_XORInst_0_0_n1 ;
    wire MCInst_MCR2_XORInst_0_1_n1 ;
    wire MCInst_MCR2_XORInst_0_2_n1 ;
    wire MCInst_MCR2_XORInst_0_3_n1 ;
    wire MCInst_MCR2_XORInst_1_0_n1 ;
    wire MCInst_MCR2_XORInst_1_1_n1 ;
    wire MCInst_MCR2_XORInst_1_2_n1 ;
    wire MCInst_MCR2_XORInst_1_3_n1 ;
    wire MCInst_MCR2_XORInst_2_0_n1 ;
    wire MCInst_MCR2_XORInst_2_1_n1 ;
    wire MCInst_MCR2_XORInst_2_2_n1 ;
    wire MCInst_MCR2_XORInst_2_3_n1 ;
    wire MCInst_MCR2_XORInst_3_0_n1 ;
    wire MCInst_MCR2_XORInst_3_1_n1 ;
    wire MCInst_MCR2_XORInst_3_2_n1 ;
    wire MCInst_MCR2_XORInst_3_3_n1 ;
    wire MCInst_MCR3_XORInst_0_0_n1 ;
    wire MCInst_MCR3_XORInst_0_1_n1 ;
    wire MCInst_MCR3_XORInst_0_2_n1 ;
    wire MCInst_MCR3_XORInst_0_3_n1 ;
    wire MCInst_MCR3_XORInst_1_0_n1 ;
    wire MCInst_MCR3_XORInst_1_1_n1 ;
    wire MCInst_MCR3_XORInst_1_2_n1 ;
    wire MCInst_MCR3_XORInst_1_3_n1 ;
    wire MCInst_MCR3_XORInst_2_0_n1 ;
    wire MCInst_MCR3_XORInst_2_1_n1 ;
    wire MCInst_MCR3_XORInst_2_2_n1 ;
    wire MCInst_MCR3_XORInst_2_3_n1 ;
    wire MCInst_MCR3_XORInst_3_0_n1 ;
    wire MCInst_MCR3_XORInst_3_1_n1 ;
    wire MCInst_MCR3_XORInst_3_2_n1 ;
    wire MCInst_MCR3_XORInst_3_3_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire FSMSignalsInst_doneInst_n1 ;
    wire [63:0] MCOutput ;
    wire [63:0] StateRegInput ;
    wire [63:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [5:0] FSMSelected ;
    wire [63:0] TweakeyGeneration_StateRegInput ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U1 ( .a ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .a ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .a ({Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR0_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, SubCellInst_SboxInst_0_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR1_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR3_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR5_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, SubCellInst_SboxInst_0_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR6_U1 ( .a ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}), .b ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, SubCellInst_SboxInst_0_Q6}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, SubCellInst_SboxInst_0_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR8_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, SubCellInst_SboxInst_0_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U1 ( .a ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .a ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, SubCellInst_SboxInst_1_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .a ({Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR0_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, SubCellInst_SboxInst_1_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR1_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, SubCellInst_SboxInst_1_XX_1_}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR3_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, SubCellInst_SboxInst_1_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR5_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR6_U1 ( .a ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, SubCellInst_SboxInst_1_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR8_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, SubCellInst_SboxInst_1_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U1 ( .a ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .a ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .a ({Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR0_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, SubCellInst_SboxInst_2_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR1_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR3_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR5_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, SubCellInst_SboxInst_2_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR6_U1 ( .a ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}), .b ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, SubCellInst_SboxInst_2_Q6}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, SubCellInst_SboxInst_2_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR8_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, SubCellInst_SboxInst_2_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U1 ( .a ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .a ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, SubCellInst_SboxInst_3_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .a ({Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR0_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, SubCellInst_SboxInst_3_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR1_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, SubCellInst_SboxInst_3_XX_1_}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR3_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, SubCellInst_SboxInst_3_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR5_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR6_U1 ( .a ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, SubCellInst_SboxInst_3_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR8_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, SubCellInst_SboxInst_3_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U1 ( .a ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .a ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .a ({Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR0_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, SubCellInst_SboxInst_4_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR1_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR3_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR5_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, SubCellInst_SboxInst_4_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR6_U1 ( .a ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}), .b ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, SubCellInst_SboxInst_4_Q6}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, SubCellInst_SboxInst_4_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR8_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, SubCellInst_SboxInst_4_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U1 ( .a ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .a ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, SubCellInst_SboxInst_5_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .a ({Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR0_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, SubCellInst_SboxInst_5_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR1_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, SubCellInst_SboxInst_5_XX_1_}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR3_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, SubCellInst_SboxInst_5_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR5_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR6_U1 ( .a ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, SubCellInst_SboxInst_5_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR8_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, SubCellInst_SboxInst_5_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U1 ( .a ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .a ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .a ({Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR0_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, SubCellInst_SboxInst_6_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR1_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR3_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR5_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, SubCellInst_SboxInst_6_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR6_U1 ( .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}), .b ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, SubCellInst_SboxInst_6_Q6}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, SubCellInst_SboxInst_6_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR8_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, SubCellInst_SboxInst_6_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U1 ( .a ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .a ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, SubCellInst_SboxInst_7_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .a ({Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR0_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, SubCellInst_SboxInst_7_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR1_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, SubCellInst_SboxInst_7_XX_1_}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR3_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, SubCellInst_SboxInst_7_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR5_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR6_U1 ( .a ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, SubCellInst_SboxInst_7_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR8_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, SubCellInst_SboxInst_7_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U1 ( .a ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .a ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .a ({Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR0_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, SubCellInst_SboxInst_8_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR1_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR3_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR5_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_8_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR6_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}), .b ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_8_Q6}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, SubCellInst_SboxInst_8_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR8_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, SubCellInst_SboxInst_8_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U1 ( .a ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .a ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, SubCellInst_SboxInst_9_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .a ({Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR0_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, SubCellInst_SboxInst_9_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR1_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, SubCellInst_SboxInst_9_XX_1_}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR3_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, SubCellInst_SboxInst_9_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR5_U1 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR6_U1 ( .a ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}), .b ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, SubCellInst_SboxInst_9_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR8_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, SubCellInst_SboxInst_9_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U1 ( .a ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .a ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .a ({Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR0_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, SubCellInst_SboxInst_10_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR1_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR3_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR5_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_10_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR6_U1 ( .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_10_Q6}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, SubCellInst_SboxInst_10_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR8_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, SubCellInst_SboxInst_10_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U1 ( .a ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .a ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, SubCellInst_SboxInst_11_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .a ({Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR0_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, SubCellInst_SboxInst_11_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR1_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, SubCellInst_SboxInst_11_XX_1_}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR3_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, SubCellInst_SboxInst_11_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR5_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR6_U1 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, SubCellInst_SboxInst_11_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR8_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, SubCellInst_SboxInst_11_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U1 ( .a ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .a ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .a ({Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR0_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, SubCellInst_SboxInst_12_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR1_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR3_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR5_U1 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_12_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR6_U1 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_12_Q6}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, SubCellInst_SboxInst_12_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR8_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, SubCellInst_SboxInst_12_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U1 ( .a ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .a ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, SubCellInst_SboxInst_13_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .a ({Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR0_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, SubCellInst_SboxInst_13_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR1_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, SubCellInst_SboxInst_13_XX_1_}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR3_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, SubCellInst_SboxInst_13_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR5_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR6_U1 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, SubCellInst_SboxInst_13_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR8_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, SubCellInst_SboxInst_13_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U1 ( .a ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .a ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .a ({Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR0_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, SubCellInst_SboxInst_14_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR1_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR3_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR5_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_14_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR6_U1 ( .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_14_Q6}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, SubCellInst_SboxInst_14_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR8_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, SubCellInst_SboxInst_14_L2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U1 ( .a ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .a ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, SubCellInst_SboxInst_15_XX_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .a ({Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR0_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, SubCellInst_SboxInst_15_Q0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR1_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, SubCellInst_SboxInst_15_XX_1_}), .c ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR3_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, SubCellInst_SboxInst_15_Q4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR5_U1 ( .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR6_U1 ( .a ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, SubCellInst_SboxInst_15_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR8_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, SubCellInst_SboxInst_15_L2}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[0]}), .a ({Key_s2[0], Key_s1[0], Key_s0[0]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, TweakeyGeneration_StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[1]}), .a ({Key_s2[1], Key_s1[1], Key_s0[1]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, TweakeyGeneration_StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[2]}), .a ({Key_s2[2], Key_s1[2], Key_s0[2]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, TweakeyGeneration_StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[3]}), .a ({Key_s2[3], Key_s1[3], Key_s0[3]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, TweakeyGeneration_StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[4]}), .a ({Key_s2[4], Key_s1[4], Key_s0[4]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, TweakeyGeneration_StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[5]}), .a ({Key_s2[5], Key_s1[5], Key_s0[5]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, TweakeyGeneration_StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[6]}), .a ({Key_s2[6], Key_s1[6], Key_s0[6]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, TweakeyGeneration_StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[7]}), .a ({Key_s2[7], Key_s1[7], Key_s0[7]}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, TweakeyGeneration_StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[8]}), .a ({Key_s2[8], Key_s1[8], Key_s0[8]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, TweakeyGeneration_StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[9]}), .a ({Key_s2[9], Key_s1[9], Key_s0[9]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, TweakeyGeneration_StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[10]}), .a ({Key_s2[10], Key_s1[10], Key_s0[10]}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, TweakeyGeneration_StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[11]}), .a ({Key_s2[11], Key_s1[11], Key_s0[11]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, TweakeyGeneration_StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[12]}), .a ({Key_s2[12], Key_s1[12], Key_s0[12]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, TweakeyGeneration_StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[13]}), .a ({Key_s2[13], Key_s1[13], Key_s0[13]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, TweakeyGeneration_StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[14]}), .a ({Key_s2[14], Key_s1[14], Key_s0[14]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, TweakeyGeneration_StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[15]}), .a ({Key_s2[15], Key_s1[15], Key_s0[15]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, TweakeyGeneration_StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[16]}), .a ({Key_s2[16], Key_s1[16], Key_s0[16]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, TweakeyGeneration_StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_key_Feedback[17]}), .a ({Key_s2[17], Key_s1[17], Key_s0[17]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, TweakeyGeneration_StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, TweakeyGeneration_key_Feedback[18]}), .a ({Key_s2[18], Key_s1[18], Key_s0[18]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, TweakeyGeneration_StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[19]}), .a ({Key_s2[19], Key_s1[19], Key_s0[19]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, TweakeyGeneration_StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_key_Feedback[20]}), .a ({Key_s2[20], Key_s1[20], Key_s0[20]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, TweakeyGeneration_StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, TweakeyGeneration_key_Feedback[21]}), .a ({Key_s2[21], Key_s1[21], Key_s0[21]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, TweakeyGeneration_StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[22]}), .a ({Key_s2[22], Key_s1[22], Key_s0[22]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, TweakeyGeneration_StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_key_Feedback[23]}), .a ({Key_s2[23], Key_s1[23], Key_s0[23]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, TweakeyGeneration_StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, TweakeyGeneration_key_Feedback[24]}), .a ({Key_s2[24], Key_s1[24], Key_s0[24]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, TweakeyGeneration_StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[25]}), .a ({Key_s2[25], Key_s1[25], Key_s0[25]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, TweakeyGeneration_StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_key_Feedback[26]}), .a ({Key_s2[26], Key_s1[26], Key_s0[26]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, TweakeyGeneration_StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, TweakeyGeneration_key_Feedback[27]}), .a ({Key_s2[27], Key_s1[27], Key_s0[27]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, TweakeyGeneration_StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[28]}), .a ({Key_s2[28], Key_s1[28], Key_s0[28]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, TweakeyGeneration_StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_key_Feedback[29]}), .a ({Key_s2[29], Key_s1[29], Key_s0[29]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, TweakeyGeneration_StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, TweakeyGeneration_key_Feedback[30]}), .a ({Key_s2[30], Key_s1[30], Key_s0[30]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, TweakeyGeneration_StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[31]}), .a ({Key_s2[31], Key_s1[31], Key_s0[31]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, TweakeyGeneration_StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_key_Feedback[32]}), .a ({Key_s2[32], Key_s1[32], Key_s0[32]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, TweakeyGeneration_StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, TweakeyGeneration_key_Feedback[33]}), .a ({Key_s2[33], Key_s1[33], Key_s0[33]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, TweakeyGeneration_StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[34]}), .a ({Key_s2[34], Key_s1[34], Key_s0[34]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, TweakeyGeneration_StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_key_Feedback[35]}), .a ({Key_s2[35], Key_s1[35], Key_s0[35]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, TweakeyGeneration_StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, TweakeyGeneration_key_Feedback[36]}), .a ({Key_s2[36], Key_s1[36], Key_s0[36]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, TweakeyGeneration_StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[37]}), .a ({Key_s2[37], Key_s1[37], Key_s0[37]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, TweakeyGeneration_StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_key_Feedback[38]}), .a ({Key_s2[38], Key_s1[38], Key_s0[38]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, TweakeyGeneration_StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, TweakeyGeneration_key_Feedback[39]}), .a ({Key_s2[39], Key_s1[39], Key_s0[39]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, TweakeyGeneration_StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[40]}), .a ({Key_s2[40], Key_s1[40], Key_s0[40]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, TweakeyGeneration_StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_key_Feedback[41]}), .a ({Key_s2[41], Key_s1[41], Key_s0[41]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, TweakeyGeneration_StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, TweakeyGeneration_key_Feedback[42]}), .a ({Key_s2[42], Key_s1[42], Key_s0[42]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, TweakeyGeneration_StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[43]}), .a ({Key_s2[43], Key_s1[43], Key_s0[43]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, TweakeyGeneration_StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_key_Feedback[44]}), .a ({Key_s2[44], Key_s1[44], Key_s0[44]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, TweakeyGeneration_StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, TweakeyGeneration_key_Feedback[45]}), .a ({Key_s2[45], Key_s1[45], Key_s0[45]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, TweakeyGeneration_StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[46]}), .a ({Key_s2[46], Key_s1[46], Key_s0[46]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, TweakeyGeneration_StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_key_Feedback[47]}), .a ({Key_s2[47], Key_s1[47], Key_s0[47]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, TweakeyGeneration_StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, TweakeyGeneration_key_Feedback[48]}), .a ({Key_s2[48], Key_s1[48], Key_s0[48]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, TweakeyGeneration_StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[49]}), .a ({Key_s2[49], Key_s1[49], Key_s0[49]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, TweakeyGeneration_StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_key_Feedback[50]}), .a ({Key_s2[50], Key_s1[50], Key_s0[50]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, TweakeyGeneration_StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, TweakeyGeneration_key_Feedback[51]}), .a ({Key_s2[51], Key_s1[51], Key_s0[51]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, TweakeyGeneration_StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[52]}), .a ({Key_s2[52], Key_s1[52], Key_s0[52]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, TweakeyGeneration_StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_key_Feedback[53]}), .a ({Key_s2[53], Key_s1[53], Key_s0[53]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, TweakeyGeneration_StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, TweakeyGeneration_key_Feedback[54]}), .a ({Key_s2[54], Key_s1[54], Key_s0[54]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, TweakeyGeneration_StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[55]}), .a ({Key_s2[55], Key_s1[55], Key_s0[55]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, TweakeyGeneration_StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_key_Feedback[56]}), .a ({Key_s2[56], Key_s1[56], Key_s0[56]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, TweakeyGeneration_StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, TweakeyGeneration_key_Feedback[57]}), .a ({Key_s2[57], Key_s1[57], Key_s0[57]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, TweakeyGeneration_StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[58]}), .a ({Key_s2[58], Key_s1[58], Key_s0[58]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, TweakeyGeneration_StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_key_Feedback[59]}), .a ({Key_s2[59], Key_s1[59], Key_s0[59]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, TweakeyGeneration_StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, TweakeyGeneration_key_Feedback[60]}), .a ({Key_s2[60], Key_s1[60], Key_s0[60]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, TweakeyGeneration_StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[61]}), .a ({Key_s2[61], Key_s1[61], Key_s0[61]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, TweakeyGeneration_StateRegInput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_key_Feedback[62]}), .a ({Key_s2[62], Key_s1[62], Key_s0[62]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, TweakeyGeneration_StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, TweakeyGeneration_key_Feedback[63]}), .a ({Key_s2[63], Key_s1[63], Key_s0[63]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, TweakeyGeneration_StateRegInput[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMUpdate[0]), .B (1'b1), .Z (FSMSelected[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMUpdate[1]), .B (1'b0), .Z (FSMSelected[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMUpdate[2]), .B (1'b0), .Z (FSMSelected[2]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMUpdate[3]), .B (1'b0), .Z (FSMSelected[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMUpdate[4]), .B (1'b0), .Z (FSMSelected[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMUpdate[5]), .B (1'b0), .Z (FSMSelected[5]) ) ;
    MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .S (FSM[4]), .A (FSMUpdateInst_StateUpdateInst_0_n4), .B (FSM[5]), .Z (FSMUpdate[0]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_0_n3), .ZN (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1 (FSMUpdateInst_StateUpdateInst_0_n2), .A2 (FSMUpdateInst_StateUpdateInst_0_n1), .ZN (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n4), .A2 (FSM[1]), .ZN (FSMUpdate[2]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n3), .A2 (FSM[5]), .ZN (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_2_n2), .ZN (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1 (FSMUpdate[1]), .A2 (FSMUpdateInst_StateUpdateInst_2_n1), .ZN (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n4), .ZN (FSMUpdate[5]) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1 (FSMUpdate[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n3), .ZN (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_5_n2), .ZN (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdateInst_StateUpdateInst_5_n1), .ZN (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1 (FSMSignalsInst_doneInst_n5), .A2 (FSMSignalsInst_doneInst_n4), .ZN (done) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1 (FSM[4]), .A2 (FSM[5]), .ZN (FSMSignalsInst_doneInst_n4) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1 (FSMSignalsInst_doneInst_n3), .A2 (FSMSignalsInst_doneInst_n2), .ZN (FSMSignalsInst_doneInst_n5) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1 (FSMUpdate[4]), .A2 (FSMSignalsInst_doneInst_n1), .ZN (FSMSignalsInst_doneInst_n2) ) ;
    INV_X1 FSMSignalsInst_doneInst_U2 ( .A (FSMUpdate[1]), .ZN (FSMSignalsInst_doneInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1 (FSM[1]), .A2 (FSMUpdate[3]), .ZN (FSMSignalsInst_doneInst_n3) ) ;
    ClockGatingController #(3) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, MCOutput[2]}), .a ({Plaintext_s2[2], Plaintext_s1[2], Plaintext_s0[2]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[3]}), .a ({Plaintext_s2[3], Plaintext_s1[3], Plaintext_s0[3]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, MCOutput[6]}), .a ({Plaintext_s2[6], Plaintext_s1[6], Plaintext_s0[6]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, MCOutput[7]}), .a ({Plaintext_s2[7], Plaintext_s1[7], Plaintext_s0[7]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, MCOutput[10]}), .a ({Plaintext_s2[10], Plaintext_s1[10], Plaintext_s0[10]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, MCOutput[11]}), .a ({Plaintext_s2[11], Plaintext_s1[11], Plaintext_s0[11]}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, MCOutput[14]}), .a ({Plaintext_s2[14], Plaintext_s1[14], Plaintext_s0[14]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCOutput[15]}), .a ({Plaintext_s2[15], Plaintext_s1[15], Plaintext_s0[15]}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, MCOutput[18]}), .a ({Plaintext_s2[18], Plaintext_s1[18], Plaintext_s0[18]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, MCOutput[19]}), .a ({Plaintext_s2[19], Plaintext_s1[19], Plaintext_s0[19]}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, MCOutput[22]}), .a ({Plaintext_s2[22], Plaintext_s1[22], Plaintext_s0[22]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, MCOutput[23]}), .a ({Plaintext_s2[23], Plaintext_s1[23], Plaintext_s0[23]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[26]}), .a ({Plaintext_s2[26], Plaintext_s1[26], Plaintext_s0[26]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCOutput[27]}), .a ({Plaintext_s2[27], Plaintext_s1[27], Plaintext_s0[27]}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, MCOutput[30]}), .a ({Plaintext_s2[30], Plaintext_s1[30], Plaintext_s0[30]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, MCOutput[31]}), .a ({Plaintext_s2[31], Plaintext_s1[31], Plaintext_s0[31]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .a ({Plaintext_s2[34], Plaintext_s1[34], Plaintext_s0[34]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .a ({Plaintext_s2[35], Plaintext_s1[35], Plaintext_s0[35]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .a ({Plaintext_s2[38], Plaintext_s1[38], Plaintext_s0[38]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .a ({Plaintext_s2[39], Plaintext_s1[39], Plaintext_s0[39]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .a ({Plaintext_s2[42], Plaintext_s1[42], Plaintext_s0[42]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .a ({Plaintext_s2[43], Plaintext_s1[43], Plaintext_s0[43]}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .a ({Plaintext_s2[46], Plaintext_s1[46], Plaintext_s0[46]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .a ({Plaintext_s2[47], Plaintext_s1[47], Plaintext_s0[47]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, MCOutput[50]}), .a ({Plaintext_s2[50], Plaintext_s1[50], Plaintext_s0[50]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[51]}), .a ({Plaintext_s2[51], Plaintext_s1[51], Plaintext_s0[51]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, MCOutput[54]}), .a ({Plaintext_s2[54], Plaintext_s1[54], Plaintext_s0[54]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[55]}), .a ({Plaintext_s2[55], Plaintext_s1[55], Plaintext_s0[55]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, MCOutput[58]}), .a ({Plaintext_s2[58], Plaintext_s1[58], Plaintext_s0[58]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, MCOutput[59]}), .a ({Plaintext_s2[59], Plaintext_s1[59], Plaintext_s0[59]}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[62]}), .a ({Plaintext_s2[62], Plaintext_s1[62], Plaintext_s0[62]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCOutput[63]}), .a ({Plaintext_s2[63], Plaintext_s1[63], Plaintext_s0[63]}), .c ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, StateRegInput[63]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, ShiftRowsOutput[7]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_U2 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_YY_0_}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, ShiftRowsOutput[6]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_AND1_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, SubCellInst_SboxInst_0_Q1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR2_U1 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, SubCellInst_SboxInst_0_Q0}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_AND3_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR7_U1 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, SubCellInst_SboxInst_0_L1}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR11_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, SubCellInst_SboxInst_0_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR12_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, SubCellInst_SboxInst_0_L3}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, SubCellInst_SboxInst_0_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR13_U1 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, ShiftRowsOutput[11]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_U2 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_1_YY_0_}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, ShiftRowsOutput[10]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_AND1_U1 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR2_U1 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, SubCellInst_SboxInst_1_Q0}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_1_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_AND3_U1 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, SubCellInst_SboxInst_1_Q4}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR7_U1 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, SubCellInst_SboxInst_1_L1}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, SubCellInst_SboxInst_1_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR11_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR12_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, SubCellInst_SboxInst_1_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR13_U1 ( .a ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, SubCellInst_SboxInst_1_XX_1_}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_1_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, ShiftRowsOutput[15]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_U2 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, SubCellInst_SboxInst_2_YY_0_}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, ShiftRowsOutput[14]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_AND1_U1 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, SubCellInst_SboxInst_2_Q1}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR2_U1 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, SubCellInst_SboxInst_2_Q0}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_AND3_U1 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR7_U1 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, SubCellInst_SboxInst_2_L1}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR11_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_2_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR12_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_2_L3}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_2_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR13_U1 ( .a ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, SubCellInst_SboxInst_2_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, ShiftRowsOutput[3]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_U2 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_3_YY_0_}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, ShiftRowsOutput[2]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_AND1_U1 ( .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR2_U1 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, SubCellInst_SboxInst_3_Q0}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_3_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_AND3_U1 ( .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, SubCellInst_SboxInst_3_Q4}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR7_U1 ( .a ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, SubCellInst_SboxInst_3_L1}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_3_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR11_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR12_U1 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, SubCellInst_SboxInst_3_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR13_U1 ( .a ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, SubCellInst_SboxInst_3_XX_1_}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_3_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_U2 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_4_YY_0_}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_AND1_U1 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, SubCellInst_SboxInst_4_Q1}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR2_U1 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, SubCellInst_SboxInst_4_Q0}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_AND3_U1 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR7_U1 ( .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, SubCellInst_SboxInst_4_L1}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR11_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, SubCellInst_SboxInst_4_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR12_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, SubCellInst_SboxInst_4_L3}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, SubCellInst_SboxInst_4_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR13_U1 ( .a ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_4_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_U2 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, SubCellInst_SboxInst_5_YY_0_}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_AND1_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR2_U1 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, SubCellInst_SboxInst_5_Q0}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, SubCellInst_SboxInst_5_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_AND3_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, SubCellInst_SboxInst_5_Q4}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR7_U1 ( .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, SubCellInst_SboxInst_5_L1}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_5_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR11_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR12_U1 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_5_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR13_U1 ( .a ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, SubCellInst_SboxInst_5_XX_1_}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, SubCellInst_SboxInst_5_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_U2 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, SubCellInst_SboxInst_6_YY_0_}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_AND1_U1 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, SubCellInst_SboxInst_6_Q1}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR2_U1 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, SubCellInst_SboxInst_6_Q0}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_AND3_U1 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR7_U1 ( .a ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, SubCellInst_SboxInst_6_L1}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR11_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, SubCellInst_SboxInst_6_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR12_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, SubCellInst_SboxInst_6_L3}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, SubCellInst_SboxInst_6_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR13_U1 ( .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, SubCellInst_SboxInst_6_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_U2 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, SubCellInst_SboxInst_7_YY_0_}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_AND1_U1 ( .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR2_U1 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, SubCellInst_SboxInst_7_Q0}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, SubCellInst_SboxInst_7_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_AND3_U1 ( .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, SubCellInst_SboxInst_7_Q4}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR7_U1 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, SubCellInst_SboxInst_7_L1}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, SubCellInst_SboxInst_7_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR11_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR12_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, SubCellInst_SboxInst_7_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR13_U1 ( .a ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, SubCellInst_SboxInst_7_XX_1_}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, SubCellInst_SboxInst_7_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, AddRoundConstantOutput[35]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_U2 ( .a ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, SubCellInst_SboxInst_8_YY_0_}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, AddRoundConstantOutput[34]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_AND1_U1 ( .a ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, SubCellInst_SboxInst_8_Q1}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR2_U1 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, SubCellInst_SboxInst_8_Q0}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_AND3_U1 ( .a ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR7_U1 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, SubCellInst_SboxInst_8_L1}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR11_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, SubCellInst_SboxInst_8_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR12_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, SubCellInst_SboxInst_8_L3}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, SubCellInst_SboxInst_8_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR13_U1 ( .a ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, SubCellInst_SboxInst_8_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, AddRoundConstantOutput[39]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_U2 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_9_YY_0_}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, AddRoundConstantOutput[38]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_AND1_U1 ( .a ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR2_U1 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, SubCellInst_SboxInst_9_Q0}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, SubCellInst_SboxInst_9_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_AND3_U1 ( .a ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, SubCellInst_SboxInst_9_Q4}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR7_U1 ( .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, SubCellInst_SboxInst_9_L1}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, SubCellInst_SboxInst_9_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR11_U1 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR12_U1 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, SubCellInst_SboxInst_9_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR13_U1 ( .a ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, SubCellInst_SboxInst_9_XX_1_}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_9_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, AddRoundConstantOutput[43]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_U2 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, SubCellInst_SboxInst_10_YY_0_}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, AddRoundConstantOutput[42]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_AND1_U1 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, SubCellInst_SboxInst_10_Q1}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR2_U1 ( .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, SubCellInst_SboxInst_10_Q0}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_AND3_U1 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR7_U1 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, SubCellInst_SboxInst_10_L1}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR11_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_10_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR12_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_10_L3}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, SubCellInst_SboxInst_10_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR13_U1 ( .a ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, SubCellInst_SboxInst_10_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellOutput[47]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_U2 ( .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, SubCellInst_SboxInst_11_YY_0_}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, SubCellOutput[46]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_AND1_U1 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR2_U1 ( .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, SubCellInst_SboxInst_11_Q0}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_AND3_U1 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, SubCellInst_SboxInst_11_Q4}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR7_U1 ( .a ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, SubCellInst_SboxInst_11_L1}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR11_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, SubCellInst_SboxInst_11_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR12_U1 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, SubCellInst_SboxInst_11_L3}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_11_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR13_U1 ( .a ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, SubCellInst_SboxInst_11_XX_1_}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, SubCellInst_SboxInst_11_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, AddRoundConstantOutput[51]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_U2 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_12_YY_0_}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, AddRoundConstantOutput[50]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_AND1_U1 ( .a ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, SubCellInst_SboxInst_12_Q1}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR2_U1 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, SubCellInst_SboxInst_12_Q0}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_12_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_AND3_U1 ( .a ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR7_U1 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, SubCellInst_SboxInst_12_L1}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, SubCellInst_SboxInst_12_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR11_U1 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR12_U1 ( .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, SubCellInst_SboxInst_12_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR13_U1 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_12_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, AddRoundConstantOutput[55]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_U2 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, SubCellInst_SboxInst_13_YY_0_}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, AddRoundConstantOutput[54]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_AND1_U1 ( .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR2_U1 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, SubCellInst_SboxInst_13_Q0}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_AND3_U1 ( .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, SubCellInst_SboxInst_13_Q4}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR7_U1 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, SubCellInst_SboxInst_13_L1}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR11_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, SubCellInst_SboxInst_13_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR12_U1 ( .a ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, SubCellInst_SboxInst_13_L3}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, SubCellInst_SboxInst_13_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR13_U1 ( .a ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, SubCellInst_SboxInst_13_XX_1_}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, SubCellInst_SboxInst_13_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, AddRoundConstantOutput[59]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_U2 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, SubCellInst_SboxInst_14_YY_0_}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, AddRoundConstantOutput[58]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_AND1_U1 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, SubCellInst_SboxInst_14_Q1}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR2_U1 ( .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, SubCellInst_SboxInst_14_Q0}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, SubCellInst_SboxInst_14_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_AND3_U1 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR7_U1 ( .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, SubCellInst_SboxInst_14_L1}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_14_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR11_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR12_U1 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_14_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR13_U1 ( .a ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, SubCellInst_SboxInst_14_YY_0_}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, SubCellOutput[63]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_U2 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, SubCellInst_SboxInst_15_YY_0_}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, SubCellOutput[62]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_AND1_U1 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR2_U1 ( .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, SubCellInst_SboxInst_15_Q0}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_AND3_U1 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, SubCellInst_SboxInst_15_Q4}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR7_U1 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, SubCellInst_SboxInst_15_L1}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR11_U1 ( .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, SubCellInst_SboxInst_15_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR12_U1 ( .a ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, SubCellInst_SboxInst_15_L3}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, SubCellInst_SboxInst_15_YY_1_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR13_U1 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, SubCellInst_SboxInst_15_XX_1_}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, SubCellInst_SboxInst_15_YY_0_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, AddConstXOR_AddConstXOR_XORInst_0_2_n1}), .b ({1'b0, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, AddRoundConstantOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, SubCellOutput[62]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, AddConstXOR_AddConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, AddConstXOR_AddConstXOR_XORInst_0_3_n1}), .b ({1'b0, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, AddRoundConstantOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, SubCellOutput[63]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, AddConstXOR_AddConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, AddConstXOR_AddConstXOR_XORInst_1_2_n1}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, AddRoundConstantOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, SubCellOutput[46]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, AddConstXOR_AddConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, AddConstXOR_AddConstXOR_XORInst_1_3_n1}), .b ({1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, AddRoundConstantOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellOutput[47]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, AddConstXOR_AddConstXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, AddRoundTweakeyXOR_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[2]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, AddRoundConstantOutput[34]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, AddRoundTweakeyXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, AddRoundTweakeyXOR_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[3]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, ShiftRowsOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, AddRoundConstantOutput[35]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, AddRoundTweakeyXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, AddRoundTweakeyXOR_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[6]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, ShiftRowsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, AddRoundConstantOutput[38]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, AddRoundTweakeyXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, AddRoundTweakeyXOR_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[7]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, AddRoundConstantOutput[39]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, AddRoundTweakeyXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, AddRoundTweakeyXOR_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[10]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, AddRoundConstantOutput[42]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, AddRoundTweakeyXOR_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, AddRoundTweakeyXOR_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[11]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, ShiftRowsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, AddRoundConstantOutput[43]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, AddRoundTweakeyXOR_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, AddRoundTweakeyXOR_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[14]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, ShiftRowsOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, AddRoundConstantOutput[46]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, AddRoundTweakeyXOR_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, AddRoundTweakeyXOR_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[15]}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, ShiftRowsOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, AddRoundConstantOutput[47]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, AddRoundTweakeyXOR_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, TweakeyGeneration_key_Feedback[18]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, AddRoundConstantOutput[50]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, AddRoundTweakeyXOR_XORInst_4_3_n1}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[19]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, AddRoundConstantOutput[51]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, AddRoundTweakeyXOR_XORInst_4_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[22]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, AddRoundConstantOutput[54]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, AddRoundTweakeyXOR_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_key_Feedback[23]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, AddRoundConstantOutput[55]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, AddRoundTweakeyXOR_XORInst_5_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_key_Feedback[26]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, AddRoundConstantOutput[58]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, AddRoundTweakeyXOR_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, TweakeyGeneration_key_Feedback[27]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, AddRoundConstantOutput[59]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, AddRoundTweakeyXOR_XORInst_6_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, TweakeyGeneration_key_Feedback[30]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, AddRoundConstantOutput[62]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, AddRoundTweakeyXOR_XORInst_7_3_n1}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[31]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, AddRoundConstantOutput[63]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, AddRoundTweakeyXOR_XORInst_7_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, MCInst_MCR0_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, MCOutput[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, MCInst_MCR0_XORInst_0_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, MCInst_MCR0_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[51]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, MCInst_MCR0_XORInst_0_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, MCInst_MCR0_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, MCOutput[54]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, MCInst_MCR0_XORInst_1_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, MCInst_MCR0_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[55]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .b ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, MCInst_MCR0_XORInst_1_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U3 ( .a ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, MCInst_MCR0_XORInst_2_2_n2}), .b ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, MCOutput[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, MCInst_MCR0_XORInst_2_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U3 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, MCInst_MCR0_XORInst_2_3_n2}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, MCOutput[59]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, MCInst_MCR0_XORInst_2_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U3 ( .a ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCInst_MCR0_XORInst_3_2_n2}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCInst_MCR0_XORInst_3_2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U3 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, MCInst_MCR0_XORInst_3_3_n2}), .b ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, MCInst_MCR0_XORInst_3_3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, MCOutput[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, MCInst_MCR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, MCOutput[19]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, MCInst_MCR2_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, MCOutput[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, MCInst_MCR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, MCOutput[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, MCInst_MCR2_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, MCInst_MCR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCOutput[27]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, MCInst_MCR2_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, MCOutput[30]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, MCInst_MCR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, MCOutput[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, MCInst_MCR2_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, MCOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, MCOutput[34]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, MCInst_MCR3_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, MCOutput[35]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, MCInst_MCR3_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, MCOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, MCOutput[38]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, MCInst_MCR3_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, MCOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, MCOutput[39]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, MCInst_MCR3_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, MCOutput[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, MCOutput[42]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, MCInst_MCR3_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, MCOutput[11]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, MCOutput[43]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, MCInst_MCR3_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, MCOutput[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, MCOutput[46]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, MCInst_MCR3_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCOutput[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, MCOutput[47]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, MCInst_MCR3_XORInst_3_3_n1}) ) ;

    /* cells in depth 2 */
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, MCOutput[0]}), .a ({Plaintext_s2[0], Plaintext_s1[0], Plaintext_s0[0]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, MCOutput[1]}), .a ({Plaintext_s2[1], Plaintext_s1[1], Plaintext_s0[1]}), .c ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCOutput[4]}), .a ({Plaintext_s2[4], Plaintext_s1[4], Plaintext_s0[4]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCOutput[5]}), .a ({Plaintext_s2[5], Plaintext_s1[5], Plaintext_s0[5]}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, MCOutput[8]}), .a ({Plaintext_s2[8], Plaintext_s1[8], Plaintext_s0[8]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, MCOutput[9]}), .a ({Plaintext_s2[9], Plaintext_s1[9], Plaintext_s0[9]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, MCOutput[12]}), .a ({Plaintext_s2[12], Plaintext_s1[12], Plaintext_s0[12]}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, MCOutput[13]}), .a ({Plaintext_s2[13], Plaintext_s1[13], Plaintext_s0[13]}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, MCOutput[16]}), .a ({Plaintext_s2[16], Plaintext_s1[16], Plaintext_s0[16]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCOutput[17]}), .a ({Plaintext_s2[17], Plaintext_s1[17], Plaintext_s0[17]}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, MCOutput[20]}), .a ({Plaintext_s2[20], Plaintext_s1[20], Plaintext_s0[20]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, MCOutput[21]}), .a ({Plaintext_s2[21], Plaintext_s1[21], Plaintext_s0[21]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, MCOutput[24]}), .a ({Plaintext_s2[24], Plaintext_s1[24], Plaintext_s0[24]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, MCOutput[25]}), .a ({Plaintext_s2[25], Plaintext_s1[25], Plaintext_s0[25]}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, MCOutput[28]}), .a ({Plaintext_s2[28], Plaintext_s1[28], Plaintext_s0[28]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, MCOutput[29]}), .a ({Plaintext_s2[29], Plaintext_s1[29], Plaintext_s0[29]}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .a ({Plaintext_s2[32], Plaintext_s1[32], Plaintext_s0[32]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .a ({Plaintext_s2[33], Plaintext_s1[33], Plaintext_s0[33]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .a ({Plaintext_s2[36], Plaintext_s1[36], Plaintext_s0[36]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .a ({Plaintext_s2[37], Plaintext_s1[37], Plaintext_s0[37]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .a ({Plaintext_s2[40], Plaintext_s1[40], Plaintext_s0[40]}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .a ({Plaintext_s2[41], Plaintext_s1[41], Plaintext_s0[41]}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .a ({Plaintext_s2[44], Plaintext_s1[44], Plaintext_s0[44]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .a ({Plaintext_s2[45], Plaintext_s1[45], Plaintext_s0[45]}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[48]}), .a ({Plaintext_s2[48], Plaintext_s1[48], Plaintext_s0[48]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, MCOutput[49]}), .a ({Plaintext_s2[49], Plaintext_s1[49], Plaintext_s0[49]}), .c ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, MCOutput[52]}), .a ({Plaintext_s2[52], Plaintext_s1[52], Plaintext_s0[52]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCOutput[53]}), .a ({Plaintext_s2[53], Plaintext_s1[53], Plaintext_s0[53]}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, MCOutput[56]}), .a ({Plaintext_s2[56], Plaintext_s1[56], Plaintext_s0[56]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCOutput[57]}), .a ({Plaintext_s2[57], Plaintext_s1[57], Plaintext_s0[57]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCOutput[60]}), .a ({Plaintext_s2[60], Plaintext_s1[60], Plaintext_s0[60]}), .c ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) PlaintextMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCOutput[61]}), .a ({Plaintext_s2[61], Plaintext_s1[61], Plaintext_s0[61]}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, StateRegInput[61]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_AND2_U1 ( .a ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, SubCellInst_SboxInst_0_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR4_U1 ( .a ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, SubCellInst_SboxInst_0_T1}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_AND4_U1 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, SubCellInst_SboxInst_0_Q6}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_0_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR9_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, SubCellInst_SboxInst_0_L2}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, SubCellInst_SboxInst_0_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR10_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_0_T3}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, ShiftRowsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, SubCellInst_SboxInst_0_YY_3}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, ShiftRowsOutput[5]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_AND2_U1 ( .a ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_1_Q2}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_1_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR4_U1 ( .a ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_1_T1}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_AND4_U1 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, SubCellInst_SboxInst_1_Q7}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, SubCellInst_SboxInst_1_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR9_U1 ( .a ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, SubCellInst_SboxInst_1_L2}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR10_U1 ( .a ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, SubCellInst_SboxInst_1_T3}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, ShiftRowsOutput[9]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_AND2_U1 ( .a ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, SubCellInst_SboxInst_2_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR4_U1 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, SubCellInst_SboxInst_2_T1}), .b ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_AND4_U1 ( .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, SubCellInst_SboxInst_2_Q6}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, SubCellInst_SboxInst_2_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR9_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, SubCellInst_SboxInst_2_L2}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR10_U1 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, SubCellInst_SboxInst_2_T3}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, ShiftRowsOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[13]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_AND2_U1 ( .a ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_3_Q2}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, SubCellInst_SboxInst_3_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR4_U1 ( .a ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, SubCellInst_SboxInst_3_T1}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_AND4_U1 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_3_Q7}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_3_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR9_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, SubCellInst_SboxInst_3_L2}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR10_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_3_T3}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, ShiftRowsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, ShiftRowsOutput[1]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_AND2_U1 ( .a ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, SubCellInst_SboxInst_4_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR4_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, SubCellInst_SboxInst_4_T1}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_AND4_U1 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, SubCellInst_SboxInst_4_Q6}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, SubCellInst_SboxInst_4_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR9_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, SubCellInst_SboxInst_4_L2}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR10_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, SubCellInst_SboxInst_4_T3}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_AND2_U1 ( .a ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, SubCellInst_SboxInst_5_Q2}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, SubCellInst_SboxInst_5_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR4_U1 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, SubCellInst_SboxInst_5_T1}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_AND4_U1 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_5_Q7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, SubCellInst_SboxInst_5_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR9_U1 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, SubCellInst_SboxInst_5_L2}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR10_U1 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, SubCellInst_SboxInst_5_T3}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_AND2_U1 ( .a ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, SubCellInst_SboxInst_6_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR4_U1 ( .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, SubCellInst_SboxInst_6_T1}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_AND4_U1 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, SubCellInst_SboxInst_6_Q6}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, SubCellInst_SboxInst_6_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR9_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, SubCellInst_SboxInst_6_L2}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR10_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, SubCellInst_SboxInst_6_T3}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_AND2_U1 ( .a ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, SubCellInst_SboxInst_7_Q2}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_7_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR4_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_7_T1}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_AND4_U1 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, SubCellInst_SboxInst_7_Q7}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, SubCellInst_SboxInst_7_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR9_U1 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, SubCellInst_SboxInst_7_L2}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR10_U1 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, SubCellInst_SboxInst_7_T3}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellOutput[29]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_AND2_U1 ( .a ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR4_U1 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_AND4_U1 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_8_Q6}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR9_U1 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, SubCellInst_SboxInst_8_L2}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, SubCellInst_SboxInst_8_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR10_U1 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, AddRoundConstantOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, SubCellInst_SboxInst_8_YY_3}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, AddRoundConstantOutput[33]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_AND2_U1 ( .a ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, SubCellInst_SboxInst_9_Q2}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, SubCellInst_SboxInst_9_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR4_U1 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, SubCellInst_SboxInst_9_T1}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_AND4_U1 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, SubCellInst_SboxInst_9_Q7}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_9_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR9_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, SubCellInst_SboxInst_9_L2}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR10_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_9_T3}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, AddRoundConstantOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, AddRoundConstantOutput[37]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_AND2_U1 ( .a ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_10_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR4_U1 ( .a ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_10_T1}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_AND4_U1 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_10_Q6}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, SubCellInst_SboxInst_10_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR9_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, SubCellInst_SboxInst_10_L2}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR10_U1 ( .a ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, SubCellInst_SboxInst_10_T3}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, AddRoundConstantOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .a ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, AddRoundConstantOutput[41]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_AND2_U1 ( .a ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, SubCellInst_SboxInst_11_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR4_U1 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, SubCellInst_SboxInst_11_T1}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_AND4_U1 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, SubCellInst_SboxInst_11_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR9_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, SubCellInst_SboxInst_11_L2}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR10_U1 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, SubCellInst_SboxInst_11_T3}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, SubCellOutput[45]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_AND2_U1 ( .a ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_12_Q2}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, SubCellInst_SboxInst_12_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR4_U1 ( .a ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, SubCellInst_SboxInst_12_T1}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_AND4_U1 ( .a ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_12_Q6}), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, SubCellInst_SboxInst_12_Q7}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR9_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, SubCellInst_SboxInst_12_L2}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR10_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_T3}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, AddRoundConstantOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, AddRoundConstantOutput[49]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_AND2_U1 ( .a ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, SubCellInst_SboxInst_13_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR4_U1 ( .a ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, SubCellInst_SboxInst_13_T1}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_AND4_U1 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, SubCellInst_SboxInst_13_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR9_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, SubCellInst_SboxInst_13_L2}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR10_U1 ( .a ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, SubCellInst_SboxInst_13_T3}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, AddRoundConstantOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, AddRoundConstantOutput[53]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_AND2_U1 ( .a ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, SubCellInst_SboxInst_14_Q2}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, SubCellInst_SboxInst_14_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR4_U1 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, SubCellInst_SboxInst_14_T1}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_AND4_U1 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_14_Q6}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_14_Q7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, SubCellInst_SboxInst_14_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR9_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, SubCellInst_SboxInst_14_L2}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR10_U1 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, SubCellInst_SboxInst_14_T3}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, AddRoundConstantOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, AddRoundConstantOutput[57]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_AND2_U1 ( .a ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, SubCellInst_SboxInst_15_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR4_U1 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, SubCellInst_SboxInst_15_T1}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_AND4_U1 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, SubCellInst_SboxInst_15_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR9_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, SubCellInst_SboxInst_15_L2}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR10_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, SubCellInst_SboxInst_15_T3}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, SubCellOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, SubCellOutput[61]}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) AddConstXOR_U2 ( .a ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellOutput[29]}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, AddConstXOR_AddConstXOR_XORInst_0_0_n1}), .b ({1'b0, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, AddRoundConstantOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, SubCellOutput[60]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, AddConstXOR_AddConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1}), .b ({1'b0, 1'b0, FSM[1]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, AddRoundConstantOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, SubCellOutput[61]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, AddConstXOR_AddConstXOR_XORInst_1_0_n1}), .b ({1'b0, 1'b0, FSM[4]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, AddRoundConstantOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellOutput[44]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, AddConstXOR_AddConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1}), .b ({1'b0, 1'b0, FSM[5]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, AddRoundConstantOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, SubCellOutput[45]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[0]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, ShiftRowsOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, AddRoundConstantOutput[32]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[1]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, ShiftRowsOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, AddRoundConstantOutput[33]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[4]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, ShiftRowsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, AddRoundConstantOutput[36]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[5]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, AddRoundConstantOutput[37]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[8]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, AddRoundConstantOutput[40]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[9]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, AddRoundConstantOutput[41]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[12]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, AddRoundConstantOutput[44]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[13]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, ShiftRowsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, AddRoundConstantOutput[45]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, AddRoundTweakeyXOR_XORInst_4_0_n1}), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[16]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, AddRoundConstantOutput[48]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, AddRoundTweakeyXOR_XORInst_4_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1}), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_key_Feedback[17]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, AddRoundConstantOutput[49]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, AddRoundTweakeyXOR_XORInst_5_0_n1}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_key_Feedback[20]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, AddRoundConstantOutput[52]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, AddRoundTweakeyXOR_XORInst_5_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, TweakeyGeneration_key_Feedback[21]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, AddRoundConstantOutput[53]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, AddRoundTweakeyXOR_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, TweakeyGeneration_key_Feedback[24]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, AddRoundConstantOutput[56]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, AddRoundTweakeyXOR_XORInst_6_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[25]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, AddRoundConstantOutput[57]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, AddRoundTweakeyXOR_XORInst_7_0_n1}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[28]}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, AddRoundConstantOutput[60]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, AddRoundTweakeyXOR_XORInst_7_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_key_Feedback[29]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, AddRoundConstantOutput[61]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, MCInst_MCR0_XORInst_0_0_n1}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, MCInst_MCR0_XORInst_0_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, MCInst_MCR0_XORInst_0_1_n1}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, MCOutput[49]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, MCInst_MCR0_XORInst_0_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, MCInst_MCR0_XORInst_1_0_n1}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, MCOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, MCInst_MCR0_XORInst_1_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, MCInst_MCR0_XORInst_1_1_n1}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCOutput[53]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, MCInst_MCR0_XORInst_1_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U3 ( .a ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2}), .b ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, MCInst_MCR0_XORInst_2_0_n1}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, MCOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, MCInst_MCR0_XORInst_2_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U3 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, MCInst_MCR0_XORInst_2_1_n1}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, MCInst_MCR0_XORInst_2_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U3 ( .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, MCInst_MCR0_XORInst_3_0_n1}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, MCInst_MCR0_XORInst_3_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U3 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, MCInst_MCR0_XORInst_3_1_n1}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, MCInst_MCR0_XORInst_3_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, MCInst_MCR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, MCOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, MCInst_MCR2_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCOutput[17]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCInst_MCR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, MCOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCInst_MCR2_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, MCOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, MCInst_MCR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, MCOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, MCInst_MCR2_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, MCOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCInst_MCR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, MCOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCInst_MCR2_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, MCOutput[29]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, MCInst_MCR3_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, MCOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, MCOutput[32]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, MCInst_MCR3_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, MCOutput[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[33]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, MCInst_MCR3_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, MCOutput[36]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, MCInst_MCR3_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, MCOutput[37]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCInst_MCR3_XORInst_2_0_n1}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, MCOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, MCOutput[40]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCInst_MCR3_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, MCOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, MCOutput[41]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, MCInst_MCR3_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, MCOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, MCOutput[44]}), .c ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, MCInst_MCR3_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, MCOutput[13]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCOutput[45]}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, StateRegInput[63]}), .Q ({Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, StateRegInput[62]}), .Q ({Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, StateRegInput[61]}), .Q ({Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, StateRegInput[60]}), .Q ({Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, StateRegInput[59]}), .Q ({Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, StateRegInput[58]}), .Q ({Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, StateRegInput[57]}), .Q ({Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, StateRegInput[56]}), .Q ({Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, StateRegInput[55]}), .Q ({Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, StateRegInput[54]}), .Q ({Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, StateRegInput[53]}), .Q ({Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, StateRegInput[52]}), .Q ({Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, StateRegInput[51]}), .Q ({Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, StateRegInput[50]}), .Q ({Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, StateRegInput[49]}), .Q ({Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, StateRegInput[48]}), .Q ({Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, StateRegInput[47]}), .Q ({Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, StateRegInput[46]}), .Q ({Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, StateRegInput[45]}), .Q ({Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, StateRegInput[44]}), .Q ({Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, StateRegInput[43]}), .Q ({Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, StateRegInput[42]}), .Q ({Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, StateRegInput[41]}), .Q ({Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, StateRegInput[40]}), .Q ({Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, StateRegInput[39]}), .Q ({Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, StateRegInput[38]}), .Q ({Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, StateRegInput[37]}), .Q ({Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, StateRegInput[36]}), .Q ({Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, StateRegInput[35]}), .Q ({Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, StateRegInput[34]}), .Q ({Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, StateRegInput[33]}), .Q ({Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, StateRegInput[32]}), .Q ({Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, StateRegInput[31]}), .Q ({Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, StateRegInput[30]}), .Q ({Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, StateRegInput[29]}), .Q ({Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, StateRegInput[28]}), .Q ({Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, StateRegInput[27]}), .Q ({Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, StateRegInput[26]}), .Q ({Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, StateRegInput[25]}), .Q ({Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, StateRegInput[24]}), .Q ({Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, StateRegInput[23]}), .Q ({Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, StateRegInput[22]}), .Q ({Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, StateRegInput[21]}), .Q ({Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, StateRegInput[20]}), .Q ({Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, StateRegInput[19]}), .Q ({Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, StateRegInput[18]}), .Q ({Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, StateRegInput[17]}), .Q ({Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, StateRegInput[16]}), .Q ({Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, StateRegInput[15]}), .Q ({Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, StateRegInput[14]}), .Q ({Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, StateRegInput[13]}), .Q ({Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, StateRegInput[12]}), .Q ({Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, StateRegInput[11]}), .Q ({Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, StateRegInput[10]}), .Q ({Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, StateRegInput[9]}), .Q ({Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, StateRegInput[8]}), .Q ({Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, StateRegInput[7]}), .Q ({Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, StateRegInput[6]}), .Q ({Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, StateRegInput[5]}), .Q ({Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, StateRegInput[4]}), .Q ({Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, StateRegInput[3]}), .Q ({Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, StateRegInput[2]}), .Q ({Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, StateRegInput[1]}), .Q ({Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, StateRegInput[0]}), .Q ({Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, TweakeyGeneration_StateRegInput[63]}), .Q ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, TweakeyGeneration_StateRegInput[62]}), .Q ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, TweakeyGeneration_key_Feedback[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, TweakeyGeneration_StateRegInput[61]}), .Q ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_key_Feedback[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, TweakeyGeneration_StateRegInput[60]}), .Q ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, TweakeyGeneration_StateRegInput[59]}), .Q ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, TweakeyGeneration_key_Feedback[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, TweakeyGeneration_StateRegInput[58]}), .Q ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_key_Feedback[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, TweakeyGeneration_StateRegInput[57]}), .Q ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, TweakeyGeneration_StateRegInput[56]}), .Q ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, TweakeyGeneration_key_Feedback[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, TweakeyGeneration_StateRegInput[55]}), .Q ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_key_Feedback[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, TweakeyGeneration_StateRegInput[54]}), .Q ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, TweakeyGeneration_StateRegInput[53]}), .Q ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, TweakeyGeneration_key_Feedback[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, TweakeyGeneration_StateRegInput[52]}), .Q ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_key_Feedback[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, TweakeyGeneration_StateRegInput[51]}), .Q ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, TweakeyGeneration_StateRegInput[50]}), .Q ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, TweakeyGeneration_key_Feedback[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, TweakeyGeneration_StateRegInput[49]}), .Q ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_key_Feedback[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, TweakeyGeneration_StateRegInput[48]}), .Q ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, TweakeyGeneration_StateRegInput[47]}), .Q ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, TweakeyGeneration_key_Feedback[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, TweakeyGeneration_StateRegInput[46]}), .Q ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, TweakeyGeneration_key_Feedback[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, TweakeyGeneration_StateRegInput[45]}), .Q ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, TweakeyGeneration_key_Feedback[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, TweakeyGeneration_StateRegInput[44]}), .Q ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, TweakeyGeneration_key_Feedback[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, TweakeyGeneration_StateRegInput[43]}), .Q ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, TweakeyGeneration_key_Feedback[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, TweakeyGeneration_StateRegInput[42]}), .Q ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, TweakeyGeneration_key_Feedback[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, TweakeyGeneration_StateRegInput[41]}), .Q ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, TweakeyGeneration_key_Feedback[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, TweakeyGeneration_StateRegInput[40]}), .Q ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, TweakeyGeneration_key_Feedback[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, TweakeyGeneration_StateRegInput[39]}), .Q ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, TweakeyGeneration_key_Feedback[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, TweakeyGeneration_StateRegInput[38]}), .Q ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, TweakeyGeneration_key_Feedback[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, TweakeyGeneration_StateRegInput[37]}), .Q ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, TweakeyGeneration_key_Feedback[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, TweakeyGeneration_StateRegInput[36]}), .Q ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, TweakeyGeneration_key_Feedback[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, TweakeyGeneration_StateRegInput[35]}), .Q ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, TweakeyGeneration_key_Feedback[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, TweakeyGeneration_StateRegInput[34]}), .Q ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, TweakeyGeneration_key_Feedback[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, TweakeyGeneration_StateRegInput[33]}), .Q ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, TweakeyGeneration_key_Feedback[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, TweakeyGeneration_StateRegInput[32]}), .Q ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, TweakeyGeneration_key_Feedback[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, TweakeyGeneration_StateRegInput[31]}), .Q ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, TweakeyGeneration_StateRegInput[30]}), .Q ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, TweakeyGeneration_key_Feedback[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, TweakeyGeneration_StateRegInput[29]}), .Q ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_key_Feedback[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, TweakeyGeneration_StateRegInput[28]}), .Q ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, TweakeyGeneration_StateRegInput[27]}), .Q ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, TweakeyGeneration_key_Feedback[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, TweakeyGeneration_StateRegInput[26]}), .Q ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_key_Feedback[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, TweakeyGeneration_StateRegInput[25]}), .Q ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, TweakeyGeneration_StateRegInput[24]}), .Q ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, TweakeyGeneration_key_Feedback[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, TweakeyGeneration_StateRegInput[23]}), .Q ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_key_Feedback[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, TweakeyGeneration_StateRegInput[22]}), .Q ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, TweakeyGeneration_StateRegInput[21]}), .Q ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, TweakeyGeneration_key_Feedback[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, TweakeyGeneration_StateRegInput[20]}), .Q ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_key_Feedback[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, TweakeyGeneration_StateRegInput[19]}), .Q ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_key_Feedback[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, TweakeyGeneration_StateRegInput[18]}), .Q ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, TweakeyGeneration_StateRegInput[17]}), .Q ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, TweakeyGeneration_key_Feedback[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, TweakeyGeneration_StateRegInput[16]}), .Q ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_key_Feedback[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, TweakeyGeneration_StateRegInput[15]}), .Q ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, TweakeyGeneration_key_Feedback[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, TweakeyGeneration_StateRegInput[14]}), .Q ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_key_Feedback[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, TweakeyGeneration_StateRegInput[13]}), .Q ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, TweakeyGeneration_StateRegInput[12]}), .Q ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, TweakeyGeneration_key_Feedback[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, TweakeyGeneration_StateRegInput[11]}), .Q ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, TweakeyGeneration_key_Feedback[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, TweakeyGeneration_StateRegInput[10]}), .Q ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_key_Feedback[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, TweakeyGeneration_StateRegInput[9]}), .Q ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, TweakeyGeneration_StateRegInput[8]}), .Q ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, TweakeyGeneration_key_Feedback[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, TweakeyGeneration_StateRegInput[7]}), .Q ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, TweakeyGeneration_StateRegInput[6]}), .Q ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, TweakeyGeneration_key_Feedback[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, TweakeyGeneration_StateRegInput[5]}), .Q ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_key_Feedback[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, TweakeyGeneration_StateRegInput[4]}), .Q ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, TweakeyGeneration_StateRegInput[3]}), .Q ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_key_Feedback[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, TweakeyGeneration_StateRegInput[2]}), .Q ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, TweakeyGeneration_StateRegInput[1]}), .Q ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, TweakeyGeneration_key_Feedback[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, TweakeyGeneration_StateRegInput[0]}), .Q ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_key_Feedback[56]}) ) ;
    DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (FSMSelected[5]), .Q (FSM[5]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (FSMSelected[4]), .Q (FSM[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (FSMSelected[3]), .Q (FSMUpdate[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (FSMSelected[2]), .Q (FSMUpdate[3]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (FSMSelected[1]), .Q (FSM[1]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (FSMSelected[0]), .Q (FSMUpdate[1]), .QN () ) ;
endmodule
