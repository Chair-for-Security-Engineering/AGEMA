/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d4 (SI_s0, clk, SI_s1, SI_s2, SI_s3, SI_s4, Fresh, SO_s0, SO_s1, SO_s2, SO_s3, SO_s4);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [7:0] SI_s4 ;
    input [8789:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    output [7:0] SO_s4 ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7783 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7786 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7789 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7792 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7795 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7798 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7801 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7804 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7807 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7810 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7813 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7816 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7819 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7822 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7825 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7828 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7831 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7834 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7837 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7840 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_17078 ;
    wire signal_17079 ;
    wire signal_17080 ;
    wire signal_17081 ;
    wire signal_17082 ;
    wire signal_17083 ;
    wire signal_17084 ;
    wire signal_17085 ;
    wire signal_17086 ;
    wire signal_17087 ;
    wire signal_17088 ;
    wire signal_17089 ;
    wire signal_17090 ;
    wire signal_17091 ;
    wire signal_17092 ;
    wire signal_17093 ;
    wire signal_17094 ;
    wire signal_17095 ;
    wire signal_17096 ;
    wire signal_17097 ;
    wire signal_17098 ;
    wire signal_17099 ;
    wire signal_17100 ;
    wire signal_17101 ;
    wire signal_17102 ;
    wire signal_17103 ;
    wire signal_17104 ;
    wire signal_17105 ;
    wire signal_17106 ;
    wire signal_17107 ;
    wire signal_17108 ;
    wire signal_17109 ;
    wire signal_17110 ;
    wire signal_17111 ;
    wire signal_17112 ;
    wire signal_17113 ;
    wire signal_17114 ;
    wire signal_17115 ;
    wire signal_17116 ;
    wire signal_17117 ;
    wire signal_17118 ;
    wire signal_17119 ;
    wire signal_17120 ;
    wire signal_17121 ;
    wire signal_17122 ;
    wire signal_17123 ;
    wire signal_17124 ;
    wire signal_17125 ;
    wire signal_17126 ;
    wire signal_17127 ;
    wire signal_17128 ;
    wire signal_17129 ;
    wire signal_17130 ;
    wire signal_17131 ;
    wire signal_17132 ;
    wire signal_17133 ;
    wire signal_17134 ;
    wire signal_17135 ;
    wire signal_17136 ;
    wire signal_17137 ;
    wire signal_17138 ;
    wire signal_17139 ;
    wire signal_17140 ;
    wire signal_17141 ;
    wire signal_17142 ;
    wire signal_17143 ;
    wire signal_17144 ;
    wire signal_17145 ;
    wire signal_17146 ;
    wire signal_17147 ;
    wire signal_17148 ;
    wire signal_17149 ;
    wire signal_17150 ;
    wire signal_17151 ;
    wire signal_17152 ;
    wire signal_17153 ;
    wire signal_17154 ;
    wire signal_17155 ;
    wire signal_17156 ;
    wire signal_17157 ;
    wire signal_17158 ;
    wire signal_17159 ;
    wire signal_17160 ;
    wire signal_17161 ;
    wire signal_17162 ;
    wire signal_17163 ;
    wire signal_17164 ;
    wire signal_17165 ;
    wire signal_17166 ;
    wire signal_17167 ;
    wire signal_17168 ;
    wire signal_17169 ;
    wire signal_17170 ;
    wire signal_17171 ;
    wire signal_17172 ;
    wire signal_17173 ;
    wire signal_17174 ;
    wire signal_17175 ;
    wire signal_17176 ;
    wire signal_17177 ;
    wire signal_17178 ;
    wire signal_17179 ;
    wire signal_17180 ;
    wire signal_17181 ;
    wire signal_17182 ;
    wire signal_17183 ;
    wire signal_17184 ;
    wire signal_17185 ;
    wire signal_17186 ;
    wire signal_17187 ;
    wire signal_17188 ;
    wire signal_17189 ;
    wire signal_17190 ;
    wire signal_17191 ;
    wire signal_17192 ;
    wire signal_17193 ;
    wire signal_17194 ;
    wire signal_17195 ;
    wire signal_17196 ;
    wire signal_17197 ;
    wire signal_17198 ;
    wire signal_17199 ;
    wire signal_17200 ;
    wire signal_17201 ;
    wire signal_17202 ;
    wire signal_17203 ;
    wire signal_17204 ;
    wire signal_17205 ;
    wire signal_17206 ;
    wire signal_17207 ;
    wire signal_17208 ;
    wire signal_17209 ;
    wire signal_17210 ;
    wire signal_17211 ;
    wire signal_17212 ;
    wire signal_17213 ;
    wire signal_17214 ;
    wire signal_17215 ;
    wire signal_17216 ;
    wire signal_17217 ;
    wire signal_17218 ;
    wire signal_17219 ;
    wire signal_17220 ;
    wire signal_17221 ;
    wire signal_17222 ;
    wire signal_17223 ;
    wire signal_17224 ;
    wire signal_17225 ;
    wire signal_17226 ;
    wire signal_17227 ;
    wire signal_17228 ;
    wire signal_17229 ;
    wire signal_17230 ;
    wire signal_17231 ;
    wire signal_17232 ;
    wire signal_17233 ;
    wire signal_17234 ;
    wire signal_17235 ;
    wire signal_17236 ;
    wire signal_17237 ;
    wire signal_17238 ;
    wire signal_17239 ;
    wire signal_17240 ;
    wire signal_17241 ;
    wire signal_17242 ;
    wire signal_17243 ;
    wire signal_17244 ;
    wire signal_17245 ;
    wire signal_17246 ;
    wire signal_17247 ;
    wire signal_17248 ;
    wire signal_17249 ;
    wire signal_17250 ;
    wire signal_17251 ;
    wire signal_17252 ;
    wire signal_17253 ;
    wire signal_17254 ;
    wire signal_17255 ;
    wire signal_17256 ;
    wire signal_17257 ;
    wire signal_17258 ;
    wire signal_17259 ;
    wire signal_17260 ;
    wire signal_17261 ;
    wire signal_17262 ;
    wire signal_17263 ;
    wire signal_17264 ;
    wire signal_17265 ;
    wire signal_17266 ;
    wire signal_17267 ;
    wire signal_17268 ;
    wire signal_17269 ;
    wire signal_17270 ;
    wire signal_17271 ;
    wire signal_17272 ;
    wire signal_17273 ;
    wire signal_17274 ;
    wire signal_17275 ;
    wire signal_17276 ;
    wire signal_17277 ;
    wire signal_17278 ;
    wire signal_17279 ;
    wire signal_17280 ;
    wire signal_17281 ;
    wire signal_17282 ;
    wire signal_17283 ;
    wire signal_17284 ;
    wire signal_17285 ;
    wire signal_17286 ;
    wire signal_17287 ;
    wire signal_17288 ;
    wire signal_17289 ;
    wire signal_17290 ;
    wire signal_17291 ;
    wire signal_17292 ;
    wire signal_17293 ;
    wire signal_17294 ;
    wire signal_17295 ;
    wire signal_17296 ;
    wire signal_17297 ;
    wire signal_17298 ;
    wire signal_17299 ;
    wire signal_17300 ;
    wire signal_17301 ;
    wire signal_17302 ;
    wire signal_17303 ;
    wire signal_17304 ;
    wire signal_17305 ;
    wire signal_17306 ;
    wire signal_17307 ;
    wire signal_17308 ;
    wire signal_17309 ;
    wire signal_17310 ;
    wire signal_17311 ;
    wire signal_17312 ;
    wire signal_17313 ;
    wire signal_17314 ;
    wire signal_17315 ;
    wire signal_17316 ;
    wire signal_17317 ;
    wire signal_17318 ;
    wire signal_17319 ;
    wire signal_17320 ;
    wire signal_17321 ;
    wire signal_17322 ;
    wire signal_17323 ;
    wire signal_17324 ;
    wire signal_17325 ;
    wire signal_17326 ;
    wire signal_17327 ;
    wire signal_17328 ;
    wire signal_17329 ;
    wire signal_17330 ;
    wire signal_17331 ;
    wire signal_17332 ;
    wire signal_17333 ;
    wire signal_17334 ;
    wire signal_17335 ;
    wire signal_17336 ;
    wire signal_17337 ;
    wire signal_17338 ;
    wire signal_17339 ;
    wire signal_17340 ;
    wire signal_17341 ;
    wire signal_17342 ;
    wire signal_17343 ;
    wire signal_17344 ;
    wire signal_17345 ;
    wire signal_17346 ;
    wire signal_17347 ;
    wire signal_17348 ;
    wire signal_17349 ;
    wire signal_17350 ;
    wire signal_17351 ;
    wire signal_17352 ;
    wire signal_17353 ;
    wire signal_17354 ;
    wire signal_17355 ;
    wire signal_17356 ;
    wire signal_17357 ;
    wire signal_17358 ;
    wire signal_17359 ;
    wire signal_17360 ;
    wire signal_17361 ;
    wire signal_17362 ;
    wire signal_17363 ;
    wire signal_17364 ;
    wire signal_17365 ;
    wire signal_17366 ;
    wire signal_17367 ;
    wire signal_17368 ;
    wire signal_17369 ;
    wire signal_17370 ;
    wire signal_17371 ;
    wire signal_17372 ;
    wire signal_17373 ;
    wire signal_17374 ;
    wire signal_17375 ;
    wire signal_17376 ;
    wire signal_17377 ;
    wire signal_17378 ;
    wire signal_17379 ;
    wire signal_17380 ;
    wire signal_17381 ;
    wire signal_17382 ;
    wire signal_17383 ;
    wire signal_17384 ;
    wire signal_17385 ;
    wire signal_17386 ;
    wire signal_17387 ;
    wire signal_17388 ;
    wire signal_17389 ;
    wire signal_17390 ;
    wire signal_17391 ;
    wire signal_17392 ;
    wire signal_17393 ;
    wire signal_17394 ;
    wire signal_17395 ;
    wire signal_17396 ;
    wire signal_17397 ;
    wire signal_17398 ;
    wire signal_17399 ;
    wire signal_17400 ;
    wire signal_17401 ;
    wire signal_17402 ;
    wire signal_17403 ;
    wire signal_17404 ;
    wire signal_17405 ;
    wire signal_17406 ;
    wire signal_17407 ;
    wire signal_17408 ;
    wire signal_17409 ;
    wire signal_17410 ;
    wire signal_17411 ;
    wire signal_17412 ;
    wire signal_17413 ;
    wire signal_17414 ;
    wire signal_17415 ;
    wire signal_17416 ;
    wire signal_17417 ;
    wire signal_17418 ;
    wire signal_17419 ;
    wire signal_17420 ;
    wire signal_17421 ;
    wire signal_17422 ;
    wire signal_17423 ;
    wire signal_17424 ;
    wire signal_17425 ;
    wire signal_17426 ;
    wire signal_17427 ;
    wire signal_17428 ;
    wire signal_17429 ;
    wire signal_17430 ;
    wire signal_17431 ;
    wire signal_17432 ;
    wire signal_17433 ;
    wire signal_17434 ;
    wire signal_17435 ;
    wire signal_17436 ;
    wire signal_17437 ;
    wire signal_17438 ;
    wire signal_17439 ;
    wire signal_17440 ;
    wire signal_17441 ;
    wire signal_17442 ;
    wire signal_17443 ;
    wire signal_17444 ;
    wire signal_17445 ;
    wire signal_17446 ;
    wire signal_17447 ;
    wire signal_17448 ;
    wire signal_17449 ;
    wire signal_17450 ;
    wire signal_17451 ;
    wire signal_17452 ;
    wire signal_17453 ;
    wire signal_17454 ;
    wire signal_17455 ;
    wire signal_17456 ;
    wire signal_17457 ;
    wire signal_17458 ;
    wire signal_17459 ;
    wire signal_17460 ;
    wire signal_17461 ;
    wire signal_17462 ;
    wire signal_17463 ;
    wire signal_17464 ;
    wire signal_17465 ;
    wire signal_17466 ;
    wire signal_17467 ;
    wire signal_17468 ;
    wire signal_17469 ;
    wire signal_17470 ;
    wire signal_17471 ;
    wire signal_17472 ;
    wire signal_17473 ;
    wire signal_17474 ;
    wire signal_17475 ;
    wire signal_17476 ;
    wire signal_17477 ;
    wire signal_17478 ;
    wire signal_17479 ;
    wire signal_17480 ;
    wire signal_17481 ;
    wire signal_17482 ;
    wire signal_17483 ;
    wire signal_17484 ;
    wire signal_17485 ;
    wire signal_17486 ;
    wire signal_17487 ;
    wire signal_17488 ;
    wire signal_17489 ;
    wire signal_17490 ;
    wire signal_17491 ;
    wire signal_17492 ;
    wire signal_17493 ;
    wire signal_17494 ;
    wire signal_17495 ;
    wire signal_17496 ;
    wire signal_17497 ;
    wire signal_17498 ;
    wire signal_17499 ;
    wire signal_17500 ;
    wire signal_17501 ;
    wire signal_17502 ;
    wire signal_17503 ;
    wire signal_17504 ;
    wire signal_17505 ;
    wire signal_17506 ;
    wire signal_17507 ;
    wire signal_17508 ;
    wire signal_17509 ;
    wire signal_17510 ;
    wire signal_17511 ;
    wire signal_17512 ;
    wire signal_17513 ;
    wire signal_17514 ;
    wire signal_17515 ;
    wire signal_17516 ;
    wire signal_17517 ;
    wire signal_17518 ;
    wire signal_17519 ;
    wire signal_17520 ;
    wire signal_17521 ;
    wire signal_17522 ;
    wire signal_17523 ;
    wire signal_17524 ;
    wire signal_17525 ;
    wire signal_17526 ;
    wire signal_17527 ;
    wire signal_17528 ;
    wire signal_17529 ;
    wire signal_17530 ;
    wire signal_17531 ;
    wire signal_17532 ;
    wire signal_17533 ;
    wire signal_17534 ;
    wire signal_17535 ;
    wire signal_17536 ;
    wire signal_17537 ;
    wire signal_17538 ;
    wire signal_17539 ;
    wire signal_17540 ;
    wire signal_17541 ;
    wire signal_17542 ;
    wire signal_17543 ;
    wire signal_17544 ;
    wire signal_17545 ;
    wire signal_17546 ;
    wire signal_17547 ;
    wire signal_17548 ;
    wire signal_17549 ;
    wire signal_17550 ;
    wire signal_17551 ;
    wire signal_17552 ;
    wire signal_17553 ;
    wire signal_17554 ;
    wire signal_17555 ;
    wire signal_17556 ;
    wire signal_17557 ;
    wire signal_17558 ;
    wire signal_17559 ;
    wire signal_17560 ;
    wire signal_17561 ;
    wire signal_17562 ;
    wire signal_17563 ;
    wire signal_17564 ;
    wire signal_17565 ;
    wire signal_17566 ;
    wire signal_17567 ;
    wire signal_17568 ;
    wire signal_17569 ;
    wire signal_17570 ;
    wire signal_17571 ;
    wire signal_17572 ;
    wire signal_17573 ;
    wire signal_17574 ;
    wire signal_17575 ;
    wire signal_17576 ;
    wire signal_17577 ;
    wire signal_17578 ;
    wire signal_17579 ;
    wire signal_17580 ;
    wire signal_17581 ;
    wire signal_17582 ;
    wire signal_17583 ;
    wire signal_17584 ;
    wire signal_17585 ;
    wire signal_17586 ;
    wire signal_17587 ;
    wire signal_17588 ;
    wire signal_17589 ;
    wire signal_17590 ;
    wire signal_17591 ;
    wire signal_17592 ;
    wire signal_17593 ;
    wire signal_17594 ;
    wire signal_17595 ;
    wire signal_17596 ;
    wire signal_17597 ;
    wire signal_17598 ;
    wire signal_17599 ;
    wire signal_17600 ;
    wire signal_17601 ;
    wire signal_17602 ;
    wire signal_17603 ;
    wire signal_17604 ;
    wire signal_17605 ;
    wire signal_17606 ;
    wire signal_17607 ;
    wire signal_17608 ;
    wire signal_17609 ;
    wire signal_17610 ;
    wire signal_17611 ;
    wire signal_17612 ;
    wire signal_17613 ;
    wire signal_17614 ;
    wire signal_17615 ;
    wire signal_17616 ;
    wire signal_17617 ;
    wire signal_17618 ;
    wire signal_17619 ;
    wire signal_17620 ;
    wire signal_17621 ;
    wire signal_17622 ;
    wire signal_17623 ;
    wire signal_17624 ;
    wire signal_17625 ;
    wire signal_17626 ;
    wire signal_17627 ;
    wire signal_17628 ;
    wire signal_17629 ;
    wire signal_17630 ;
    wire signal_17631 ;
    wire signal_17632 ;
    wire signal_17633 ;
    wire signal_17634 ;
    wire signal_17635 ;
    wire signal_17636 ;
    wire signal_17637 ;
    wire signal_17638 ;
    wire signal_17639 ;
    wire signal_17640 ;
    wire signal_17641 ;
    wire signal_17642 ;
    wire signal_17643 ;
    wire signal_17644 ;
    wire signal_17645 ;
    wire signal_17646 ;
    wire signal_17647 ;
    wire signal_17648 ;
    wire signal_17649 ;
    wire signal_17650 ;
    wire signal_17651 ;
    wire signal_17652 ;
    wire signal_17653 ;
    wire signal_17654 ;
    wire signal_17655 ;
    wire signal_17656 ;
    wire signal_17657 ;
    wire signal_17658 ;
    wire signal_17659 ;
    wire signal_17660 ;
    wire signal_17661 ;
    wire signal_17662 ;
    wire signal_17663 ;
    wire signal_17664 ;
    wire signal_17665 ;
    wire signal_17666 ;
    wire signal_17667 ;
    wire signal_17668 ;
    wire signal_17669 ;
    wire signal_17670 ;
    wire signal_17671 ;
    wire signal_17672 ;
    wire signal_17673 ;
    wire signal_17674 ;
    wire signal_17675 ;
    wire signal_17676 ;
    wire signal_17677 ;
    wire signal_17678 ;
    wire signal_17679 ;
    wire signal_17680 ;
    wire signal_17681 ;
    wire signal_17682 ;
    wire signal_17683 ;
    wire signal_17684 ;
    wire signal_17685 ;
    wire signal_17686 ;
    wire signal_17687 ;
    wire signal_17688 ;
    wire signal_17689 ;
    wire signal_17690 ;
    wire signal_17691 ;
    wire signal_17692 ;
    wire signal_17693 ;
    wire signal_17694 ;
    wire signal_17695 ;
    wire signal_17696 ;
    wire signal_17697 ;
    wire signal_17698 ;
    wire signal_17699 ;
    wire signal_17700 ;
    wire signal_17701 ;
    wire signal_17702 ;
    wire signal_17703 ;
    wire signal_17704 ;
    wire signal_17705 ;
    wire signal_17706 ;
    wire signal_17707 ;
    wire signal_17708 ;
    wire signal_17709 ;
    wire signal_17710 ;
    wire signal_17711 ;
    wire signal_17712 ;
    wire signal_17713 ;
    wire signal_17714 ;
    wire signal_17715 ;
    wire signal_17716 ;
    wire signal_17717 ;
    wire signal_17718 ;
    wire signal_17719 ;
    wire signal_17720 ;
    wire signal_17721 ;
    wire signal_17722 ;
    wire signal_17723 ;
    wire signal_17724 ;
    wire signal_17725 ;
    wire signal_17726 ;
    wire signal_17727 ;
    wire signal_17728 ;
    wire signal_17729 ;
    wire signal_17730 ;
    wire signal_17731 ;
    wire signal_17732 ;
    wire signal_17733 ;
    wire signal_17734 ;
    wire signal_17735 ;
    wire signal_17736 ;
    wire signal_17737 ;
    wire signal_17738 ;
    wire signal_17739 ;
    wire signal_17740 ;
    wire signal_17741 ;
    wire signal_17742 ;
    wire signal_17743 ;
    wire signal_17744 ;
    wire signal_17745 ;
    wire signal_17746 ;
    wire signal_17747 ;
    wire signal_17748 ;
    wire signal_17749 ;
    wire signal_17750 ;
    wire signal_17751 ;
    wire signal_17752 ;
    wire signal_17753 ;
    wire signal_17754 ;
    wire signal_17755 ;
    wire signal_17756 ;
    wire signal_17757 ;
    wire signal_17758 ;
    wire signal_17759 ;
    wire signal_17760 ;
    wire signal_17761 ;
    wire signal_17762 ;
    wire signal_17763 ;
    wire signal_17764 ;
    wire signal_17765 ;
    wire signal_17766 ;
    wire signal_17767 ;
    wire signal_17768 ;
    wire signal_17769 ;
    wire signal_17770 ;
    wire signal_17771 ;
    wire signal_17772 ;
    wire signal_17773 ;
    wire signal_17774 ;
    wire signal_17775 ;
    wire signal_17776 ;
    wire signal_17777 ;
    wire signal_17778 ;
    wire signal_17779 ;
    wire signal_17780 ;
    wire signal_17781 ;
    wire signal_17782 ;
    wire signal_17783 ;
    wire signal_17784 ;
    wire signal_17785 ;
    wire signal_17786 ;
    wire signal_17787 ;
    wire signal_17788 ;
    wire signal_17789 ;
    wire signal_17790 ;
    wire signal_17791 ;
    wire signal_17792 ;
    wire signal_17793 ;
    wire signal_17794 ;
    wire signal_17795 ;
    wire signal_17796 ;
    wire signal_17797 ;
    wire signal_17798 ;
    wire signal_17799 ;
    wire signal_17800 ;
    wire signal_17801 ;
    wire signal_17802 ;
    wire signal_17803 ;
    wire signal_17804 ;
    wire signal_17805 ;
    wire signal_17806 ;
    wire signal_17807 ;
    wire signal_17808 ;
    wire signal_17809 ;
    wire signal_17810 ;
    wire signal_17811 ;
    wire signal_17812 ;
    wire signal_17813 ;
    wire signal_17814 ;
    wire signal_17815 ;
    wire signal_17816 ;
    wire signal_17817 ;
    wire signal_17818 ;
    wire signal_17819 ;
    wire signal_17820 ;
    wire signal_17821 ;
    wire signal_17822 ;
    wire signal_17823 ;
    wire signal_17824 ;
    wire signal_17825 ;
    wire signal_17826 ;
    wire signal_17827 ;
    wire signal_17828 ;
    wire signal_17829 ;
    wire signal_17830 ;
    wire signal_17831 ;
    wire signal_17832 ;
    wire signal_17833 ;
    wire signal_17834 ;
    wire signal_17835 ;
    wire signal_17836 ;
    wire signal_17837 ;
    wire signal_17838 ;
    wire signal_17839 ;
    wire signal_17840 ;
    wire signal_17841 ;
    wire signal_17842 ;
    wire signal_17843 ;
    wire signal_17844 ;
    wire signal_17845 ;
    wire signal_17846 ;
    wire signal_17847 ;
    wire signal_17848 ;
    wire signal_17849 ;
    wire signal_17850 ;
    wire signal_17851 ;
    wire signal_17852 ;
    wire signal_17853 ;
    wire signal_17854 ;
    wire signal_17855 ;
    wire signal_17856 ;
    wire signal_17857 ;
    wire signal_17858 ;
    wire signal_17859 ;
    wire signal_17860 ;
    wire signal_17861 ;
    wire signal_17862 ;
    wire signal_17863 ;
    wire signal_17864 ;
    wire signal_17865 ;
    wire signal_17866 ;
    wire signal_17867 ;
    wire signal_17868 ;
    wire signal_17869 ;
    wire signal_17870 ;
    wire signal_17871 ;
    wire signal_17872 ;
    wire signal_17873 ;
    wire signal_17874 ;
    wire signal_17875 ;
    wire signal_17876 ;
    wire signal_17877 ;
    wire signal_17878 ;
    wire signal_17879 ;
    wire signal_17880 ;
    wire signal_17881 ;
    wire signal_17882 ;
    wire signal_17883 ;
    wire signal_17884 ;
    wire signal_17885 ;
    wire signal_17886 ;
    wire signal_17887 ;
    wire signal_17888 ;
    wire signal_17889 ;
    wire signal_17890 ;
    wire signal_17891 ;
    wire signal_17892 ;
    wire signal_17893 ;
    wire signal_17894 ;
    wire signal_17895 ;
    wire signal_17896 ;
    wire signal_17897 ;
    wire signal_17898 ;
    wire signal_17899 ;
    wire signal_17900 ;
    wire signal_17901 ;
    wire signal_17902 ;
    wire signal_17903 ;
    wire signal_17904 ;
    wire signal_17905 ;
    wire signal_17906 ;
    wire signal_17907 ;
    wire signal_17908 ;
    wire signal_17909 ;
    wire signal_17910 ;
    wire signal_17911 ;
    wire signal_17912 ;
    wire signal_17913 ;
    wire signal_17914 ;
    wire signal_17915 ;
    wire signal_17916 ;
    wire signal_17917 ;
    wire signal_17918 ;
    wire signal_17919 ;
    wire signal_17920 ;
    wire signal_17921 ;
    wire signal_17922 ;
    wire signal_17923 ;
    wire signal_17924 ;
    wire signal_17925 ;
    wire signal_17926 ;
    wire signal_17927 ;
    wire signal_17928 ;
    wire signal_17929 ;
    wire signal_17930 ;
    wire signal_17931 ;
    wire signal_17932 ;
    wire signal_17933 ;
    wire signal_17934 ;
    wire signal_17935 ;
    wire signal_17936 ;
    wire signal_17937 ;
    wire signal_17938 ;
    wire signal_17939 ;
    wire signal_17940 ;
    wire signal_17941 ;
    wire signal_17942 ;
    wire signal_17943 ;
    wire signal_17944 ;
    wire signal_17945 ;
    wire signal_17946 ;
    wire signal_17947 ;
    wire signal_17948 ;
    wire signal_17949 ;
    wire signal_17950 ;
    wire signal_17951 ;
    wire signal_17952 ;
    wire signal_17953 ;
    wire signal_17954 ;
    wire signal_17955 ;
    wire signal_17956 ;
    wire signal_17957 ;
    wire signal_17958 ;
    wire signal_17959 ;
    wire signal_17960 ;
    wire signal_17961 ;
    wire signal_17962 ;
    wire signal_17963 ;
    wire signal_17964 ;
    wire signal_17965 ;
    wire signal_17966 ;
    wire signal_17967 ;
    wire signal_17968 ;
    wire signal_17969 ;
    wire signal_17970 ;
    wire signal_17971 ;
    wire signal_17972 ;
    wire signal_17973 ;
    wire signal_17974 ;
    wire signal_17975 ;
    wire signal_17976 ;
    wire signal_17977 ;
    wire signal_17978 ;
    wire signal_17979 ;
    wire signal_17980 ;
    wire signal_17981 ;
    wire signal_17982 ;
    wire signal_17983 ;
    wire signal_17984 ;
    wire signal_17985 ;
    wire signal_17986 ;
    wire signal_17987 ;
    wire signal_17988 ;
    wire signal_17989 ;
    wire signal_17990 ;
    wire signal_17991 ;
    wire signal_17992 ;
    wire signal_17993 ;
    wire signal_17994 ;
    wire signal_17995 ;
    wire signal_17996 ;
    wire signal_17997 ;
    wire signal_17998 ;
    wire signal_17999 ;
    wire signal_18000 ;
    wire signal_18001 ;
    wire signal_18002 ;
    wire signal_18003 ;
    wire signal_18004 ;
    wire signal_18005 ;
    wire signal_18006 ;
    wire signal_18007 ;
    wire signal_18008 ;
    wire signal_18009 ;
    wire signal_18010 ;
    wire signal_18011 ;
    wire signal_18012 ;
    wire signal_18013 ;
    wire signal_18014 ;
    wire signal_18015 ;
    wire signal_18016 ;
    wire signal_18017 ;
    wire signal_18018 ;
    wire signal_18019 ;
    wire signal_18020 ;
    wire signal_18021 ;
    wire signal_18022 ;
    wire signal_18023 ;
    wire signal_18024 ;
    wire signal_18025 ;
    wire signal_18026 ;
    wire signal_18027 ;
    wire signal_18028 ;
    wire signal_18029 ;
    wire signal_18030 ;
    wire signal_18031 ;
    wire signal_18032 ;
    wire signal_18033 ;
    wire signal_18034 ;
    wire signal_18035 ;
    wire signal_18036 ;
    wire signal_18037 ;
    wire signal_18038 ;
    wire signal_18039 ;
    wire signal_18040 ;
    wire signal_18041 ;
    wire signal_18042 ;
    wire signal_18043 ;
    wire signal_18044 ;
    wire signal_18045 ;
    wire signal_18046 ;
    wire signal_18047 ;
    wire signal_18048 ;
    wire signal_18049 ;
    wire signal_18050 ;
    wire signal_18051 ;
    wire signal_18052 ;
    wire signal_18053 ;
    wire signal_18054 ;
    wire signal_18055 ;
    wire signal_18056 ;
    wire signal_18057 ;
    wire signal_18058 ;
    wire signal_18059 ;
    wire signal_18060 ;
    wire signal_18061 ;
    wire signal_18062 ;
    wire signal_18063 ;
    wire signal_18064 ;
    wire signal_18065 ;
    wire signal_18066 ;
    wire signal_18067 ;
    wire signal_18068 ;
    wire signal_18069 ;
    wire signal_18070 ;
    wire signal_18071 ;
    wire signal_18072 ;
    wire signal_18073 ;
    wire signal_18074 ;
    wire signal_18075 ;
    wire signal_18076 ;
    wire signal_18077 ;
    wire signal_18078 ;
    wire signal_18079 ;
    wire signal_18080 ;
    wire signal_18081 ;
    wire signal_18082 ;
    wire signal_18083 ;
    wire signal_18084 ;
    wire signal_18085 ;
    wire signal_18086 ;
    wire signal_18087 ;
    wire signal_18088 ;
    wire signal_18089 ;
    wire signal_18090 ;
    wire signal_18091 ;
    wire signal_18092 ;
    wire signal_18093 ;
    wire signal_18094 ;
    wire signal_18095 ;
    wire signal_18096 ;
    wire signal_18097 ;
    wire signal_18098 ;
    wire signal_18099 ;
    wire signal_18100 ;
    wire signal_18101 ;
    wire signal_18102 ;
    wire signal_18103 ;
    wire signal_18104 ;
    wire signal_18105 ;
    wire signal_18106 ;
    wire signal_18107 ;
    wire signal_18108 ;
    wire signal_18109 ;
    wire signal_18110 ;
    wire signal_18111 ;
    wire signal_18112 ;
    wire signal_18113 ;
    wire signal_18114 ;
    wire signal_18115 ;
    wire signal_18116 ;
    wire signal_18117 ;
    wire signal_18118 ;
    wire signal_18119 ;
    wire signal_18120 ;
    wire signal_18121 ;
    wire signal_18122 ;
    wire signal_18123 ;
    wire signal_18124 ;
    wire signal_18125 ;
    wire signal_18126 ;
    wire signal_18127 ;
    wire signal_18128 ;
    wire signal_18129 ;
    wire signal_18130 ;
    wire signal_18131 ;
    wire signal_18132 ;
    wire signal_18133 ;
    wire signal_18134 ;
    wire signal_18135 ;
    wire signal_18136 ;
    wire signal_18137 ;
    wire signal_18138 ;
    wire signal_18139 ;
    wire signal_18140 ;
    wire signal_18141 ;
    wire signal_18142 ;
    wire signal_18143 ;
    wire signal_18144 ;
    wire signal_18145 ;
    wire signal_18146 ;
    wire signal_18147 ;
    wire signal_18148 ;
    wire signal_18149 ;
    wire signal_18150 ;
    wire signal_18151 ;
    wire signal_18152 ;
    wire signal_18153 ;
    wire signal_18154 ;
    wire signal_18155 ;
    wire signal_18156 ;
    wire signal_18157 ;
    wire signal_18158 ;
    wire signal_18159 ;
    wire signal_18160 ;
    wire signal_18161 ;
    wire signal_18162 ;
    wire signal_18163 ;
    wire signal_18164 ;
    wire signal_18165 ;
    wire signal_18166 ;
    wire signal_18167 ;
    wire signal_18168 ;
    wire signal_18169 ;
    wire signal_18170 ;
    wire signal_18171 ;
    wire signal_18172 ;
    wire signal_18173 ;
    wire signal_18174 ;
    wire signal_18175 ;
    wire signal_18176 ;
    wire signal_18177 ;
    wire signal_18178 ;
    wire signal_18179 ;
    wire signal_18180 ;
    wire signal_18181 ;
    wire signal_18182 ;
    wire signal_18183 ;
    wire signal_18184 ;
    wire signal_18185 ;
    wire signal_18186 ;
    wire signal_18187 ;
    wire signal_18188 ;
    wire signal_18189 ;
    wire signal_18190 ;
    wire signal_18191 ;
    wire signal_18192 ;
    wire signal_18193 ;
    wire signal_18194 ;
    wire signal_18195 ;
    wire signal_18196 ;
    wire signal_18197 ;
    wire signal_18198 ;
    wire signal_18199 ;
    wire signal_18200 ;
    wire signal_18201 ;
    wire signal_18202 ;
    wire signal_18203 ;
    wire signal_18204 ;
    wire signal_18205 ;
    wire signal_18206 ;
    wire signal_18207 ;
    wire signal_18208 ;
    wire signal_18209 ;
    wire signal_18210 ;
    wire signal_18211 ;
    wire signal_18212 ;
    wire signal_18213 ;
    wire signal_18214 ;
    wire signal_18215 ;
    wire signal_18216 ;
    wire signal_18217 ;
    wire signal_18218 ;
    wire signal_18219 ;
    wire signal_18220 ;
    wire signal_18221 ;
    wire signal_18222 ;
    wire signal_18223 ;
    wire signal_18224 ;
    wire signal_18225 ;
    wire signal_18226 ;
    wire signal_18227 ;
    wire signal_18228 ;
    wire signal_18229 ;
    wire signal_18230 ;
    wire signal_18231 ;
    wire signal_18232 ;
    wire signal_18233 ;
    wire signal_18234 ;
    wire signal_18235 ;
    wire signal_18236 ;
    wire signal_18237 ;
    wire signal_18238 ;
    wire signal_18239 ;
    wire signal_18240 ;
    wire signal_18241 ;
    wire signal_18242 ;
    wire signal_18243 ;
    wire signal_18244 ;
    wire signal_18245 ;
    wire signal_18246 ;
    wire signal_18247 ;
    wire signal_18248 ;
    wire signal_18249 ;
    wire signal_18250 ;
    wire signal_18251 ;
    wire signal_18252 ;
    wire signal_18253 ;
    wire signal_18254 ;
    wire signal_18255 ;
    wire signal_18256 ;
    wire signal_18257 ;
    wire signal_18258 ;
    wire signal_18259 ;
    wire signal_18260 ;
    wire signal_18261 ;
    wire signal_18262 ;
    wire signal_18263 ;
    wire signal_18264 ;
    wire signal_18265 ;
    wire signal_18266 ;
    wire signal_18267 ;
    wire signal_18268 ;
    wire signal_18269 ;
    wire signal_18270 ;
    wire signal_18271 ;
    wire signal_18272 ;
    wire signal_18273 ;
    wire signal_18274 ;
    wire signal_18275 ;
    wire signal_18276 ;
    wire signal_18277 ;
    wire signal_18278 ;
    wire signal_18279 ;
    wire signal_18280 ;
    wire signal_18281 ;
    wire signal_18282 ;
    wire signal_18283 ;
    wire signal_18284 ;
    wire signal_18285 ;
    wire signal_18286 ;
    wire signal_18287 ;
    wire signal_18288 ;
    wire signal_18289 ;
    wire signal_18290 ;
    wire signal_18291 ;
    wire signal_18292 ;
    wire signal_18293 ;
    wire signal_18294 ;
    wire signal_18295 ;
    wire signal_18296 ;
    wire signal_18297 ;
    wire signal_18298 ;
    wire signal_18299 ;
    wire signal_18300 ;
    wire signal_18301 ;
    wire signal_18302 ;
    wire signal_18303 ;
    wire signal_18304 ;
    wire signal_18305 ;
    wire signal_18306 ;
    wire signal_18307 ;
    wire signal_18308 ;
    wire signal_18309 ;
    wire signal_18310 ;
    wire signal_18311 ;
    wire signal_18312 ;
    wire signal_18313 ;
    wire signal_18314 ;
    wire signal_18315 ;
    wire signal_18316 ;
    wire signal_18317 ;
    wire signal_18318 ;
    wire signal_18319 ;
    wire signal_18320 ;
    wire signal_18321 ;
    wire signal_18322 ;
    wire signal_18323 ;
    wire signal_18324 ;
    wire signal_18325 ;
    wire signal_18326 ;
    wire signal_18327 ;
    wire signal_18328 ;
    wire signal_18329 ;
    wire signal_18330 ;
    wire signal_18331 ;
    wire signal_18332 ;
    wire signal_18333 ;
    wire signal_18334 ;
    wire signal_18335 ;
    wire signal_18336 ;
    wire signal_18337 ;
    wire signal_18338 ;
    wire signal_18339 ;
    wire signal_18340 ;
    wire signal_18341 ;
    wire signal_18342 ;
    wire signal_18343 ;
    wire signal_18344 ;
    wire signal_18345 ;
    wire signal_18346 ;
    wire signal_18347 ;
    wire signal_18348 ;
    wire signal_18349 ;
    wire signal_18350 ;
    wire signal_18351 ;
    wire signal_18352 ;
    wire signal_18353 ;
    wire signal_18354 ;
    wire signal_18355 ;
    wire signal_18356 ;
    wire signal_18357 ;
    wire signal_18358 ;
    wire signal_18359 ;
    wire signal_18360 ;
    wire signal_18361 ;
    wire signal_18362 ;
    wire signal_18363 ;
    wire signal_18364 ;
    wire signal_18365 ;
    wire signal_18366 ;
    wire signal_18367 ;
    wire signal_18368 ;
    wire signal_18369 ;
    wire signal_18370 ;
    wire signal_18371 ;
    wire signal_18372 ;
    wire signal_18373 ;
    wire signal_18374 ;
    wire signal_18375 ;
    wire signal_18376 ;
    wire signal_18377 ;
    wire signal_18378 ;
    wire signal_18379 ;
    wire signal_18380 ;
    wire signal_18381 ;
    wire signal_18382 ;
    wire signal_18383 ;
    wire signal_18384 ;
    wire signal_18385 ;
    wire signal_18386 ;
    wire signal_18387 ;
    wire signal_18388 ;
    wire signal_18389 ;
    wire signal_18390 ;
    wire signal_18391 ;
    wire signal_18392 ;
    wire signal_18393 ;
    wire signal_18394 ;
    wire signal_18395 ;
    wire signal_18396 ;
    wire signal_18397 ;
    wire signal_18398 ;
    wire signal_18399 ;
    wire signal_18400 ;
    wire signal_18401 ;
    wire signal_18402 ;
    wire signal_18403 ;
    wire signal_18404 ;
    wire signal_18405 ;
    wire signal_18406 ;
    wire signal_18407 ;
    wire signal_18408 ;
    wire signal_18409 ;
    wire signal_18410 ;
    wire signal_18411 ;
    wire signal_18412 ;
    wire signal_18413 ;
    wire signal_18414 ;
    wire signal_18415 ;
    wire signal_18416 ;
    wire signal_18417 ;
    wire signal_18418 ;
    wire signal_18419 ;
    wire signal_18420 ;
    wire signal_18421 ;
    wire signal_18422 ;
    wire signal_18423 ;
    wire signal_18424 ;
    wire signal_18425 ;
    wire signal_18426 ;
    wire signal_18427 ;
    wire signal_18428 ;
    wire signal_18429 ;
    wire signal_18430 ;
    wire signal_18431 ;
    wire signal_18432 ;
    wire signal_18433 ;
    wire signal_18434 ;
    wire signal_18435 ;
    wire signal_18436 ;
    wire signal_18437 ;
    wire signal_18438 ;
    wire signal_18439 ;
    wire signal_18440 ;
    wire signal_18441 ;
    wire signal_18442 ;
    wire signal_18443 ;
    wire signal_18444 ;
    wire signal_18445 ;
    wire signal_18446 ;
    wire signal_18447 ;
    wire signal_18448 ;
    wire signal_18449 ;
    wire signal_18450 ;
    wire signal_18451 ;
    wire signal_18452 ;
    wire signal_18453 ;
    wire signal_18454 ;
    wire signal_18455 ;
    wire signal_18456 ;
    wire signal_18457 ;
    wire signal_18458 ;
    wire signal_18459 ;
    wire signal_18460 ;
    wire signal_18461 ;
    wire signal_18462 ;
    wire signal_18463 ;
    wire signal_18464 ;
    wire signal_18465 ;
    wire signal_18466 ;
    wire signal_18467 ;
    wire signal_18468 ;
    wire signal_18469 ;
    wire signal_18470 ;
    wire signal_18471 ;
    wire signal_18472 ;
    wire signal_18473 ;
    wire signal_18474 ;
    wire signal_18475 ;
    wire signal_18476 ;
    wire signal_18477 ;
    wire signal_18478 ;
    wire signal_18479 ;
    wire signal_18480 ;
    wire signal_18481 ;
    wire signal_18482 ;
    wire signal_18483 ;
    wire signal_18484 ;
    wire signal_18485 ;
    wire signal_18486 ;
    wire signal_18487 ;
    wire signal_18488 ;
    wire signal_18489 ;
    wire signal_18490 ;
    wire signal_18491 ;
    wire signal_18492 ;
    wire signal_18493 ;
    wire signal_18494 ;
    wire signal_18495 ;
    wire signal_18496 ;
    wire signal_18497 ;
    wire signal_18498 ;
    wire signal_18499 ;
    wire signal_18500 ;
    wire signal_18501 ;
    wire signal_18502 ;
    wire signal_18503 ;
    wire signal_18504 ;
    wire signal_18505 ;
    wire signal_18506 ;
    wire signal_18507 ;
    wire signal_18508 ;
    wire signal_18509 ;
    wire signal_18510 ;
    wire signal_18511 ;
    wire signal_18512 ;
    wire signal_18513 ;
    wire signal_18514 ;
    wire signal_18515 ;
    wire signal_18516 ;
    wire signal_18517 ;
    wire signal_18518 ;
    wire signal_18519 ;
    wire signal_18520 ;
    wire signal_18521 ;
    wire signal_18522 ;
    wire signal_18523 ;
    wire signal_18524 ;
    wire signal_18525 ;
    wire signal_18526 ;
    wire signal_18527 ;
    wire signal_18528 ;
    wire signal_18529 ;
    wire signal_18530 ;
    wire signal_18531 ;
    wire signal_18532 ;
    wire signal_18533 ;
    wire signal_18534 ;
    wire signal_18535 ;
    wire signal_18536 ;
    wire signal_18537 ;
    wire signal_18538 ;
    wire signal_18539 ;
    wire signal_18540 ;
    wire signal_18541 ;
    wire signal_18542 ;
    wire signal_18543 ;
    wire signal_18544 ;
    wire signal_18545 ;
    wire signal_18546 ;
    wire signal_18547 ;
    wire signal_18548 ;
    wire signal_18549 ;
    wire signal_18550 ;
    wire signal_18551 ;
    wire signal_18552 ;
    wire signal_18553 ;
    wire signal_18554 ;
    wire signal_18555 ;
    wire signal_18556 ;
    wire signal_18557 ;
    wire signal_18558 ;
    wire signal_18559 ;
    wire signal_18560 ;
    wire signal_18561 ;
    wire signal_18562 ;
    wire signal_18563 ;
    wire signal_18564 ;
    wire signal_18565 ;
    wire signal_18566 ;
    wire signal_18567 ;
    wire signal_18568 ;
    wire signal_18569 ;
    wire signal_18570 ;
    wire signal_18571 ;
    wire signal_18572 ;
    wire signal_18573 ;
    wire signal_18574 ;
    wire signal_18575 ;
    wire signal_18576 ;
    wire signal_18577 ;
    wire signal_18578 ;
    wire signal_18579 ;
    wire signal_18580 ;
    wire signal_18581 ;
    wire signal_18582 ;
    wire signal_18583 ;
    wire signal_18584 ;
    wire signal_18585 ;
    wire signal_18586 ;
    wire signal_18587 ;
    wire signal_18588 ;
    wire signal_18589 ;
    wire signal_18590 ;
    wire signal_18591 ;
    wire signal_18592 ;
    wire signal_18593 ;
    wire signal_18594 ;
    wire signal_18595 ;
    wire signal_18596 ;
    wire signal_18597 ;
    wire signal_18598 ;
    wire signal_18599 ;
    wire signal_18600 ;
    wire signal_18601 ;
    wire signal_18602 ;
    wire signal_18603 ;
    wire signal_18604 ;
    wire signal_18605 ;
    wire signal_18606 ;
    wire signal_18607 ;
    wire signal_18608 ;
    wire signal_18609 ;
    wire signal_18610 ;
    wire signal_18611 ;
    wire signal_18612 ;
    wire signal_18613 ;
    wire signal_18614 ;
    wire signal_18615 ;
    wire signal_18616 ;
    wire signal_18617 ;
    wire signal_18618 ;
    wire signal_18619 ;
    wire signal_18620 ;
    wire signal_18621 ;
    wire signal_18622 ;
    wire signal_18623 ;
    wire signal_18624 ;
    wire signal_18625 ;
    wire signal_18626 ;
    wire signal_18627 ;
    wire signal_18628 ;
    wire signal_18629 ;
    wire signal_18630 ;
    wire signal_18631 ;
    wire signal_18632 ;
    wire signal_18633 ;
    wire signal_18634 ;
    wire signal_18635 ;
    wire signal_18636 ;
    wire signal_18637 ;
    wire signal_18638 ;
    wire signal_18639 ;
    wire signal_18640 ;
    wire signal_18641 ;
    wire signal_18642 ;
    wire signal_18643 ;
    wire signal_18644 ;
    wire signal_18645 ;
    wire signal_18646 ;
    wire signal_18647 ;
    wire signal_18648 ;
    wire signal_18649 ;
    wire signal_18650 ;
    wire signal_18651 ;
    wire signal_18652 ;
    wire signal_18653 ;
    wire signal_18654 ;
    wire signal_18655 ;
    wire signal_18656 ;
    wire signal_18657 ;
    wire signal_18658 ;
    wire signal_18659 ;
    wire signal_18660 ;
    wire signal_18661 ;
    wire signal_18662 ;
    wire signal_18663 ;
    wire signal_18664 ;
    wire signal_18665 ;
    wire signal_18666 ;
    wire signal_18667 ;
    wire signal_18668 ;
    wire signal_18669 ;
    wire signal_18670 ;
    wire signal_18671 ;
    wire signal_18672 ;
    wire signal_18673 ;
    wire signal_18674 ;
    wire signal_18675 ;
    wire signal_18676 ;
    wire signal_18677 ;
    wire signal_18678 ;
    wire signal_18679 ;
    wire signal_18680 ;
    wire signal_18681 ;
    wire signal_18682 ;
    wire signal_18683 ;
    wire signal_18684 ;
    wire signal_18685 ;
    wire signal_18686 ;
    wire signal_18687 ;
    wire signal_18688 ;
    wire signal_18689 ;
    wire signal_18690 ;
    wire signal_18691 ;
    wire signal_18692 ;
    wire signal_18693 ;
    wire signal_18694 ;
    wire signal_18695 ;
    wire signal_18696 ;
    wire signal_18697 ;
    wire signal_18698 ;
    wire signal_18699 ;
    wire signal_18700 ;
    wire signal_18701 ;
    wire signal_18702 ;
    wire signal_18703 ;
    wire signal_18704 ;
    wire signal_18705 ;
    wire signal_18706 ;
    wire signal_18707 ;
    wire signal_18708 ;
    wire signal_18709 ;
    wire signal_18710 ;
    wire signal_18711 ;
    wire signal_18712 ;
    wire signal_18713 ;
    wire signal_18714 ;
    wire signal_18715 ;
    wire signal_18716 ;
    wire signal_18717 ;
    wire signal_18718 ;
    wire signal_18719 ;
    wire signal_18720 ;
    wire signal_18721 ;
    wire signal_18722 ;
    wire signal_18723 ;
    wire signal_18724 ;
    wire signal_18725 ;
    wire signal_18726 ;
    wire signal_18727 ;
    wire signal_18728 ;
    wire signal_18729 ;
    wire signal_18730 ;
    wire signal_18731 ;
    wire signal_18732 ;
    wire signal_18733 ;
    wire signal_18734 ;
    wire signal_18735 ;
    wire signal_18736 ;
    wire signal_18737 ;
    wire signal_18738 ;
    wire signal_18739 ;
    wire signal_18740 ;
    wire signal_18741 ;
    wire signal_18742 ;
    wire signal_18743 ;
    wire signal_18744 ;
    wire signal_18745 ;
    wire signal_18746 ;
    wire signal_18747 ;
    wire signal_18748 ;
    wire signal_18749 ;
    wire signal_18750 ;
    wire signal_18751 ;
    wire signal_18752 ;
    wire signal_18753 ;
    wire signal_18754 ;
    wire signal_18755 ;
    wire signal_18756 ;
    wire signal_18757 ;
    wire signal_18758 ;
    wire signal_18759 ;
    wire signal_18760 ;
    wire signal_18761 ;
    wire signal_18762 ;
    wire signal_18763 ;
    wire signal_18764 ;
    wire signal_18765 ;
    wire signal_18766 ;
    wire signal_18767 ;
    wire signal_18768 ;
    wire signal_18769 ;
    wire signal_18770 ;
    wire signal_18771 ;
    wire signal_18772 ;
    wire signal_18773 ;
    wire signal_18774 ;
    wire signal_18775 ;
    wire signal_18776 ;
    wire signal_18777 ;
    wire signal_18778 ;
    wire signal_18779 ;
    wire signal_18780 ;
    wire signal_18781 ;
    wire signal_18782 ;
    wire signal_18783 ;
    wire signal_18784 ;
    wire signal_18785 ;
    wire signal_18786 ;
    wire signal_18787 ;
    wire signal_18788 ;
    wire signal_18789 ;
    wire signal_18790 ;
    wire signal_18791 ;
    wire signal_18792 ;
    wire signal_18793 ;
    wire signal_18794 ;
    wire signal_18795 ;
    wire signal_18796 ;
    wire signal_18797 ;
    wire signal_18798 ;
    wire signal_18799 ;
    wire signal_18800 ;
    wire signal_18801 ;
    wire signal_18802 ;
    wire signal_18803 ;
    wire signal_18804 ;
    wire signal_18805 ;
    wire signal_18806 ;
    wire signal_18807 ;
    wire signal_18808 ;
    wire signal_18809 ;
    wire signal_18810 ;
    wire signal_18811 ;
    wire signal_18812 ;
    wire signal_18813 ;
    wire signal_18814 ;
    wire signal_18815 ;
    wire signal_18816 ;
    wire signal_18817 ;
    wire signal_18818 ;
    wire signal_18819 ;
    wire signal_18820 ;
    wire signal_18821 ;
    wire signal_18822 ;
    wire signal_18823 ;
    wire signal_18824 ;
    wire signal_18825 ;
    wire signal_18826 ;
    wire signal_18827 ;
    wire signal_18828 ;
    wire signal_18829 ;
    wire signal_18830 ;
    wire signal_18831 ;
    wire signal_18832 ;
    wire signal_18833 ;
    wire signal_18834 ;
    wire signal_18835 ;
    wire signal_18836 ;
    wire signal_18837 ;
    wire signal_18838 ;
    wire signal_18839 ;
    wire signal_18840 ;
    wire signal_18841 ;
    wire signal_18842 ;
    wire signal_18843 ;
    wire signal_18844 ;
    wire signal_18845 ;
    wire signal_18846 ;
    wire signal_18847 ;
    wire signal_18848 ;
    wire signal_18849 ;
    wire signal_18850 ;
    wire signal_18851 ;
    wire signal_18852 ;
    wire signal_18853 ;
    wire signal_18854 ;
    wire signal_18855 ;
    wire signal_18856 ;
    wire signal_18857 ;
    wire signal_18858 ;
    wire signal_18859 ;
    wire signal_18860 ;
    wire signal_18861 ;
    wire signal_18862 ;
    wire signal_18863 ;
    wire signal_18864 ;
    wire signal_18865 ;
    wire signal_18866 ;
    wire signal_18867 ;
    wire signal_18868 ;
    wire signal_18869 ;
    wire signal_18870 ;
    wire signal_18871 ;
    wire signal_18872 ;
    wire signal_18873 ;
    wire signal_18874 ;
    wire signal_18875 ;
    wire signal_18876 ;
    wire signal_18877 ;
    wire signal_18878 ;
    wire signal_18879 ;
    wire signal_18880 ;
    wire signal_18881 ;
    wire signal_18882 ;
    wire signal_18883 ;
    wire signal_18884 ;
    wire signal_18885 ;
    wire signal_18886 ;
    wire signal_18887 ;
    wire signal_18888 ;
    wire signal_18889 ;
    wire signal_18890 ;
    wire signal_18891 ;
    wire signal_18892 ;
    wire signal_18893 ;
    wire signal_18894 ;
    wire signal_18895 ;
    wire signal_18896 ;
    wire signal_18897 ;
    wire signal_18898 ;
    wire signal_18899 ;
    wire signal_18900 ;
    wire signal_18901 ;
    wire signal_18902 ;
    wire signal_18903 ;
    wire signal_18904 ;
    wire signal_18905 ;
    wire signal_18906 ;
    wire signal_18907 ;
    wire signal_18908 ;
    wire signal_18909 ;
    wire signal_18910 ;
    wire signal_18911 ;
    wire signal_18912 ;
    wire signal_18913 ;
    wire signal_18914 ;
    wire signal_18915 ;
    wire signal_18916 ;
    wire signal_18917 ;
    wire signal_18918 ;
    wire signal_18919 ;
    wire signal_18920 ;
    wire signal_18921 ;
    wire signal_18922 ;
    wire signal_18923 ;
    wire signal_18924 ;
    wire signal_18925 ;
    wire signal_18926 ;
    wire signal_18927 ;
    wire signal_18928 ;
    wire signal_18929 ;
    wire signal_18930 ;
    wire signal_18931 ;
    wire signal_18932 ;
    wire signal_18933 ;
    wire signal_18934 ;
    wire signal_18935 ;
    wire signal_18936 ;
    wire signal_18937 ;
    wire signal_18938 ;
    wire signal_18939 ;
    wire signal_18940 ;
    wire signal_18941 ;
    wire signal_18942 ;
    wire signal_18943 ;
    wire signal_18944 ;
    wire signal_18945 ;
    wire signal_18946 ;
    wire signal_18947 ;
    wire signal_18948 ;
    wire signal_18949 ;
    wire signal_18950 ;
    wire signal_18951 ;
    wire signal_18952 ;
    wire signal_18953 ;
    wire signal_18954 ;
    wire signal_18955 ;
    wire signal_18956 ;
    wire signal_18957 ;
    wire signal_18958 ;
    wire signal_18959 ;
    wire signal_18960 ;
    wire signal_18961 ;
    wire signal_18962 ;
    wire signal_18963 ;
    wire signal_18964 ;
    wire signal_18965 ;
    wire signal_18966 ;
    wire signal_18967 ;
    wire signal_18968 ;
    wire signal_18969 ;
    wire signal_18970 ;
    wire signal_18971 ;
    wire signal_18972 ;
    wire signal_18973 ;
    wire signal_18974 ;
    wire signal_18975 ;
    wire signal_18976 ;
    wire signal_18977 ;
    wire signal_18978 ;
    wire signal_18979 ;
    wire signal_18980 ;
    wire signal_18981 ;
    wire signal_18982 ;
    wire signal_18983 ;
    wire signal_18984 ;
    wire signal_18985 ;
    wire signal_18986 ;
    wire signal_18987 ;
    wire signal_18988 ;
    wire signal_18989 ;
    wire signal_18990 ;
    wire signal_18991 ;
    wire signal_18992 ;
    wire signal_18993 ;
    wire signal_18994 ;
    wire signal_18995 ;
    wire signal_18996 ;
    wire signal_18997 ;
    wire signal_18998 ;
    wire signal_18999 ;
    wire signal_19000 ;
    wire signal_19001 ;
    wire signal_19002 ;
    wire signal_19003 ;
    wire signal_19004 ;
    wire signal_19005 ;
    wire signal_19006 ;
    wire signal_19007 ;
    wire signal_19008 ;
    wire signal_19009 ;
    wire signal_19010 ;
    wire signal_19011 ;
    wire signal_19012 ;
    wire signal_19013 ;
    wire signal_19014 ;
    wire signal_19015 ;
    wire signal_19016 ;
    wire signal_19017 ;
    wire signal_19018 ;
    wire signal_19019 ;
    wire signal_19020 ;
    wire signal_19021 ;
    wire signal_19022 ;
    wire signal_19023 ;
    wire signal_19024 ;
    wire signal_19025 ;
    wire signal_19026 ;
    wire signal_19027 ;
    wire signal_19028 ;
    wire signal_19029 ;
    wire signal_19030 ;
    wire signal_19031 ;
    wire signal_19032 ;
    wire signal_19033 ;
    wire signal_19034 ;
    wire signal_19035 ;
    wire signal_19036 ;
    wire signal_19037 ;
    wire signal_19038 ;
    wire signal_19039 ;
    wire signal_19040 ;
    wire signal_19041 ;
    wire signal_19042 ;
    wire signal_19043 ;
    wire signal_19044 ;
    wire signal_19045 ;
    wire signal_19046 ;
    wire signal_19047 ;
    wire signal_19048 ;
    wire signal_19049 ;
    wire signal_19050 ;
    wire signal_19051 ;
    wire signal_19052 ;
    wire signal_19053 ;
    wire signal_19054 ;
    wire signal_19055 ;
    wire signal_19056 ;
    wire signal_19057 ;
    wire signal_19058 ;
    wire signal_19059 ;
    wire signal_19060 ;
    wire signal_19061 ;
    wire signal_19062 ;
    wire signal_19063 ;
    wire signal_19064 ;
    wire signal_19065 ;
    wire signal_19066 ;
    wire signal_19067 ;
    wire signal_19068 ;
    wire signal_19069 ;
    wire signal_19070 ;
    wire signal_19071 ;
    wire signal_19072 ;
    wire signal_19073 ;
    wire signal_19074 ;
    wire signal_19075 ;
    wire signal_19076 ;
    wire signal_19077 ;
    wire signal_19078 ;
    wire signal_19079 ;
    wire signal_19080 ;
    wire signal_19081 ;
    wire signal_19082 ;
    wire signal_19083 ;
    wire signal_19084 ;
    wire signal_19085 ;
    wire signal_19086 ;
    wire signal_19087 ;
    wire signal_19088 ;
    wire signal_19089 ;
    wire signal_19090 ;
    wire signal_19091 ;
    wire signal_19092 ;
    wire signal_19093 ;
    wire signal_19094 ;
    wire signal_19095 ;
    wire signal_19096 ;
    wire signal_19097 ;
    wire signal_19098 ;
    wire signal_19099 ;
    wire signal_19100 ;
    wire signal_19101 ;
    wire signal_19102 ;
    wire signal_19103 ;
    wire signal_19104 ;
    wire signal_19105 ;
    wire signal_19106 ;
    wire signal_19107 ;
    wire signal_19108 ;
    wire signal_19109 ;
    wire signal_19110 ;
    wire signal_19111 ;
    wire signal_19112 ;
    wire signal_19113 ;
    wire signal_19114 ;
    wire signal_19115 ;
    wire signal_19116 ;
    wire signal_19117 ;
    wire signal_19118 ;
    wire signal_19119 ;
    wire signal_19120 ;
    wire signal_19121 ;
    wire signal_19122 ;
    wire signal_19123 ;
    wire signal_19124 ;
    wire signal_19125 ;
    wire signal_19126 ;
    wire signal_19127 ;
    wire signal_19128 ;
    wire signal_19129 ;
    wire signal_19130 ;
    wire signal_19131 ;
    wire signal_19132 ;
    wire signal_19133 ;
    wire signal_19134 ;
    wire signal_19135 ;
    wire signal_19136 ;
    wire signal_19137 ;
    wire signal_19138 ;
    wire signal_19139 ;
    wire signal_19140 ;
    wire signal_19141 ;
    wire signal_19142 ;
    wire signal_19143 ;
    wire signal_19144 ;
    wire signal_19145 ;
    wire signal_19146 ;
    wire signal_19147 ;
    wire signal_19148 ;
    wire signal_19149 ;
    wire signal_19150 ;
    wire signal_19151 ;
    wire signal_19152 ;
    wire signal_19153 ;
    wire signal_19154 ;
    wire signal_19155 ;
    wire signal_19156 ;
    wire signal_19157 ;
    wire signal_19158 ;
    wire signal_19159 ;
    wire signal_19160 ;
    wire signal_19161 ;
    wire signal_19162 ;
    wire signal_19163 ;
    wire signal_19164 ;
    wire signal_19165 ;
    wire signal_19166 ;
    wire signal_19167 ;
    wire signal_19168 ;
    wire signal_19169 ;
    wire signal_19170 ;
    wire signal_19171 ;
    wire signal_19172 ;
    wire signal_19173 ;
    wire signal_19174 ;
    wire signal_19175 ;
    wire signal_19176 ;
    wire signal_19177 ;
    wire signal_19178 ;
    wire signal_19179 ;
    wire signal_19180 ;
    wire signal_19181 ;
    wire signal_19182 ;
    wire signal_19183 ;
    wire signal_19184 ;
    wire signal_19185 ;
    wire signal_19186 ;
    wire signal_19187 ;
    wire signal_19188 ;
    wire signal_19189 ;
    wire signal_19190 ;
    wire signal_19191 ;
    wire signal_19192 ;
    wire signal_19193 ;
    wire signal_19194 ;
    wire signal_19195 ;
    wire signal_19196 ;
    wire signal_19197 ;
    wire signal_19198 ;
    wire signal_19199 ;
    wire signal_19200 ;
    wire signal_19201 ;
    wire signal_19202 ;
    wire signal_19203 ;
    wire signal_19204 ;
    wire signal_19205 ;
    wire signal_19206 ;
    wire signal_19207 ;
    wire signal_19208 ;
    wire signal_19209 ;
    wire signal_19210 ;
    wire signal_19211 ;
    wire signal_19212 ;
    wire signal_19213 ;
    wire signal_19214 ;
    wire signal_19215 ;
    wire signal_19216 ;
    wire signal_19217 ;
    wire signal_19218 ;
    wire signal_19219 ;
    wire signal_19220 ;
    wire signal_19221 ;
    wire signal_19222 ;
    wire signal_19223 ;
    wire signal_19224 ;
    wire signal_19225 ;
    wire signal_19226 ;
    wire signal_19227 ;
    wire signal_19228 ;
    wire signal_19229 ;
    wire signal_19230 ;
    wire signal_19231 ;
    wire signal_19232 ;
    wire signal_19233 ;
    wire signal_19234 ;
    wire signal_19235 ;
    wire signal_19236 ;
    wire signal_19237 ;
    wire signal_19238 ;
    wire signal_19239 ;
    wire signal_19240 ;
    wire signal_19241 ;
    wire signal_19242 ;
    wire signal_19243 ;
    wire signal_19244 ;
    wire signal_19245 ;
    wire signal_19246 ;
    wire signal_19247 ;
    wire signal_19248 ;
    wire signal_19249 ;
    wire signal_19250 ;
    wire signal_19251 ;
    wire signal_19252 ;
    wire signal_19253 ;
    wire signal_19254 ;
    wire signal_19255 ;
    wire signal_19256 ;
    wire signal_19257 ;
    wire signal_19258 ;
    wire signal_19259 ;
    wire signal_19260 ;
    wire signal_19261 ;
    wire signal_19262 ;
    wire signal_19263 ;
    wire signal_19264 ;
    wire signal_19265 ;
    wire signal_19266 ;
    wire signal_19267 ;
    wire signal_19268 ;
    wire signal_19269 ;
    wire signal_19270 ;
    wire signal_19271 ;
    wire signal_19272 ;
    wire signal_19273 ;
    wire signal_19274 ;
    wire signal_19275 ;
    wire signal_19276 ;
    wire signal_19277 ;
    wire signal_19278 ;
    wire signal_19279 ;
    wire signal_19280 ;
    wire signal_19281 ;
    wire signal_19282 ;
    wire signal_19283 ;
    wire signal_19284 ;
    wire signal_19285 ;
    wire signal_19286 ;
    wire signal_19287 ;
    wire signal_19288 ;
    wire signal_19289 ;
    wire signal_19290 ;
    wire signal_19291 ;
    wire signal_19292 ;
    wire signal_19293 ;
    wire signal_19294 ;
    wire signal_19295 ;
    wire signal_19296 ;
    wire signal_19297 ;
    wire signal_19298 ;
    wire signal_19299 ;
    wire signal_19300 ;
    wire signal_19301 ;
    wire signal_19302 ;
    wire signal_19303 ;
    wire signal_19304 ;
    wire signal_19305 ;
    wire signal_19306 ;
    wire signal_19307 ;
    wire signal_19308 ;
    wire signal_19309 ;
    wire signal_19310 ;
    wire signal_19311 ;
    wire signal_19312 ;
    wire signal_19313 ;
    wire signal_19314 ;
    wire signal_19315 ;
    wire signal_19316 ;
    wire signal_19317 ;
    wire signal_19318 ;
    wire signal_19319 ;
    wire signal_19320 ;
    wire signal_19321 ;
    wire signal_19322 ;
    wire signal_19323 ;
    wire signal_19324 ;
    wire signal_19325 ;
    wire signal_19326 ;
    wire signal_19327 ;
    wire signal_19328 ;
    wire signal_19329 ;
    wire signal_19330 ;
    wire signal_19331 ;
    wire signal_19332 ;
    wire signal_19333 ;
    wire signal_19334 ;
    wire signal_19335 ;
    wire signal_19336 ;
    wire signal_19337 ;
    wire signal_19338 ;
    wire signal_19339 ;
    wire signal_19340 ;
    wire signal_19341 ;
    wire signal_19342 ;
    wire signal_19343 ;
    wire signal_19344 ;
    wire signal_19345 ;
    wire signal_19346 ;
    wire signal_19347 ;
    wire signal_19348 ;
    wire signal_19349 ;
    wire signal_19350 ;
    wire signal_19351 ;
    wire signal_19352 ;
    wire signal_19353 ;
    wire signal_19354 ;
    wire signal_19355 ;
    wire signal_19356 ;
    wire signal_19357 ;
    wire signal_19358 ;
    wire signal_19359 ;
    wire signal_19360 ;
    wire signal_19361 ;
    wire signal_19362 ;
    wire signal_19363 ;
    wire signal_19364 ;
    wire signal_19365 ;
    wire signal_19366 ;
    wire signal_19367 ;
    wire signal_19368 ;
    wire signal_19369 ;
    wire signal_19370 ;
    wire signal_19371 ;
    wire signal_19372 ;
    wire signal_19373 ;
    wire signal_19374 ;
    wire signal_19375 ;
    wire signal_19376 ;
    wire signal_19377 ;
    wire signal_19378 ;
    wire signal_19379 ;
    wire signal_19380 ;
    wire signal_19381 ;
    wire signal_19382 ;
    wire signal_19383 ;
    wire signal_19384 ;
    wire signal_19385 ;
    wire signal_19386 ;
    wire signal_19387 ;
    wire signal_19388 ;
    wire signal_19389 ;
    wire signal_19390 ;
    wire signal_19391 ;
    wire signal_19392 ;
    wire signal_19393 ;
    wire signal_19394 ;
    wire signal_19395 ;
    wire signal_19396 ;
    wire signal_19397 ;
    wire signal_19398 ;
    wire signal_19399 ;
    wire signal_19400 ;
    wire signal_19401 ;
    wire signal_19402 ;
    wire signal_19403 ;
    wire signal_19404 ;
    wire signal_19405 ;
    wire signal_19406 ;
    wire signal_19407 ;
    wire signal_19408 ;
    wire signal_19409 ;
    wire signal_19410 ;
    wire signal_19411 ;
    wire signal_19412 ;
    wire signal_19413 ;
    wire signal_19414 ;
    wire signal_19415 ;
    wire signal_19416 ;
    wire signal_19417 ;
    wire signal_19418 ;
    wire signal_19419 ;
    wire signal_19420 ;
    wire signal_19421 ;
    wire signal_19422 ;
    wire signal_19423 ;
    wire signal_19424 ;
    wire signal_19425 ;
    wire signal_19426 ;
    wire signal_19427 ;
    wire signal_19428 ;
    wire signal_19429 ;
    wire signal_19430 ;
    wire signal_19431 ;
    wire signal_19432 ;
    wire signal_19433 ;
    wire signal_19434 ;
    wire signal_19435 ;
    wire signal_19436 ;
    wire signal_19437 ;
    wire signal_19438 ;
    wire signal_19439 ;
    wire signal_19440 ;
    wire signal_19441 ;
    wire signal_19442 ;
    wire signal_19443 ;
    wire signal_19444 ;
    wire signal_19445 ;
    wire signal_19446 ;
    wire signal_19447 ;
    wire signal_19448 ;
    wire signal_19449 ;
    wire signal_19450 ;
    wire signal_19451 ;
    wire signal_19452 ;
    wire signal_19453 ;
    wire signal_19454 ;
    wire signal_19455 ;
    wire signal_19456 ;
    wire signal_19457 ;
    wire signal_19458 ;
    wire signal_19459 ;
    wire signal_19460 ;
    wire signal_19461 ;
    wire signal_19462 ;
    wire signal_19463 ;
    wire signal_19464 ;
    wire signal_19465 ;
    wire signal_19466 ;
    wire signal_19467 ;
    wire signal_19468 ;
    wire signal_19469 ;
    wire signal_19470 ;
    wire signal_19471 ;
    wire signal_19472 ;
    wire signal_19473 ;
    wire signal_19474 ;
    wire signal_19475 ;
    wire signal_19476 ;
    wire signal_19477 ;
    wire signal_19478 ;
    wire signal_19479 ;
    wire signal_19480 ;
    wire signal_19481 ;
    wire signal_19482 ;
    wire signal_19483 ;
    wire signal_19484 ;
    wire signal_19485 ;
    wire signal_19486 ;
    wire signal_19487 ;
    wire signal_19488 ;
    wire signal_19489 ;
    wire signal_19490 ;
    wire signal_19491 ;
    wire signal_19492 ;
    wire signal_19493 ;
    wire signal_19494 ;
    wire signal_19495 ;
    wire signal_19496 ;
    wire signal_19497 ;
    wire signal_19498 ;
    wire signal_19499 ;
    wire signal_19500 ;
    wire signal_19501 ;
    wire signal_19502 ;
    wire signal_19503 ;
    wire signal_19504 ;
    wire signal_19505 ;
    wire signal_19506 ;
    wire signal_19507 ;
    wire signal_19508 ;
    wire signal_19509 ;
    wire signal_19510 ;
    wire signal_19511 ;
    wire signal_19512 ;
    wire signal_19513 ;
    wire signal_19514 ;
    wire signal_19515 ;
    wire signal_19516 ;
    wire signal_19517 ;
    wire signal_19518 ;
    wire signal_19519 ;
    wire signal_19520 ;
    wire signal_19521 ;
    wire signal_19522 ;
    wire signal_19523 ;
    wire signal_19524 ;
    wire signal_19525 ;
    wire signal_19526 ;
    wire signal_19527 ;
    wire signal_19528 ;
    wire signal_19529 ;
    wire signal_19530 ;
    wire signal_19531 ;
    wire signal_19532 ;
    wire signal_19533 ;
    wire signal_19534 ;
    wire signal_19535 ;
    wire signal_19536 ;
    wire signal_19537 ;
    wire signal_19538 ;
    wire signal_19539 ;
    wire signal_19540 ;
    wire signal_19541 ;
    wire signal_19542 ;
    wire signal_19543 ;
    wire signal_19544 ;
    wire signal_19545 ;
    wire signal_19546 ;
    wire signal_19547 ;
    wire signal_19548 ;
    wire signal_19549 ;
    wire signal_19550 ;
    wire signal_19551 ;
    wire signal_19552 ;
    wire signal_19553 ;
    wire signal_19554 ;
    wire signal_19555 ;
    wire signal_19556 ;
    wire signal_19557 ;
    wire signal_19558 ;
    wire signal_19559 ;
    wire signal_19560 ;
    wire signal_19561 ;
    wire signal_19562 ;
    wire signal_19563 ;
    wire signal_19564 ;
    wire signal_19565 ;
    wire signal_19566 ;
    wire signal_19567 ;
    wire signal_19568 ;
    wire signal_19569 ;
    wire signal_19570 ;
    wire signal_19571 ;
    wire signal_19572 ;
    wire signal_19573 ;
    wire signal_19574 ;
    wire signal_19575 ;
    wire signal_19576 ;
    wire signal_19577 ;
    wire signal_19578 ;
    wire signal_19579 ;
    wire signal_19580 ;
    wire signal_19581 ;
    wire signal_19582 ;
    wire signal_19583 ;
    wire signal_19584 ;
    wire signal_19585 ;
    wire signal_19586 ;
    wire signal_19587 ;
    wire signal_19588 ;
    wire signal_19589 ;
    wire signal_19590 ;
    wire signal_19591 ;
    wire signal_19592 ;
    wire signal_19593 ;
    wire signal_19594 ;
    wire signal_19595 ;
    wire signal_19596 ;
    wire signal_19597 ;
    wire signal_19598 ;
    wire signal_19599 ;
    wire signal_19600 ;
    wire signal_19601 ;
    wire signal_19602 ;
    wire signal_19603 ;
    wire signal_19604 ;
    wire signal_19605 ;
    wire signal_19606 ;
    wire signal_19607 ;
    wire signal_19608 ;
    wire signal_19609 ;
    wire signal_19610 ;
    wire signal_19611 ;
    wire signal_19612 ;
    wire signal_19613 ;
    wire signal_19614 ;
    wire signal_19615 ;
    wire signal_19616 ;
    wire signal_19617 ;
    wire signal_19618 ;
    wire signal_19619 ;
    wire signal_19620 ;
    wire signal_19621 ;
    wire signal_19622 ;
    wire signal_19623 ;
    wire signal_19624 ;
    wire signal_19625 ;
    wire signal_19626 ;
    wire signal_19627 ;
    wire signal_19628 ;
    wire signal_19629 ;
    wire signal_19630 ;
    wire signal_19631 ;
    wire signal_19632 ;
    wire signal_19633 ;
    wire signal_19634 ;
    wire signal_19635 ;
    wire signal_19636 ;
    wire signal_19637 ;
    wire signal_19638 ;
    wire signal_19639 ;
    wire signal_19640 ;
    wire signal_19641 ;
    wire signal_19642 ;
    wire signal_19643 ;
    wire signal_19644 ;
    wire signal_19645 ;
    wire signal_19646 ;
    wire signal_19647 ;
    wire signal_19648 ;
    wire signal_19649 ;
    wire signal_19650 ;
    wire signal_19651 ;
    wire signal_19652 ;
    wire signal_19653 ;
    wire signal_19654 ;
    wire signal_19655 ;
    wire signal_19656 ;
    wire signal_19657 ;
    wire signal_19658 ;
    wire signal_19659 ;
    wire signal_19660 ;
    wire signal_19661 ;
    wire signal_19662 ;
    wire signal_19663 ;
    wire signal_19664 ;
    wire signal_19665 ;
    wire signal_19666 ;
    wire signal_19667 ;
    wire signal_19668 ;
    wire signal_19669 ;
    wire signal_19670 ;
    wire signal_19671 ;
    wire signal_19672 ;
    wire signal_19673 ;
    wire signal_19674 ;
    wire signal_19675 ;
    wire signal_19676 ;
    wire signal_19677 ;
    wire signal_19678 ;
    wire signal_19679 ;
    wire signal_19680 ;
    wire signal_19681 ;
    wire signal_19682 ;
    wire signal_19683 ;
    wire signal_19684 ;
    wire signal_19685 ;
    wire signal_19686 ;
    wire signal_19687 ;
    wire signal_19688 ;
    wire signal_19689 ;
    wire signal_19690 ;
    wire signal_19691 ;
    wire signal_19692 ;
    wire signal_19693 ;
    wire signal_19694 ;
    wire signal_19695 ;
    wire signal_19696 ;
    wire signal_19697 ;
    wire signal_19698 ;
    wire signal_19699 ;
    wire signal_19700 ;
    wire signal_19701 ;
    wire signal_19702 ;
    wire signal_19703 ;
    wire signal_19704 ;
    wire signal_19705 ;
    wire signal_19706 ;
    wire signal_19707 ;
    wire signal_19708 ;
    wire signal_19709 ;
    wire signal_19710 ;
    wire signal_19711 ;
    wire signal_19712 ;
    wire signal_19713 ;
    wire signal_19714 ;
    wire signal_19715 ;
    wire signal_19716 ;
    wire signal_19717 ;
    wire signal_19718 ;
    wire signal_19719 ;
    wire signal_19720 ;
    wire signal_19721 ;
    wire signal_19722 ;
    wire signal_19723 ;
    wire signal_19724 ;
    wire signal_19725 ;
    wire signal_19726 ;
    wire signal_19727 ;
    wire signal_19728 ;
    wire signal_19729 ;
    wire signal_19730 ;
    wire signal_19731 ;
    wire signal_19732 ;
    wire signal_19733 ;
    wire signal_19734 ;
    wire signal_19735 ;
    wire signal_19736 ;
    wire signal_19737 ;
    wire signal_19738 ;
    wire signal_19739 ;
    wire signal_19740 ;
    wire signal_19741 ;
    wire signal_19742 ;
    wire signal_19743 ;
    wire signal_19744 ;
    wire signal_19745 ;
    wire signal_19746 ;
    wire signal_19747 ;
    wire signal_19748 ;
    wire signal_19749 ;
    wire signal_19750 ;
    wire signal_19751 ;
    wire signal_19752 ;
    wire signal_19753 ;
    wire signal_19754 ;
    wire signal_19755 ;
    wire signal_19756 ;
    wire signal_19757 ;
    wire signal_19758 ;
    wire signal_19759 ;
    wire signal_19760 ;
    wire signal_19761 ;
    wire signal_19762 ;
    wire signal_19763 ;
    wire signal_19764 ;
    wire signal_19765 ;
    wire signal_19766 ;
    wire signal_19767 ;
    wire signal_19768 ;
    wire signal_19769 ;
    wire signal_19770 ;
    wire signal_19771 ;
    wire signal_19772 ;
    wire signal_19773 ;
    wire signal_19774 ;
    wire signal_19775 ;
    wire signal_19776 ;
    wire signal_19777 ;
    wire signal_19778 ;
    wire signal_19779 ;
    wire signal_19780 ;
    wire signal_19781 ;
    wire signal_19782 ;
    wire signal_19783 ;
    wire signal_19784 ;
    wire signal_19785 ;
    wire signal_19786 ;
    wire signal_19787 ;
    wire signal_19788 ;
    wire signal_19789 ;
    wire signal_19790 ;
    wire signal_19791 ;
    wire signal_19792 ;
    wire signal_19793 ;
    wire signal_19794 ;
    wire signal_19795 ;
    wire signal_19796 ;
    wire signal_19797 ;
    wire signal_19798 ;
    wire signal_19799 ;
    wire signal_19800 ;
    wire signal_19801 ;
    wire signal_19802 ;
    wire signal_19803 ;
    wire signal_19804 ;
    wire signal_19805 ;
    wire signal_19806 ;
    wire signal_19807 ;
    wire signal_19808 ;
    wire signal_19809 ;
    wire signal_19810 ;
    wire signal_19811 ;
    wire signal_19812 ;
    wire signal_19813 ;
    wire signal_19814 ;
    wire signal_19815 ;
    wire signal_19816 ;
    wire signal_19817 ;
    wire signal_19818 ;
    wire signal_19819 ;
    wire signal_19820 ;
    wire signal_19821 ;
    wire signal_19822 ;
    wire signal_19823 ;
    wire signal_19824 ;
    wire signal_19825 ;
    wire signal_19826 ;
    wire signal_19827 ;
    wire signal_19828 ;
    wire signal_19829 ;
    wire signal_19830 ;
    wire signal_19831 ;
    wire signal_19832 ;
    wire signal_19833 ;
    wire signal_19834 ;
    wire signal_19835 ;
    wire signal_19836 ;
    wire signal_19837 ;
    wire signal_19838 ;
    wire signal_19839 ;
    wire signal_19840 ;
    wire signal_19841 ;
    wire signal_19842 ;
    wire signal_19843 ;
    wire signal_19844 ;
    wire signal_19845 ;
    wire signal_19846 ;
    wire signal_19847 ;
    wire signal_19848 ;
    wire signal_19849 ;
    wire signal_19850 ;
    wire signal_19851 ;
    wire signal_19852 ;
    wire signal_19853 ;
    wire signal_19854 ;
    wire signal_19855 ;
    wire signal_19856 ;
    wire signal_19857 ;
    wire signal_19858 ;
    wire signal_19859 ;
    wire signal_19860 ;
    wire signal_19861 ;
    wire signal_19862 ;
    wire signal_19863 ;
    wire signal_19864 ;
    wire signal_19865 ;
    wire signal_19866 ;
    wire signal_19867 ;
    wire signal_19868 ;
    wire signal_19869 ;
    wire signal_19870 ;
    wire signal_19871 ;
    wire signal_19872 ;
    wire signal_19873 ;
    wire signal_19874 ;
    wire signal_19875 ;
    wire signal_19876 ;
    wire signal_19877 ;
    wire signal_19878 ;
    wire signal_19879 ;
    wire signal_19880 ;
    wire signal_19881 ;
    wire signal_19882 ;
    wire signal_19883 ;
    wire signal_19884 ;
    wire signal_19885 ;
    wire signal_19886 ;
    wire signal_19887 ;
    wire signal_19888 ;
    wire signal_19889 ;
    wire signal_19890 ;
    wire signal_19891 ;
    wire signal_19892 ;
    wire signal_19893 ;
    wire signal_19894 ;
    wire signal_19895 ;
    wire signal_19896 ;
    wire signal_19897 ;
    wire signal_19898 ;
    wire signal_19899 ;
    wire signal_19900 ;
    wire signal_19901 ;
    wire signal_19902 ;
    wire signal_19903 ;
    wire signal_19904 ;
    wire signal_19905 ;
    wire signal_19906 ;
    wire signal_19907 ;
    wire signal_19908 ;
    wire signal_19909 ;
    wire signal_19910 ;
    wire signal_19911 ;
    wire signal_19912 ;
    wire signal_19913 ;
    wire signal_19914 ;
    wire signal_19915 ;
    wire signal_19916 ;
    wire signal_19917 ;
    wire signal_19918 ;
    wire signal_19919 ;
    wire signal_19920 ;
    wire signal_19921 ;
    wire signal_19922 ;
    wire signal_19923 ;
    wire signal_19924 ;
    wire signal_19925 ;
    wire signal_19926 ;
    wire signal_19927 ;
    wire signal_19928 ;
    wire signal_19929 ;
    wire signal_19930 ;
    wire signal_19931 ;
    wire signal_19932 ;
    wire signal_19933 ;
    wire signal_19934 ;
    wire signal_19935 ;
    wire signal_19936 ;
    wire signal_19937 ;
    wire signal_19938 ;
    wire signal_19939 ;
    wire signal_19940 ;
    wire signal_19941 ;
    wire signal_19942 ;
    wire signal_19943 ;
    wire signal_19944 ;
    wire signal_19945 ;
    wire signal_19946 ;
    wire signal_19947 ;
    wire signal_19948 ;
    wire signal_19949 ;
    wire signal_19950 ;
    wire signal_19951 ;
    wire signal_19952 ;
    wire signal_19953 ;
    wire signal_19954 ;
    wire signal_19955 ;
    wire signal_19956 ;
    wire signal_19957 ;
    wire signal_19958 ;
    wire signal_19959 ;
    wire signal_19960 ;
    wire signal_19961 ;
    wire signal_19962 ;
    wire signal_19963 ;
    wire signal_19964 ;
    wire signal_19965 ;
    wire signal_19966 ;
    wire signal_19967 ;
    wire signal_19968 ;
    wire signal_19969 ;
    wire signal_19970 ;
    wire signal_19971 ;
    wire signal_19972 ;
    wire signal_19973 ;
    wire signal_19974 ;
    wire signal_19975 ;
    wire signal_19976 ;
    wire signal_19977 ;
    wire signal_19978 ;
    wire signal_19979 ;
    wire signal_19980 ;
    wire signal_19981 ;
    wire signal_19982 ;
    wire signal_19983 ;
    wire signal_19984 ;
    wire signal_19985 ;
    wire signal_19986 ;
    wire signal_19987 ;
    wire signal_19988 ;
    wire signal_19989 ;
    wire signal_19990 ;
    wire signal_19991 ;
    wire signal_19992 ;
    wire signal_19993 ;
    wire signal_19994 ;
    wire signal_19995 ;
    wire signal_19996 ;
    wire signal_19997 ;
    wire signal_19998 ;
    wire signal_19999 ;
    wire signal_20000 ;
    wire signal_20001 ;
    wire signal_20002 ;
    wire signal_20003 ;
    wire signal_20004 ;
    wire signal_20005 ;
    wire signal_20006 ;
    wire signal_20007 ;
    wire signal_20008 ;
    wire signal_20009 ;
    wire signal_20010 ;
    wire signal_20011 ;
    wire signal_20012 ;
    wire signal_20013 ;
    wire signal_20014 ;
    wire signal_20015 ;
    wire signal_20016 ;
    wire signal_20017 ;
    wire signal_20018 ;
    wire signal_20019 ;
    wire signal_20020 ;
    wire signal_20021 ;
    wire signal_20022 ;
    wire signal_20023 ;
    wire signal_20024 ;
    wire signal_20025 ;
    wire signal_20026 ;
    wire signal_20027 ;
    wire signal_20028 ;
    wire signal_20029 ;
    wire signal_20030 ;
    wire signal_20031 ;
    wire signal_20032 ;
    wire signal_20033 ;
    wire signal_20034 ;
    wire signal_20035 ;
    wire signal_20036 ;
    wire signal_20037 ;
    wire signal_20038 ;
    wire signal_20039 ;
    wire signal_20040 ;
    wire signal_20041 ;
    wire signal_20042 ;
    wire signal_20043 ;
    wire signal_20044 ;
    wire signal_20045 ;
    wire signal_20046 ;
    wire signal_20047 ;
    wire signal_20048 ;
    wire signal_20049 ;
    wire signal_20050 ;
    wire signal_20051 ;
    wire signal_20052 ;
    wire signal_20053 ;
    wire signal_20054 ;
    wire signal_20055 ;
    wire signal_20056 ;
    wire signal_20057 ;
    wire signal_20058 ;
    wire signal_20059 ;
    wire signal_20060 ;
    wire signal_20061 ;
    wire signal_20062 ;
    wire signal_20063 ;
    wire signal_20064 ;
    wire signal_20065 ;
    wire signal_20066 ;
    wire signal_20067 ;
    wire signal_20068 ;
    wire signal_20069 ;
    wire signal_20070 ;
    wire signal_20071 ;
    wire signal_20072 ;
    wire signal_20073 ;
    wire signal_20074 ;
    wire signal_20075 ;
    wire signal_20076 ;
    wire signal_20077 ;
    wire signal_20078 ;
    wire signal_20079 ;
    wire signal_20080 ;
    wire signal_20081 ;
    wire signal_20082 ;
    wire signal_20083 ;
    wire signal_20084 ;
    wire signal_20085 ;
    wire signal_20086 ;
    wire signal_20087 ;
    wire signal_20088 ;
    wire signal_20089 ;
    wire signal_20090 ;
    wire signal_20091 ;
    wire signal_20092 ;
    wire signal_20093 ;
    wire signal_20094 ;
    wire signal_20095 ;
    wire signal_20096 ;
    wire signal_20097 ;
    wire signal_20098 ;
    wire signal_20099 ;
    wire signal_20100 ;
    wire signal_20101 ;
    wire signal_20102 ;
    wire signal_20103 ;
    wire signal_20104 ;
    wire signal_20105 ;
    wire signal_20106 ;
    wire signal_20107 ;
    wire signal_20108 ;
    wire signal_20109 ;
    wire signal_20110 ;
    wire signal_20111 ;
    wire signal_20112 ;
    wire signal_20113 ;
    wire signal_20114 ;
    wire signal_20115 ;
    wire signal_20116 ;
    wire signal_20117 ;
    wire signal_20118 ;
    wire signal_20119 ;
    wire signal_20120 ;
    wire signal_20121 ;
    wire signal_20122 ;
    wire signal_20123 ;
    wire signal_20124 ;
    wire signal_20125 ;
    wire signal_20126 ;
    wire signal_20127 ;
    wire signal_20128 ;
    wire signal_20129 ;
    wire signal_20130 ;
    wire signal_20131 ;
    wire signal_20132 ;
    wire signal_20133 ;
    wire signal_20134 ;
    wire signal_20135 ;
    wire signal_20136 ;
    wire signal_20137 ;
    wire signal_20138 ;
    wire signal_20139 ;
    wire signal_20140 ;
    wire signal_20141 ;
    wire signal_20142 ;
    wire signal_20143 ;
    wire signal_20144 ;
    wire signal_20145 ;
    wire signal_20146 ;
    wire signal_20147 ;
    wire signal_20148 ;
    wire signal_20149 ;
    wire signal_20150 ;
    wire signal_20151 ;
    wire signal_20152 ;
    wire signal_20153 ;
    wire signal_20154 ;
    wire signal_20155 ;
    wire signal_20156 ;
    wire signal_20157 ;
    wire signal_20158 ;
    wire signal_20159 ;
    wire signal_20160 ;
    wire signal_20161 ;
    wire signal_20162 ;
    wire signal_20163 ;
    wire signal_20164 ;
    wire signal_20165 ;
    wire signal_20166 ;
    wire signal_20167 ;
    wire signal_20168 ;
    wire signal_20169 ;
    wire signal_20170 ;
    wire signal_20171 ;
    wire signal_20172 ;
    wire signal_20173 ;
    wire signal_20174 ;
    wire signal_20175 ;
    wire signal_20176 ;
    wire signal_20177 ;
    wire signal_20178 ;
    wire signal_20179 ;
    wire signal_20180 ;
    wire signal_20181 ;
    wire signal_20182 ;
    wire signal_20183 ;
    wire signal_20184 ;
    wire signal_20185 ;
    wire signal_20186 ;
    wire signal_20187 ;
    wire signal_20188 ;
    wire signal_20189 ;
    wire signal_20190 ;
    wire signal_20191 ;
    wire signal_20192 ;
    wire signal_20193 ;
    wire signal_20194 ;
    wire signal_20195 ;
    wire signal_20196 ;
    wire signal_20197 ;
    wire signal_20198 ;
    wire signal_20199 ;
    wire signal_20200 ;
    wire signal_20201 ;
    wire signal_20202 ;
    wire signal_20203 ;
    wire signal_20204 ;
    wire signal_20205 ;
    wire signal_20206 ;
    wire signal_20207 ;
    wire signal_20208 ;
    wire signal_20209 ;
    wire signal_20210 ;
    wire signal_20211 ;
    wire signal_20212 ;
    wire signal_20213 ;
    wire signal_20214 ;
    wire signal_20215 ;
    wire signal_20216 ;
    wire signal_20217 ;
    wire signal_20218 ;
    wire signal_20219 ;
    wire signal_20220 ;
    wire signal_20221 ;
    wire signal_20222 ;
    wire signal_20223 ;
    wire signal_20224 ;
    wire signal_20225 ;
    wire signal_20226 ;
    wire signal_20227 ;
    wire signal_20228 ;
    wire signal_20229 ;
    wire signal_20230 ;
    wire signal_20231 ;
    wire signal_20232 ;
    wire signal_20233 ;
    wire signal_20234 ;
    wire signal_20235 ;
    wire signal_20236 ;
    wire signal_20237 ;
    wire signal_20238 ;
    wire signal_20239 ;
    wire signal_20240 ;
    wire signal_20241 ;
    wire signal_20242 ;
    wire signal_20243 ;
    wire signal_20244 ;
    wire signal_20245 ;
    wire signal_20246 ;
    wire signal_20247 ;
    wire signal_20248 ;
    wire signal_20249 ;
    wire signal_20250 ;
    wire signal_20251 ;
    wire signal_20252 ;
    wire signal_20253 ;
    wire signal_20254 ;
    wire signal_20255 ;
    wire signal_20256 ;
    wire signal_20257 ;
    wire signal_20258 ;
    wire signal_20259 ;
    wire signal_20260 ;
    wire signal_20261 ;
    wire signal_20262 ;
    wire signal_20263 ;
    wire signal_20264 ;
    wire signal_20265 ;
    wire signal_20266 ;
    wire signal_20267 ;
    wire signal_20268 ;
    wire signal_20269 ;
    wire signal_20270 ;
    wire signal_20271 ;
    wire signal_20272 ;
    wire signal_20273 ;
    wire signal_20274 ;
    wire signal_20275 ;
    wire signal_20276 ;
    wire signal_20277 ;
    wire signal_20278 ;
    wire signal_20279 ;
    wire signal_20280 ;
    wire signal_20281 ;
    wire signal_20282 ;
    wire signal_20283 ;
    wire signal_20284 ;
    wire signal_20285 ;
    wire signal_20286 ;
    wire signal_20287 ;
    wire signal_20288 ;
    wire signal_20289 ;
    wire signal_20290 ;
    wire signal_20291 ;
    wire signal_20292 ;
    wire signal_20293 ;
    wire signal_20294 ;
    wire signal_20295 ;
    wire signal_20296 ;
    wire signal_20297 ;
    wire signal_20298 ;
    wire signal_20299 ;
    wire signal_20300 ;
    wire signal_20301 ;
    wire signal_20302 ;
    wire signal_20303 ;
    wire signal_20304 ;
    wire signal_20305 ;
    wire signal_20306 ;
    wire signal_20307 ;
    wire signal_20308 ;
    wire signal_20309 ;
    wire signal_20310 ;
    wire signal_20311 ;
    wire signal_20312 ;
    wire signal_20313 ;
    wire signal_20314 ;
    wire signal_20315 ;
    wire signal_20316 ;
    wire signal_20317 ;
    wire signal_20318 ;
    wire signal_20319 ;
    wire signal_20320 ;
    wire signal_20321 ;
    wire signal_20322 ;
    wire signal_20323 ;
    wire signal_20324 ;
    wire signal_20325 ;
    wire signal_20326 ;
    wire signal_20327 ;
    wire signal_20328 ;
    wire signal_20329 ;
    wire signal_20330 ;
    wire signal_20331 ;
    wire signal_20332 ;
    wire signal_20333 ;
    wire signal_20334 ;
    wire signal_20335 ;
    wire signal_20336 ;
    wire signal_20337 ;
    wire signal_20338 ;
    wire signal_20339 ;
    wire signal_20340 ;
    wire signal_20341 ;
    wire signal_20342 ;
    wire signal_20343 ;
    wire signal_20344 ;
    wire signal_20345 ;
    wire signal_20346 ;
    wire signal_20347 ;
    wire signal_20348 ;
    wire signal_20349 ;
    wire signal_20350 ;
    wire signal_20351 ;
    wire signal_20352 ;
    wire signal_20353 ;
    wire signal_20354 ;
    wire signal_20355 ;
    wire signal_20356 ;
    wire signal_20357 ;
    wire signal_20358 ;
    wire signal_20359 ;
    wire signal_20360 ;
    wire signal_20361 ;
    wire signal_20362 ;
    wire signal_20363 ;
    wire signal_20364 ;
    wire signal_20365 ;
    wire signal_20366 ;
    wire signal_20367 ;
    wire signal_20368 ;
    wire signal_20369 ;
    wire signal_20370 ;
    wire signal_20371 ;
    wire signal_20372 ;
    wire signal_20373 ;
    wire signal_20374 ;
    wire signal_20375 ;
    wire signal_20376 ;
    wire signal_20377 ;
    wire signal_20378 ;
    wire signal_20379 ;
    wire signal_20380 ;
    wire signal_20381 ;
    wire signal_20382 ;
    wire signal_20383 ;
    wire signal_20384 ;
    wire signal_20385 ;
    wire signal_20386 ;
    wire signal_20387 ;
    wire signal_20388 ;
    wire signal_20389 ;
    wire signal_20390 ;
    wire signal_20391 ;
    wire signal_20392 ;
    wire signal_20393 ;
    wire signal_20394 ;
    wire signal_20395 ;
    wire signal_20396 ;
    wire signal_20397 ;
    wire signal_20398 ;
    wire signal_20399 ;
    wire signal_20400 ;
    wire signal_20401 ;
    wire signal_20402 ;
    wire signal_20403 ;
    wire signal_20404 ;
    wire signal_20405 ;
    wire signal_20406 ;
    wire signal_20407 ;
    wire signal_20408 ;
    wire signal_20409 ;
    wire signal_20410 ;
    wire signal_20411 ;
    wire signal_20412 ;
    wire signal_20413 ;
    wire signal_20414 ;
    wire signal_20415 ;
    wire signal_20416 ;
    wire signal_20417 ;
    wire signal_20418 ;
    wire signal_20419 ;
    wire signal_20420 ;
    wire signal_20421 ;
    wire signal_20422 ;
    wire signal_20423 ;
    wire signal_20424 ;
    wire signal_20425 ;
    wire signal_20426 ;
    wire signal_20427 ;
    wire signal_20428 ;
    wire signal_20429 ;
    wire signal_20430 ;
    wire signal_20431 ;
    wire signal_20432 ;
    wire signal_20433 ;
    wire signal_20434 ;
    wire signal_20435 ;
    wire signal_20436 ;
    wire signal_20437 ;
    wire signal_20438 ;
    wire signal_20439 ;
    wire signal_20440 ;
    wire signal_20441 ;
    wire signal_20442 ;
    wire signal_20443 ;
    wire signal_20444 ;
    wire signal_20445 ;
    wire signal_20446 ;
    wire signal_20447 ;
    wire signal_20448 ;
    wire signal_20449 ;
    wire signal_20450 ;
    wire signal_20451 ;
    wire signal_20452 ;
    wire signal_20453 ;
    wire signal_20454 ;
    wire signal_20455 ;
    wire signal_20456 ;
    wire signal_20457 ;
    wire signal_20458 ;
    wire signal_20459 ;
    wire signal_20460 ;
    wire signal_20461 ;
    wire signal_20462 ;
    wire signal_20463 ;
    wire signal_20464 ;
    wire signal_20465 ;
    wire signal_20466 ;
    wire signal_20467 ;
    wire signal_20468 ;
    wire signal_20469 ;
    wire signal_20470 ;
    wire signal_20471 ;
    wire signal_20472 ;
    wire signal_20473 ;
    wire signal_20474 ;
    wire signal_20475 ;
    wire signal_20476 ;
    wire signal_20477 ;
    wire signal_20478 ;
    wire signal_20479 ;
    wire signal_20480 ;
    wire signal_20481 ;
    wire signal_20482 ;
    wire signal_20483 ;
    wire signal_20484 ;
    wire signal_20485 ;
    wire signal_20486 ;
    wire signal_20487 ;
    wire signal_20488 ;
    wire signal_20489 ;
    wire signal_20490 ;
    wire signal_20491 ;
    wire signal_20492 ;
    wire signal_20493 ;
    wire signal_20494 ;
    wire signal_20495 ;
    wire signal_20496 ;
    wire signal_20497 ;
    wire signal_20498 ;
    wire signal_20499 ;
    wire signal_20500 ;
    wire signal_20501 ;
    wire signal_20502 ;
    wire signal_20503 ;
    wire signal_20504 ;
    wire signal_20505 ;
    wire signal_20506 ;
    wire signal_20507 ;
    wire signal_20508 ;
    wire signal_20509 ;
    wire signal_20510 ;
    wire signal_20511 ;
    wire signal_20512 ;
    wire signal_20513 ;
    wire signal_20514 ;
    wire signal_20515 ;
    wire signal_20516 ;
    wire signal_20517 ;
    wire signal_20518 ;
    wire signal_20519 ;
    wire signal_20520 ;
    wire signal_20521 ;
    wire signal_20522 ;
    wire signal_20523 ;
    wire signal_20524 ;
    wire signal_20525 ;
    wire signal_20526 ;
    wire signal_20527 ;
    wire signal_20528 ;
    wire signal_20529 ;
    wire signal_20530 ;
    wire signal_20531 ;
    wire signal_20532 ;
    wire signal_20533 ;
    wire signal_20534 ;
    wire signal_20535 ;
    wire signal_20536 ;
    wire signal_20537 ;
    wire signal_20538 ;
    wire signal_20539 ;
    wire signal_20540 ;
    wire signal_20541 ;
    wire signal_20542 ;
    wire signal_20543 ;
    wire signal_20544 ;
    wire signal_20545 ;
    wire signal_20546 ;
    wire signal_20547 ;
    wire signal_20548 ;
    wire signal_20549 ;
    wire signal_20550 ;
    wire signal_20551 ;
    wire signal_20552 ;
    wire signal_20553 ;
    wire signal_20554 ;
    wire signal_20555 ;
    wire signal_20556 ;
    wire signal_20557 ;
    wire signal_20558 ;
    wire signal_20559 ;
    wire signal_20560 ;
    wire signal_20561 ;
    wire signal_20562 ;
    wire signal_20563 ;
    wire signal_20564 ;
    wire signal_20565 ;
    wire signal_20566 ;
    wire signal_20567 ;
    wire signal_20568 ;
    wire signal_20569 ;
    wire signal_20570 ;
    wire signal_20571 ;
    wire signal_20572 ;
    wire signal_20573 ;
    wire signal_20574 ;
    wire signal_20575 ;
    wire signal_20576 ;
    wire signal_20577 ;
    wire signal_20578 ;
    wire signal_20579 ;
    wire signal_20580 ;
    wire signal_20581 ;
    wire signal_20582 ;
    wire signal_20583 ;
    wire signal_20584 ;
    wire signal_20585 ;
    wire signal_20586 ;
    wire signal_20587 ;
    wire signal_20588 ;
    wire signal_20589 ;
    wire signal_20590 ;
    wire signal_20591 ;
    wire signal_20592 ;
    wire signal_20593 ;
    wire signal_20594 ;
    wire signal_20595 ;
    wire signal_20596 ;
    wire signal_20597 ;
    wire signal_20598 ;
    wire signal_20599 ;
    wire signal_20600 ;
    wire signal_20601 ;
    wire signal_20602 ;
    wire signal_20603 ;
    wire signal_20604 ;
    wire signal_20605 ;
    wire signal_20606 ;
    wire signal_20607 ;
    wire signal_20608 ;
    wire signal_20609 ;
    wire signal_20610 ;
    wire signal_20611 ;
    wire signal_20612 ;
    wire signal_20613 ;
    wire signal_20614 ;
    wire signal_20615 ;
    wire signal_20616 ;
    wire signal_20617 ;
    wire signal_20618 ;
    wire signal_20619 ;
    wire signal_20620 ;
    wire signal_20621 ;
    wire signal_20622 ;
    wire signal_20623 ;
    wire signal_20624 ;
    wire signal_20625 ;
    wire signal_20626 ;
    wire signal_20627 ;
    wire signal_20628 ;
    wire signal_20629 ;
    wire signal_20630 ;
    wire signal_20631 ;
    wire signal_20632 ;
    wire signal_20633 ;
    wire signal_20634 ;
    wire signal_20635 ;
    wire signal_20636 ;
    wire signal_20637 ;
    wire signal_20638 ;
    wire signal_20639 ;
    wire signal_20640 ;
    wire signal_20641 ;
    wire signal_20642 ;
    wire signal_20643 ;
    wire signal_20644 ;
    wire signal_20645 ;
    wire signal_20646 ;
    wire signal_20647 ;
    wire signal_20648 ;
    wire signal_20649 ;
    wire signal_20650 ;
    wire signal_20651 ;
    wire signal_20652 ;
    wire signal_20653 ;
    wire signal_20654 ;
    wire signal_20655 ;
    wire signal_20656 ;
    wire signal_20657 ;
    wire signal_20658 ;
    wire signal_20659 ;
    wire signal_20660 ;
    wire signal_20661 ;
    wire signal_20662 ;
    wire signal_20663 ;
    wire signal_20664 ;
    wire signal_20665 ;
    wire signal_20666 ;
    wire signal_20667 ;
    wire signal_20668 ;
    wire signal_20669 ;
    wire signal_20670 ;
    wire signal_20671 ;
    wire signal_20672 ;
    wire signal_20673 ;
    wire signal_20674 ;
    wire signal_20675 ;
    wire signal_20676 ;
    wire signal_20677 ;
    wire signal_20678 ;
    wire signal_20679 ;
    wire signal_20680 ;
    wire signal_20681 ;
    wire signal_20682 ;
    wire signal_20683 ;
    wire signal_20684 ;
    wire signal_20685 ;
    wire signal_20686 ;
    wire signal_20687 ;
    wire signal_20688 ;
    wire signal_20689 ;
    wire signal_20690 ;
    wire signal_20691 ;
    wire signal_20692 ;
    wire signal_20693 ;
    wire signal_20694 ;
    wire signal_20695 ;
    wire signal_20696 ;
    wire signal_20697 ;
    wire signal_20698 ;
    wire signal_20699 ;
    wire signal_20700 ;
    wire signal_20701 ;
    wire signal_20702 ;
    wire signal_20703 ;
    wire signal_20704 ;
    wire signal_20705 ;
    wire signal_20706 ;
    wire signal_20707 ;
    wire signal_20708 ;
    wire signal_20709 ;
    wire signal_20710 ;
    wire signal_20711 ;
    wire signal_20712 ;
    wire signal_20713 ;
    wire signal_20714 ;
    wire signal_20715 ;
    wire signal_20716 ;
    wire signal_20717 ;
    wire signal_20718 ;
    wire signal_20719 ;
    wire signal_20720 ;
    wire signal_20721 ;
    wire signal_20722 ;
    wire signal_20723 ;
    wire signal_20724 ;
    wire signal_20725 ;
    wire signal_20726 ;
    wire signal_20727 ;
    wire signal_20728 ;
    wire signal_20729 ;
    wire signal_20730 ;
    wire signal_20731 ;
    wire signal_20732 ;
    wire signal_20733 ;
    wire signal_20734 ;
    wire signal_20735 ;
    wire signal_20736 ;
    wire signal_20737 ;
    wire signal_20738 ;
    wire signal_20739 ;
    wire signal_20740 ;
    wire signal_20741 ;
    wire signal_20742 ;
    wire signal_20743 ;
    wire signal_20744 ;
    wire signal_20745 ;
    wire signal_20746 ;
    wire signal_20747 ;
    wire signal_20748 ;
    wire signal_20749 ;
    wire signal_20750 ;
    wire signal_20751 ;
    wire signal_20752 ;
    wire signal_20753 ;
    wire signal_20754 ;
    wire signal_20755 ;
    wire signal_20756 ;
    wire signal_20757 ;
    wire signal_20758 ;
    wire signal_20759 ;
    wire signal_20760 ;
    wire signal_20761 ;
    wire signal_20762 ;
    wire signal_20763 ;
    wire signal_20764 ;
    wire signal_20765 ;
    wire signal_20766 ;
    wire signal_20767 ;
    wire signal_20768 ;
    wire signal_20769 ;
    wire signal_20770 ;
    wire signal_20771 ;
    wire signal_20772 ;
    wire signal_20773 ;
    wire signal_20774 ;
    wire signal_20775 ;
    wire signal_20776 ;
    wire signal_20777 ;
    wire signal_20778 ;
    wire signal_20779 ;
    wire signal_20780 ;
    wire signal_20781 ;
    wire signal_20782 ;
    wire signal_20783 ;
    wire signal_20784 ;
    wire signal_20785 ;
    wire signal_20786 ;
    wire signal_20787 ;
    wire signal_20788 ;
    wire signal_20789 ;
    wire signal_20790 ;
    wire signal_20791 ;
    wire signal_20792 ;
    wire signal_20793 ;
    wire signal_20794 ;
    wire signal_20795 ;
    wire signal_20796 ;
    wire signal_20797 ;
    wire signal_20798 ;
    wire signal_20799 ;
    wire signal_20800 ;
    wire signal_20801 ;
    wire signal_20802 ;
    wire signal_20803 ;
    wire signal_20804 ;
    wire signal_20805 ;
    wire signal_20806 ;
    wire signal_20807 ;
    wire signal_20808 ;
    wire signal_20809 ;
    wire signal_20810 ;
    wire signal_20811 ;
    wire signal_20812 ;
    wire signal_20813 ;
    wire signal_20814 ;
    wire signal_20815 ;
    wire signal_20816 ;
    wire signal_20817 ;
    wire signal_20818 ;
    wire signal_20819 ;
    wire signal_20820 ;
    wire signal_20821 ;
    wire signal_20822 ;
    wire signal_20823 ;
    wire signal_20824 ;
    wire signal_20825 ;
    wire signal_20826 ;
    wire signal_20827 ;
    wire signal_20828 ;
    wire signal_20829 ;
    wire signal_20830 ;
    wire signal_20831 ;
    wire signal_20832 ;
    wire signal_20833 ;
    wire signal_20834 ;
    wire signal_20835 ;
    wire signal_20836 ;
    wire signal_20837 ;
    wire signal_20838 ;
    wire signal_20839 ;
    wire signal_20840 ;
    wire signal_20841 ;
    wire signal_20842 ;
    wire signal_20843 ;
    wire signal_20844 ;
    wire signal_20845 ;
    wire signal_20846 ;
    wire signal_20847 ;
    wire signal_20848 ;
    wire signal_20849 ;
    wire signal_20850 ;
    wire signal_20851 ;
    wire signal_20852 ;
    wire signal_20853 ;
    wire signal_20854 ;
    wire signal_20855 ;
    wire signal_20856 ;
    wire signal_20857 ;
    wire signal_20858 ;
    wire signal_20859 ;
    wire signal_20860 ;
    wire signal_20861 ;
    wire signal_20862 ;
    wire signal_20863 ;
    wire signal_20864 ;
    wire signal_20865 ;
    wire signal_20866 ;
    wire signal_20867 ;
    wire signal_20868 ;
    wire signal_20869 ;
    wire signal_20870 ;
    wire signal_20871 ;
    wire signal_20872 ;
    wire signal_20873 ;
    wire signal_20874 ;
    wire signal_20875 ;
    wire signal_20876 ;
    wire signal_20877 ;
    wire signal_20878 ;
    wire signal_20879 ;
    wire signal_20880 ;
    wire signal_20881 ;
    wire signal_20882 ;
    wire signal_20883 ;
    wire signal_20884 ;
    wire signal_20885 ;
    wire signal_20886 ;
    wire signal_20887 ;
    wire signal_20888 ;
    wire signal_20889 ;
    wire signal_20890 ;
    wire signal_20891 ;
    wire signal_20892 ;
    wire signal_20893 ;
    wire signal_20894 ;
    wire signal_20895 ;
    wire signal_20896 ;
    wire signal_20897 ;
    wire signal_20898 ;
    wire signal_20899 ;
    wire signal_20900 ;
    wire signal_20901 ;
    wire signal_20902 ;
    wire signal_20903 ;
    wire signal_20904 ;
    wire signal_20905 ;
    wire signal_20906 ;
    wire signal_20907 ;
    wire signal_20908 ;
    wire signal_20909 ;
    wire signal_20910 ;
    wire signal_20911 ;
    wire signal_20912 ;
    wire signal_20913 ;
    wire signal_20914 ;
    wire signal_20915 ;
    wire signal_20916 ;
    wire signal_20917 ;
    wire signal_20918 ;
    wire signal_20919 ;
    wire signal_20920 ;
    wire signal_20921 ;
    wire signal_20922 ;
    wire signal_20923 ;
    wire signal_20924 ;
    wire signal_20925 ;
    wire signal_20926 ;
    wire signal_20927 ;
    wire signal_20928 ;
    wire signal_20929 ;
    wire signal_20930 ;
    wire signal_20931 ;
    wire signal_20932 ;
    wire signal_20933 ;
    wire signal_20934 ;
    wire signal_20935 ;
    wire signal_20936 ;
    wire signal_20937 ;
    wire signal_20938 ;
    wire signal_20939 ;
    wire signal_20940 ;
    wire signal_20941 ;
    wire signal_20942 ;
    wire signal_20943 ;
    wire signal_20944 ;
    wire signal_20945 ;
    wire signal_20946 ;
    wire signal_20947 ;
    wire signal_20948 ;
    wire signal_20949 ;
    wire signal_20950 ;
    wire signal_20951 ;
    wire signal_20952 ;
    wire signal_20953 ;
    wire signal_20954 ;
    wire signal_20955 ;
    wire signal_20956 ;
    wire signal_20957 ;
    wire signal_20958 ;
    wire signal_20959 ;
    wire signal_20960 ;
    wire signal_20961 ;
    wire signal_20962 ;
    wire signal_20963 ;
    wire signal_20964 ;
    wire signal_20965 ;
    wire signal_20966 ;
    wire signal_20967 ;
    wire signal_20968 ;
    wire signal_20969 ;
    wire signal_20970 ;
    wire signal_20971 ;
    wire signal_20972 ;
    wire signal_20973 ;
    wire signal_20974 ;
    wire signal_20975 ;
    wire signal_20976 ;
    wire signal_20977 ;
    wire signal_20978 ;
    wire signal_20979 ;
    wire signal_20980 ;
    wire signal_20981 ;
    wire signal_20982 ;
    wire signal_20983 ;
    wire signal_20984 ;
    wire signal_20985 ;
    wire signal_20986 ;
    wire signal_20987 ;
    wire signal_20988 ;
    wire signal_20989 ;
    wire signal_20990 ;
    wire signal_20991 ;
    wire signal_20992 ;
    wire signal_20993 ;
    wire signal_20994 ;
    wire signal_20995 ;
    wire signal_20996 ;
    wire signal_20997 ;
    wire signal_20998 ;
    wire signal_20999 ;
    wire signal_21000 ;
    wire signal_21001 ;
    wire signal_21002 ;
    wire signal_21003 ;
    wire signal_21004 ;
    wire signal_21005 ;
    wire signal_21006 ;
    wire signal_21007 ;
    wire signal_21008 ;
    wire signal_21009 ;
    wire signal_21010 ;
    wire signal_21011 ;
    wire signal_21012 ;
    wire signal_21013 ;
    wire signal_21014 ;
    wire signal_21015 ;
    wire signal_21016 ;
    wire signal_21017 ;
    wire signal_21018 ;
    wire signal_21019 ;
    wire signal_21020 ;
    wire signal_21021 ;
    wire signal_21022 ;
    wire signal_21023 ;
    wire signal_21024 ;
    wire signal_21025 ;
    wire signal_21026 ;
    wire signal_21027 ;
    wire signal_21028 ;
    wire signal_21029 ;
    wire signal_21030 ;
    wire signal_21031 ;
    wire signal_21032 ;
    wire signal_21033 ;
    wire signal_21034 ;
    wire signal_21035 ;
    wire signal_21036 ;
    wire signal_21037 ;
    wire signal_21038 ;
    wire signal_21039 ;
    wire signal_21040 ;
    wire signal_21041 ;
    wire signal_21042 ;
    wire signal_21043 ;
    wire signal_21044 ;
    wire signal_21045 ;
    wire signal_21046 ;
    wire signal_21047 ;
    wire signal_21048 ;
    wire signal_21049 ;
    wire signal_21050 ;
    wire signal_21051 ;
    wire signal_21052 ;
    wire signal_21053 ;
    wire signal_21054 ;
    wire signal_21055 ;
    wire signal_21056 ;
    wire signal_21057 ;
    wire signal_21058 ;
    wire signal_21059 ;
    wire signal_21060 ;
    wire signal_21061 ;
    wire signal_21062 ;
    wire signal_21063 ;
    wire signal_21064 ;
    wire signal_21065 ;
    wire signal_21066 ;
    wire signal_21067 ;
    wire signal_21068 ;
    wire signal_21069 ;
    wire signal_21070 ;
    wire signal_21071 ;
    wire signal_21072 ;
    wire signal_21073 ;
    wire signal_21074 ;
    wire signal_21075 ;
    wire signal_21076 ;
    wire signal_21077 ;
    wire signal_21078 ;
    wire signal_21079 ;
    wire signal_21080 ;
    wire signal_21081 ;
    wire signal_21082 ;
    wire signal_21083 ;
    wire signal_21084 ;
    wire signal_21085 ;
    wire signal_21086 ;
    wire signal_21087 ;
    wire signal_21088 ;
    wire signal_21089 ;
    wire signal_21090 ;
    wire signal_21091 ;
    wire signal_21092 ;
    wire signal_21093 ;
    wire signal_21094 ;
    wire signal_21095 ;
    wire signal_21096 ;
    wire signal_21097 ;
    wire signal_21098 ;
    wire signal_21099 ;
    wire signal_21100 ;
    wire signal_21101 ;
    wire signal_21102 ;
    wire signal_21103 ;
    wire signal_21104 ;
    wire signal_21105 ;
    wire signal_21106 ;
    wire signal_21107 ;
    wire signal_21108 ;
    wire signal_21109 ;
    wire signal_21110 ;
    wire signal_21111 ;
    wire signal_21112 ;
    wire signal_21113 ;
    wire signal_21114 ;
    wire signal_21115 ;
    wire signal_21116 ;
    wire signal_21117 ;
    wire signal_21118 ;
    wire signal_21119 ;
    wire signal_21120 ;
    wire signal_21121 ;
    wire signal_21122 ;
    wire signal_21123 ;
    wire signal_21124 ;
    wire signal_21125 ;
    wire signal_21126 ;
    wire signal_21127 ;
    wire signal_21128 ;
    wire signal_21129 ;
    wire signal_21130 ;
    wire signal_21131 ;
    wire signal_21132 ;
    wire signal_21133 ;
    wire signal_21134 ;
    wire signal_21135 ;
    wire signal_21136 ;
    wire signal_21137 ;
    wire signal_21138 ;
    wire signal_21139 ;
    wire signal_21140 ;
    wire signal_21141 ;
    wire signal_21142 ;
    wire signal_21143 ;
    wire signal_21144 ;
    wire signal_21145 ;
    wire signal_21146 ;
    wire signal_21147 ;
    wire signal_21148 ;
    wire signal_21149 ;
    wire signal_21150 ;
    wire signal_21151 ;
    wire signal_21152 ;
    wire signal_21153 ;
    wire signal_21154 ;
    wire signal_21155 ;
    wire signal_21156 ;
    wire signal_21157 ;
    wire signal_21158 ;
    wire signal_21159 ;
    wire signal_21160 ;
    wire signal_21161 ;
    wire signal_21162 ;
    wire signal_21163 ;
    wire signal_21164 ;
    wire signal_21165 ;
    wire signal_21166 ;
    wire signal_21167 ;
    wire signal_21168 ;
    wire signal_21169 ;
    wire signal_21170 ;
    wire signal_21171 ;
    wire signal_21172 ;
    wire signal_21173 ;
    wire signal_21174 ;
    wire signal_21175 ;
    wire signal_21176 ;
    wire signal_21177 ;
    wire signal_21178 ;
    wire signal_21179 ;
    wire signal_21180 ;
    wire signal_21181 ;
    wire signal_21182 ;
    wire signal_21183 ;
    wire signal_21184 ;
    wire signal_21185 ;
    wire signal_21186 ;
    wire signal_21187 ;
    wire signal_21188 ;
    wire signal_21189 ;
    wire signal_21190 ;
    wire signal_21191 ;
    wire signal_21192 ;
    wire signal_21193 ;
    wire signal_21194 ;
    wire signal_21195 ;
    wire signal_21196 ;
    wire signal_21197 ;
    wire signal_21198 ;
    wire signal_21199 ;
    wire signal_21200 ;
    wire signal_21201 ;
    wire signal_21202 ;
    wire signal_21203 ;
    wire signal_21204 ;
    wire signal_21205 ;
    wire signal_21206 ;
    wire signal_21207 ;
    wire signal_21208 ;
    wire signal_21209 ;
    wire signal_21210 ;
    wire signal_21211 ;
    wire signal_21212 ;
    wire signal_21213 ;
    wire signal_21214 ;
    wire signal_21215 ;
    wire signal_21216 ;
    wire signal_21217 ;
    wire signal_21218 ;
    wire signal_21219 ;
    wire signal_21220 ;
    wire signal_21221 ;
    wire signal_21222 ;
    wire signal_21223 ;
    wire signal_21224 ;
    wire signal_21225 ;
    wire signal_21226 ;
    wire signal_21227 ;
    wire signal_21228 ;
    wire signal_21229 ;
    wire signal_21230 ;
    wire signal_21231 ;
    wire signal_21232 ;
    wire signal_21233 ;
    wire signal_21234 ;
    wire signal_21235 ;
    wire signal_21236 ;
    wire signal_21237 ;
    wire signal_21238 ;
    wire signal_21239 ;
    wire signal_21240 ;
    wire signal_21241 ;
    wire signal_21242 ;
    wire signal_21243 ;
    wire signal_21244 ;
    wire signal_21245 ;
    wire signal_21246 ;
    wire signal_21247 ;
    wire signal_21248 ;
    wire signal_21249 ;
    wire signal_21250 ;
    wire signal_21251 ;
    wire signal_21252 ;
    wire signal_21253 ;
    wire signal_21254 ;
    wire signal_21255 ;
    wire signal_21256 ;
    wire signal_21257 ;
    wire signal_21258 ;
    wire signal_21259 ;
    wire signal_21260 ;
    wire signal_21261 ;
    wire signal_21262 ;
    wire signal_21263 ;
    wire signal_21264 ;
    wire signal_21265 ;
    wire signal_21266 ;
    wire signal_21267 ;
    wire signal_21268 ;
    wire signal_21269 ;
    wire signal_21270 ;
    wire signal_21271 ;
    wire signal_21272 ;
    wire signal_21273 ;
    wire signal_21274 ;
    wire signal_21275 ;
    wire signal_21276 ;
    wire signal_21277 ;
    wire signal_21278 ;
    wire signal_21279 ;
    wire signal_21280 ;
    wire signal_21281 ;
    wire signal_21282 ;
    wire signal_21283 ;
    wire signal_21284 ;
    wire signal_21285 ;
    wire signal_21286 ;
    wire signal_21287 ;
    wire signal_21288 ;
    wire signal_21289 ;
    wire signal_21290 ;
    wire signal_21291 ;
    wire signal_21292 ;
    wire signal_21293 ;
    wire signal_21294 ;
    wire signal_21295 ;
    wire signal_21296 ;
    wire signal_21297 ;
    wire signal_21298 ;
    wire signal_21299 ;
    wire signal_21300 ;
    wire signal_21301 ;
    wire signal_21302 ;
    wire signal_21303 ;
    wire signal_21304 ;
    wire signal_21305 ;
    wire signal_21306 ;
    wire signal_21307 ;
    wire signal_21308 ;
    wire signal_21309 ;
    wire signal_21310 ;
    wire signal_21311 ;
    wire signal_21312 ;
    wire signal_21313 ;
    wire signal_21314 ;
    wire signal_21315 ;
    wire signal_21316 ;
    wire signal_21317 ;
    wire signal_21318 ;
    wire signal_21319 ;
    wire signal_21320 ;
    wire signal_21321 ;
    wire signal_21322 ;
    wire signal_21323 ;
    wire signal_21324 ;
    wire signal_21325 ;
    wire signal_21326 ;
    wire signal_21327 ;
    wire signal_21328 ;
    wire signal_21329 ;
    wire signal_21330 ;
    wire signal_21331 ;
    wire signal_21332 ;
    wire signal_21333 ;
    wire signal_21334 ;
    wire signal_21335 ;
    wire signal_21336 ;
    wire signal_21337 ;
    wire signal_21338 ;
    wire signal_21339 ;
    wire signal_21340 ;
    wire signal_21341 ;
    wire signal_21342 ;
    wire signal_21343 ;
    wire signal_21344 ;
    wire signal_21345 ;
    wire signal_21346 ;
    wire signal_21347 ;
    wire signal_21348 ;
    wire signal_21349 ;
    wire signal_21350 ;
    wire signal_21351 ;
    wire signal_21352 ;
    wire signal_21353 ;
    wire signal_21354 ;
    wire signal_21355 ;
    wire signal_21356 ;
    wire signal_21357 ;
    wire signal_21358 ;
    wire signal_21359 ;
    wire signal_21360 ;
    wire signal_21361 ;
    wire signal_21362 ;
    wire signal_21363 ;
    wire signal_21364 ;
    wire signal_21365 ;
    wire signal_21366 ;
    wire signal_21367 ;
    wire signal_21368 ;
    wire signal_21369 ;
    wire signal_21370 ;
    wire signal_21371 ;
    wire signal_21372 ;
    wire signal_21373 ;
    wire signal_21374 ;
    wire signal_21375 ;
    wire signal_21376 ;
    wire signal_21377 ;
    wire signal_21378 ;
    wire signal_21379 ;
    wire signal_21380 ;
    wire signal_21381 ;
    wire signal_21382 ;
    wire signal_21383 ;
    wire signal_21384 ;
    wire signal_21385 ;
    wire signal_21386 ;
    wire signal_21387 ;
    wire signal_21388 ;
    wire signal_21389 ;
    wire signal_21390 ;
    wire signal_21391 ;
    wire signal_21392 ;
    wire signal_21393 ;
    wire signal_21394 ;
    wire signal_21395 ;
    wire signal_21396 ;
    wire signal_21397 ;
    wire signal_21398 ;
    wire signal_21399 ;
    wire signal_21400 ;
    wire signal_21401 ;
    wire signal_21402 ;
    wire signal_21403 ;
    wire signal_21404 ;
    wire signal_21405 ;
    wire signal_21406 ;
    wire signal_21407 ;
    wire signal_21408 ;
    wire signal_21409 ;
    wire signal_21410 ;
    wire signal_21411 ;
    wire signal_21412 ;
    wire signal_21413 ;
    wire signal_21414 ;
    wire signal_21415 ;
    wire signal_21416 ;
    wire signal_21417 ;
    wire signal_21418 ;
    wire signal_21419 ;
    wire signal_21420 ;
    wire signal_21421 ;
    wire signal_21422 ;
    wire signal_21423 ;
    wire signal_21424 ;
    wire signal_21425 ;
    wire signal_21426 ;
    wire signal_21427 ;
    wire signal_21428 ;
    wire signal_21429 ;
    wire signal_21430 ;
    wire signal_21431 ;
    wire signal_21432 ;
    wire signal_21433 ;
    wire signal_21434 ;
    wire signal_21435 ;
    wire signal_21436 ;
    wire signal_21437 ;
    wire signal_21438 ;
    wire signal_21439 ;
    wire signal_21440 ;
    wire signal_21441 ;
    wire signal_21442 ;
    wire signal_21443 ;
    wire signal_21444 ;
    wire signal_21445 ;
    wire signal_21446 ;
    wire signal_21447 ;
    wire signal_21448 ;
    wire signal_21449 ;
    wire signal_21450 ;
    wire signal_21451 ;
    wire signal_21452 ;
    wire signal_21453 ;
    wire signal_21454 ;
    wire signal_21455 ;
    wire signal_21456 ;
    wire signal_21457 ;
    wire signal_21458 ;
    wire signal_21459 ;
    wire signal_21460 ;
    wire signal_21461 ;
    wire signal_21462 ;
    wire signal_21463 ;
    wire signal_21464 ;
    wire signal_21465 ;
    wire signal_21466 ;
    wire signal_21467 ;
    wire signal_21468 ;
    wire signal_21469 ;
    wire signal_21470 ;
    wire signal_21471 ;
    wire signal_21472 ;
    wire signal_21473 ;
    wire signal_21474 ;
    wire signal_21475 ;
    wire signal_21476 ;
    wire signal_21477 ;
    wire signal_21478 ;
    wire signal_21479 ;
    wire signal_21480 ;
    wire signal_21481 ;
    wire signal_21482 ;
    wire signal_21483 ;
    wire signal_21484 ;
    wire signal_21485 ;
    wire signal_21486 ;
    wire signal_21487 ;
    wire signal_21488 ;
    wire signal_21489 ;
    wire signal_21490 ;
    wire signal_21491 ;
    wire signal_21492 ;
    wire signal_21493 ;
    wire signal_21494 ;
    wire signal_21495 ;
    wire signal_21496 ;
    wire signal_21497 ;
    wire signal_21498 ;
    wire signal_21499 ;
    wire signal_21500 ;
    wire signal_21501 ;
    wire signal_21502 ;
    wire signal_21503 ;
    wire signal_21504 ;
    wire signal_21505 ;
    wire signal_21506 ;
    wire signal_21507 ;
    wire signal_21508 ;
    wire signal_21509 ;
    wire signal_21510 ;
    wire signal_21511 ;
    wire signal_21512 ;
    wire signal_21513 ;
    wire signal_21514 ;
    wire signal_21515 ;
    wire signal_21516 ;
    wire signal_21517 ;
    wire signal_21518 ;
    wire signal_21519 ;
    wire signal_21520 ;
    wire signal_21521 ;
    wire signal_21522 ;
    wire signal_21523 ;
    wire signal_21524 ;
    wire signal_21525 ;
    wire signal_21526 ;
    wire signal_21527 ;
    wire signal_21528 ;
    wire signal_21529 ;
    wire signal_21530 ;
    wire signal_21531 ;
    wire signal_21532 ;
    wire signal_21533 ;
    wire signal_21534 ;
    wire signal_21535 ;
    wire signal_21536 ;
    wire signal_21537 ;
    wire signal_21538 ;
    wire signal_21539 ;
    wire signal_21540 ;
    wire signal_21541 ;
    wire signal_21542 ;
    wire signal_21543 ;
    wire signal_21544 ;
    wire signal_21545 ;
    wire signal_21546 ;
    wire signal_21547 ;
    wire signal_21548 ;
    wire signal_21549 ;
    wire signal_21550 ;
    wire signal_21551 ;
    wire signal_21552 ;
    wire signal_21553 ;
    wire signal_21554 ;
    wire signal_21555 ;
    wire signal_21556 ;
    wire signal_21557 ;
    wire signal_21558 ;
    wire signal_21559 ;
    wire signal_21560 ;
    wire signal_21561 ;
    wire signal_21562 ;
    wire signal_21563 ;
    wire signal_21564 ;
    wire signal_21565 ;
    wire signal_21566 ;
    wire signal_21567 ;
    wire signal_21568 ;
    wire signal_21569 ;
    wire signal_21570 ;
    wire signal_21571 ;
    wire signal_21572 ;
    wire signal_21573 ;
    wire signal_21574 ;
    wire signal_21575 ;
    wire signal_21576 ;
    wire signal_21577 ;
    wire signal_21578 ;
    wire signal_21579 ;
    wire signal_21580 ;
    wire signal_21581 ;
    wire signal_21582 ;
    wire signal_21583 ;
    wire signal_21584 ;
    wire signal_21585 ;
    wire signal_21586 ;
    wire signal_21587 ;
    wire signal_21588 ;
    wire signal_21589 ;
    wire signal_21590 ;
    wire signal_21591 ;
    wire signal_21592 ;
    wire signal_21593 ;
    wire signal_21594 ;
    wire signal_21595 ;
    wire signal_21596 ;
    wire signal_21597 ;
    wire signal_21598 ;
    wire signal_21599 ;
    wire signal_21600 ;
    wire signal_21601 ;
    wire signal_21602 ;
    wire signal_21603 ;
    wire signal_21604 ;
    wire signal_21605 ;
    wire signal_21606 ;
    wire signal_21607 ;
    wire signal_21608 ;
    wire signal_21609 ;
    wire signal_21610 ;
    wire signal_21611 ;
    wire signal_21612 ;
    wire signal_21613 ;
    wire signal_21614 ;
    wire signal_21615 ;
    wire signal_21616 ;
    wire signal_21617 ;
    wire signal_21618 ;
    wire signal_21619 ;
    wire signal_21620 ;
    wire signal_21621 ;
    wire signal_21622 ;
    wire signal_21623 ;
    wire signal_21624 ;
    wire signal_21625 ;
    wire signal_21626 ;
    wire signal_21627 ;
    wire signal_21628 ;
    wire signal_21629 ;
    wire signal_21630 ;
    wire signal_21631 ;
    wire signal_21632 ;
    wire signal_21633 ;
    wire signal_21634 ;
    wire signal_21635 ;
    wire signal_21636 ;
    wire signal_21637 ;
    wire signal_21638 ;
    wire signal_21639 ;
    wire signal_21640 ;
    wire signal_21641 ;
    wire signal_21642 ;
    wire signal_21643 ;
    wire signal_21644 ;
    wire signal_21645 ;
    wire signal_21646 ;
    wire signal_21647 ;
    wire signal_21648 ;
    wire signal_21649 ;
    wire signal_21650 ;
    wire signal_21651 ;
    wire signal_21652 ;
    wire signal_21653 ;
    wire signal_21654 ;
    wire signal_21655 ;
    wire signal_21656 ;
    wire signal_21657 ;
    wire signal_21658 ;
    wire signal_21659 ;
    wire signal_21660 ;
    wire signal_21661 ;
    wire signal_21662 ;
    wire signal_21663 ;
    wire signal_21664 ;
    wire signal_21665 ;
    wire signal_21666 ;
    wire signal_21667 ;
    wire signal_21668 ;
    wire signal_21669 ;
    wire signal_21670 ;
    wire signal_21671 ;
    wire signal_21672 ;
    wire signal_21673 ;
    wire signal_21674 ;
    wire signal_21675 ;
    wire signal_21676 ;
    wire signal_21677 ;
    wire signal_21678 ;
    wire signal_21679 ;
    wire signal_21680 ;
    wire signal_21681 ;
    wire signal_21682 ;
    wire signal_21683 ;
    wire signal_21684 ;
    wire signal_21685 ;
    wire signal_21686 ;
    wire signal_21687 ;
    wire signal_21688 ;
    wire signal_21689 ;
    wire signal_21690 ;
    wire signal_21691 ;
    wire signal_21692 ;
    wire signal_21693 ;
    wire signal_21694 ;
    wire signal_21695 ;
    wire signal_21696 ;
    wire signal_21697 ;
    wire signal_21698 ;
    wire signal_21699 ;
    wire signal_21700 ;
    wire signal_21701 ;
    wire signal_21702 ;
    wire signal_21703 ;
    wire signal_21704 ;
    wire signal_21705 ;
    wire signal_21706 ;
    wire signal_21707 ;
    wire signal_21708 ;
    wire signal_21709 ;
    wire signal_21710 ;
    wire signal_21711 ;
    wire signal_21712 ;
    wire signal_21713 ;
    wire signal_21714 ;
    wire signal_21715 ;
    wire signal_21716 ;
    wire signal_21717 ;
    wire signal_21718 ;
    wire signal_21719 ;
    wire signal_21720 ;
    wire signal_21721 ;
    wire signal_21722 ;
    wire signal_21723 ;
    wire signal_21724 ;
    wire signal_21725 ;
    wire signal_21726 ;
    wire signal_21727 ;
    wire signal_21728 ;
    wire signal_21729 ;
    wire signal_21730 ;
    wire signal_21731 ;
    wire signal_21732 ;
    wire signal_21733 ;
    wire signal_21734 ;
    wire signal_21735 ;
    wire signal_21736 ;
    wire signal_21737 ;
    wire signal_21738 ;
    wire signal_21739 ;
    wire signal_21740 ;
    wire signal_21741 ;
    wire signal_21742 ;
    wire signal_21743 ;
    wire signal_21744 ;
    wire signal_21745 ;
    wire signal_21746 ;
    wire signal_21747 ;
    wire signal_21748 ;
    wire signal_21749 ;
    wire signal_21750 ;
    wire signal_21751 ;
    wire signal_21752 ;
    wire signal_21753 ;
    wire signal_21754 ;
    wire signal_21755 ;
    wire signal_21756 ;
    wire signal_21757 ;
    wire signal_21758 ;
    wire signal_21759 ;
    wire signal_21760 ;
    wire signal_21761 ;
    wire signal_21762 ;
    wire signal_21763 ;
    wire signal_21764 ;
    wire signal_21765 ;
    wire signal_21766 ;
    wire signal_21767 ;
    wire signal_21768 ;
    wire signal_21769 ;
    wire signal_21770 ;
    wire signal_21771 ;
    wire signal_21772 ;
    wire signal_21773 ;
    wire signal_21774 ;
    wire signal_21775 ;
    wire signal_21776 ;
    wire signal_21777 ;
    wire signal_21778 ;
    wire signal_21779 ;
    wire signal_21780 ;
    wire signal_21781 ;
    wire signal_21782 ;
    wire signal_21783 ;
    wire signal_21784 ;
    wire signal_21785 ;
    wire signal_21786 ;
    wire signal_21787 ;
    wire signal_21788 ;
    wire signal_21789 ;
    wire signal_21790 ;
    wire signal_21791 ;
    wire signal_21792 ;
    wire signal_21793 ;
    wire signal_21794 ;
    wire signal_21795 ;
    wire signal_21796 ;
    wire signal_21797 ;
    wire signal_21798 ;
    wire signal_21799 ;
    wire signal_21800 ;
    wire signal_21801 ;
    wire signal_21802 ;
    wire signal_21803 ;
    wire signal_21804 ;
    wire signal_21805 ;
    wire signal_21806 ;
    wire signal_21807 ;
    wire signal_21808 ;
    wire signal_21809 ;
    wire signal_21810 ;
    wire signal_21811 ;
    wire signal_21812 ;
    wire signal_21813 ;
    wire signal_21814 ;
    wire signal_21815 ;
    wire signal_21816 ;
    wire signal_21817 ;
    wire signal_21818 ;
    wire signal_21819 ;
    wire signal_21820 ;
    wire signal_21821 ;
    wire signal_21822 ;
    wire signal_21823 ;
    wire signal_21824 ;
    wire signal_21825 ;
    wire signal_21826 ;
    wire signal_21827 ;
    wire signal_21828 ;
    wire signal_21829 ;
    wire signal_21830 ;
    wire signal_21831 ;
    wire signal_21832 ;
    wire signal_21833 ;
    wire signal_21834 ;
    wire signal_21835 ;
    wire signal_21836 ;
    wire signal_21837 ;
    wire signal_21838 ;
    wire signal_21839 ;
    wire signal_21840 ;
    wire signal_21841 ;
    wire signal_21842 ;
    wire signal_21843 ;
    wire signal_21844 ;
    wire signal_21845 ;
    wire signal_21846 ;
    wire signal_21847 ;
    wire signal_21848 ;
    wire signal_21849 ;
    wire signal_21850 ;
    wire signal_21851 ;
    wire signal_21852 ;
    wire signal_21853 ;
    wire signal_21854 ;
    wire signal_21855 ;
    wire signal_21856 ;
    wire signal_21857 ;
    wire signal_21858 ;
    wire signal_21859 ;
    wire signal_21860 ;
    wire signal_21861 ;
    wire signal_21862 ;
    wire signal_21863 ;
    wire signal_21864 ;
    wire signal_21865 ;
    wire signal_21866 ;
    wire signal_21867 ;
    wire signal_21868 ;
    wire signal_21869 ;
    wire signal_21870 ;
    wire signal_21871 ;
    wire signal_21872 ;
    wire signal_21873 ;
    wire signal_21874 ;
    wire signal_21875 ;
    wire signal_21876 ;
    wire signal_21877 ;
    wire signal_21878 ;
    wire signal_21879 ;
    wire signal_21880 ;
    wire signal_21881 ;
    wire signal_21882 ;
    wire signal_21883 ;
    wire signal_21884 ;
    wire signal_21885 ;
    wire signal_21886 ;
    wire signal_21887 ;
    wire signal_21888 ;
    wire signal_21889 ;
    wire signal_21890 ;
    wire signal_21891 ;
    wire signal_21892 ;
    wire signal_21893 ;
    wire signal_21894 ;
    wire signal_21895 ;
    wire signal_21896 ;
    wire signal_21897 ;
    wire signal_21898 ;
    wire signal_21899 ;
    wire signal_21900 ;
    wire signal_21901 ;
    wire signal_21902 ;
    wire signal_21903 ;
    wire signal_21904 ;
    wire signal_21905 ;
    wire signal_21906 ;
    wire signal_21907 ;
    wire signal_21908 ;
    wire signal_21909 ;
    wire signal_21910 ;
    wire signal_21911 ;
    wire signal_21912 ;
    wire signal_21913 ;
    wire signal_21914 ;
    wire signal_21915 ;
    wire signal_21916 ;
    wire signal_21917 ;
    wire signal_21918 ;
    wire signal_21919 ;
    wire signal_21920 ;
    wire signal_21921 ;
    wire signal_21922 ;
    wire signal_21923 ;
    wire signal_21924 ;
    wire signal_21925 ;
    wire signal_21926 ;
    wire signal_21927 ;
    wire signal_21928 ;
    wire signal_21929 ;
    wire signal_21930 ;
    wire signal_21931 ;
    wire signal_21932 ;
    wire signal_21933 ;
    wire signal_21934 ;
    wire signal_21935 ;
    wire signal_21936 ;
    wire signal_21937 ;
    wire signal_21938 ;
    wire signal_21939 ;
    wire signal_21940 ;
    wire signal_21941 ;
    wire signal_21942 ;
    wire signal_21943 ;
    wire signal_21944 ;
    wire signal_21945 ;
    wire signal_21946 ;
    wire signal_21947 ;
    wire signal_21948 ;
    wire signal_21949 ;
    wire signal_21950 ;
    wire signal_21951 ;
    wire signal_21952 ;
    wire signal_21953 ;
    wire signal_21954 ;
    wire signal_21955 ;
    wire signal_21956 ;
    wire signal_21957 ;
    wire signal_21958 ;
    wire signal_21959 ;
    wire signal_21960 ;
    wire signal_21961 ;
    wire signal_21962 ;
    wire signal_21963 ;
    wire signal_21964 ;
    wire signal_21965 ;
    wire signal_21966 ;
    wire signal_21967 ;
    wire signal_21968 ;
    wire signal_21969 ;
    wire signal_21970 ;
    wire signal_21971 ;
    wire signal_21972 ;
    wire signal_21973 ;
    wire signal_21974 ;
    wire signal_21975 ;
    wire signal_21976 ;
    wire signal_21977 ;
    wire signal_21978 ;
    wire signal_21979 ;
    wire signal_21980 ;
    wire signal_21981 ;
    wire signal_21982 ;
    wire signal_21983 ;
    wire signal_21984 ;
    wire signal_21985 ;
    wire signal_21986 ;
    wire signal_21987 ;
    wire signal_21988 ;
    wire signal_21989 ;
    wire signal_21990 ;
    wire signal_21991 ;
    wire signal_21992 ;
    wire signal_21993 ;
    wire signal_21994 ;
    wire signal_21995 ;
    wire signal_21996 ;
    wire signal_21997 ;
    wire signal_21998 ;
    wire signal_21999 ;
    wire signal_22000 ;
    wire signal_22001 ;
    wire signal_22002 ;
    wire signal_22003 ;
    wire signal_22004 ;
    wire signal_22005 ;
    wire signal_22006 ;
    wire signal_22007 ;
    wire signal_22008 ;
    wire signal_22009 ;
    wire signal_22010 ;
    wire signal_22011 ;
    wire signal_22012 ;
    wire signal_22013 ;
    wire signal_22014 ;
    wire signal_22015 ;
    wire signal_22016 ;
    wire signal_22017 ;
    wire signal_22018 ;
    wire signal_22019 ;
    wire signal_22020 ;
    wire signal_22021 ;
    wire signal_22022 ;
    wire signal_22023 ;
    wire signal_22024 ;
    wire signal_22025 ;
    wire signal_22026 ;
    wire signal_22027 ;
    wire signal_22028 ;
    wire signal_22029 ;
    wire signal_22030 ;
    wire signal_22031 ;
    wire signal_22032 ;
    wire signal_22033 ;
    wire signal_22034 ;
    wire signal_22035 ;
    wire signal_22036 ;
    wire signal_22037 ;
    wire signal_22038 ;
    wire signal_22039 ;
    wire signal_22040 ;
    wire signal_22041 ;
    wire signal_22042 ;
    wire signal_22043 ;
    wire signal_22044 ;
    wire signal_22045 ;
    wire signal_22046 ;
    wire signal_22047 ;
    wire signal_22048 ;
    wire signal_22049 ;
    wire signal_22050 ;
    wire signal_22051 ;
    wire signal_22052 ;
    wire signal_22053 ;
    wire signal_22054 ;
    wire signal_22055 ;
    wire signal_22056 ;
    wire signal_22057 ;
    wire signal_22058 ;
    wire signal_22059 ;
    wire signal_22060 ;
    wire signal_22061 ;
    wire signal_22062 ;
    wire signal_22063 ;
    wire signal_22064 ;
    wire signal_22065 ;
    wire signal_22066 ;
    wire signal_22067 ;
    wire signal_22068 ;
    wire signal_22069 ;
    wire signal_22070 ;
    wire signal_22071 ;
    wire signal_22072 ;
    wire signal_22073 ;
    wire signal_22074 ;
    wire signal_22075 ;
    wire signal_22076 ;
    wire signal_22077 ;
    wire signal_22078 ;
    wire signal_22079 ;
    wire signal_22080 ;
    wire signal_22081 ;
    wire signal_22082 ;
    wire signal_22083 ;
    wire signal_22084 ;
    wire signal_22085 ;
    wire signal_22086 ;
    wire signal_22087 ;
    wire signal_22088 ;
    wire signal_22089 ;
    wire signal_22090 ;
    wire signal_22091 ;
    wire signal_22092 ;
    wire signal_22093 ;
    wire signal_22094 ;
    wire signal_22095 ;
    wire signal_22096 ;
    wire signal_22097 ;
    wire signal_22098 ;
    wire signal_22099 ;
    wire signal_22100 ;
    wire signal_22101 ;
    wire signal_22102 ;
    wire signal_22103 ;
    wire signal_22104 ;
    wire signal_22105 ;
    wire signal_22106 ;
    wire signal_22107 ;
    wire signal_22108 ;
    wire signal_22109 ;
    wire signal_22110 ;
    wire signal_22111 ;
    wire signal_22112 ;
    wire signal_22113 ;
    wire signal_22114 ;
    wire signal_22115 ;
    wire signal_22116 ;
    wire signal_22117 ;
    wire signal_22118 ;
    wire signal_22119 ;
    wire signal_22120 ;
    wire signal_22121 ;
    wire signal_22122 ;
    wire signal_22123 ;
    wire signal_22124 ;
    wire signal_22125 ;
    wire signal_22126 ;
    wire signal_22127 ;
    wire signal_22128 ;
    wire signal_22129 ;
    wire signal_22130 ;
    wire signal_22131 ;
    wire signal_22132 ;
    wire signal_22133 ;
    wire signal_22134 ;
    wire signal_22135 ;
    wire signal_22136 ;
    wire signal_22137 ;
    wire signal_22138 ;
    wire signal_22139 ;
    wire signal_22140 ;
    wire signal_22141 ;
    wire signal_22142 ;
    wire signal_22143 ;
    wire signal_22144 ;
    wire signal_22145 ;
    wire signal_22146 ;
    wire signal_22147 ;
    wire signal_22148 ;
    wire signal_22149 ;
    wire signal_22150 ;
    wire signal_22151 ;
    wire signal_22152 ;
    wire signal_22153 ;
    wire signal_22154 ;
    wire signal_22155 ;
    wire signal_22156 ;
    wire signal_22157 ;
    wire signal_22158 ;
    wire signal_22159 ;
    wire signal_22160 ;
    wire signal_22161 ;
    wire signal_22162 ;
    wire signal_22163 ;
    wire signal_22164 ;
    wire signal_22165 ;
    wire signal_22166 ;
    wire signal_22167 ;
    wire signal_22168 ;
    wire signal_22169 ;
    wire signal_22170 ;
    wire signal_22171 ;
    wire signal_22172 ;
    wire signal_22173 ;
    wire signal_22174 ;
    wire signal_22175 ;
    wire signal_22176 ;
    wire signal_22177 ;
    wire signal_22178 ;
    wire signal_22179 ;
    wire signal_22180 ;
    wire signal_22181 ;
    wire signal_22182 ;
    wire signal_22183 ;
    wire signal_22184 ;
    wire signal_22185 ;
    wire signal_22186 ;
    wire signal_22187 ;
    wire signal_22188 ;
    wire signal_22189 ;
    wire signal_22190 ;
    wire signal_22191 ;
    wire signal_22192 ;
    wire signal_22193 ;
    wire signal_22194 ;
    wire signal_22195 ;
    wire signal_22196 ;
    wire signal_22197 ;
    wire signal_22198 ;
    wire signal_22199 ;
    wire signal_22200 ;
    wire signal_22201 ;
    wire signal_22202 ;
    wire signal_22203 ;
    wire signal_22204 ;
    wire signal_22205 ;
    wire signal_22206 ;
    wire signal_22207 ;
    wire signal_22208 ;
    wire signal_22209 ;
    wire signal_22210 ;
    wire signal_22211 ;
    wire signal_22212 ;
    wire signal_22213 ;
    wire signal_22214 ;
    wire signal_22215 ;
    wire signal_22216 ;
    wire signal_22217 ;
    wire signal_22218 ;
    wire signal_22219 ;
    wire signal_22220 ;
    wire signal_22221 ;
    wire signal_22222 ;
    wire signal_22223 ;
    wire signal_22224 ;
    wire signal_22225 ;
    wire signal_22226 ;
    wire signal_22227 ;
    wire signal_22228 ;
    wire signal_22229 ;
    wire signal_22230 ;
    wire signal_22231 ;
    wire signal_22232 ;
    wire signal_22233 ;
    wire signal_22234 ;
    wire signal_22235 ;
    wire signal_22236 ;
    wire signal_22237 ;
    wire signal_22238 ;
    wire signal_22239 ;
    wire signal_22240 ;
    wire signal_22241 ;
    wire signal_22242 ;
    wire signal_22243 ;
    wire signal_22244 ;
    wire signal_22245 ;
    wire signal_22246 ;
    wire signal_22247 ;
    wire signal_22248 ;
    wire signal_22249 ;
    wire signal_22250 ;
    wire signal_22251 ;
    wire signal_22252 ;
    wire signal_22253 ;
    wire signal_22254 ;
    wire signal_22255 ;
    wire signal_22256 ;
    wire signal_22257 ;
    wire signal_22258 ;
    wire signal_22259 ;
    wire signal_22260 ;
    wire signal_22261 ;
    wire signal_22262 ;
    wire signal_22263 ;
    wire signal_22264 ;
    wire signal_22265 ;
    wire signal_22266 ;
    wire signal_22267 ;
    wire signal_22268 ;
    wire signal_22269 ;
    wire signal_22270 ;
    wire signal_22271 ;
    wire signal_22272 ;
    wire signal_22273 ;
    wire signal_22274 ;
    wire signal_22275 ;
    wire signal_22276 ;
    wire signal_22277 ;
    wire signal_22278 ;
    wire signal_22279 ;
    wire signal_22280 ;
    wire signal_22281 ;
    wire signal_22282 ;
    wire signal_22283 ;
    wire signal_22284 ;
    wire signal_22285 ;
    wire signal_22286 ;
    wire signal_22287 ;
    wire signal_22288 ;
    wire signal_22289 ;
    wire signal_22290 ;
    wire signal_22291 ;
    wire signal_22292 ;
    wire signal_22293 ;
    wire signal_22294 ;
    wire signal_22295 ;
    wire signal_22296 ;
    wire signal_22297 ;
    wire signal_22298 ;
    wire signal_22299 ;
    wire signal_22300 ;
    wire signal_22301 ;
    wire signal_22302 ;
    wire signal_22303 ;
    wire signal_22304 ;
    wire signal_22305 ;
    wire signal_22306 ;
    wire signal_22307 ;
    wire signal_22308 ;
    wire signal_22309 ;
    wire signal_22310 ;
    wire signal_22311 ;
    wire signal_22312 ;
    wire signal_22313 ;
    wire signal_22314 ;
    wire signal_22315 ;
    wire signal_22316 ;
    wire signal_22317 ;
    wire signal_22318 ;
    wire signal_22319 ;
    wire signal_22320 ;
    wire signal_22321 ;
    wire signal_22322 ;
    wire signal_22323 ;
    wire signal_22324 ;
    wire signal_22325 ;
    wire signal_22326 ;
    wire signal_22327 ;
    wire signal_22328 ;
    wire signal_22329 ;
    wire signal_22330 ;
    wire signal_22331 ;
    wire signal_22332 ;
    wire signal_22333 ;
    wire signal_22334 ;
    wire signal_22335 ;
    wire signal_22336 ;
    wire signal_22337 ;
    wire signal_22338 ;
    wire signal_22339 ;
    wire signal_22340 ;
    wire signal_22341 ;
    wire signal_22342 ;
    wire signal_22343 ;
    wire signal_22344 ;
    wire signal_22345 ;
    wire signal_22346 ;
    wire signal_22347 ;
    wire signal_22348 ;
    wire signal_22349 ;
    wire signal_22350 ;
    wire signal_22351 ;
    wire signal_22352 ;
    wire signal_22353 ;
    wire signal_22354 ;
    wire signal_22355 ;
    wire signal_22356 ;
    wire signal_22357 ;
    wire signal_22358 ;
    wire signal_22359 ;
    wire signal_22360 ;
    wire signal_22361 ;
    wire signal_22362 ;
    wire signal_22363 ;
    wire signal_22364 ;
    wire signal_22365 ;
    wire signal_22366 ;
    wire signal_22367 ;
    wire signal_22368 ;
    wire signal_22369 ;
    wire signal_22370 ;
    wire signal_22371 ;
    wire signal_22372 ;
    wire signal_22373 ;
    wire signal_22374 ;
    wire signal_22375 ;
    wire signal_22376 ;
    wire signal_22377 ;
    wire signal_22378 ;
    wire signal_22379 ;
    wire signal_22380 ;
    wire signal_22381 ;
    wire signal_22382 ;
    wire signal_22383 ;
    wire signal_22384 ;
    wire signal_22385 ;
    wire signal_22386 ;
    wire signal_22387 ;
    wire signal_22388 ;
    wire signal_22389 ;
    wire signal_22390 ;
    wire signal_22391 ;
    wire signal_22392 ;
    wire signal_22393 ;
    wire signal_22394 ;
    wire signal_22395 ;
    wire signal_22396 ;
    wire signal_22397 ;
    wire signal_22398 ;
    wire signal_22399 ;
    wire signal_22400 ;
    wire signal_22401 ;
    wire signal_22402 ;
    wire signal_22403 ;
    wire signal_22404 ;
    wire signal_22405 ;
    wire signal_22406 ;
    wire signal_22407 ;
    wire signal_22408 ;
    wire signal_22409 ;
    wire signal_22410 ;
    wire signal_22411 ;
    wire signal_22412 ;
    wire signal_22413 ;
    wire signal_22414 ;
    wire signal_22415 ;
    wire signal_22416 ;
    wire signal_22417 ;
    wire signal_22418 ;
    wire signal_22419 ;
    wire signal_22420 ;
    wire signal_22421 ;
    wire signal_22422 ;
    wire signal_22423 ;
    wire signal_22424 ;
    wire signal_22425 ;
    wire signal_22426 ;
    wire signal_22427 ;
    wire signal_22428 ;
    wire signal_22429 ;
    wire signal_22430 ;
    wire signal_22431 ;
    wire signal_22432 ;
    wire signal_22433 ;
    wire signal_22434 ;
    wire signal_22435 ;
    wire signal_22436 ;
    wire signal_22437 ;
    wire signal_22438 ;
    wire signal_22439 ;
    wire signal_22440 ;
    wire signal_22441 ;
    wire signal_22442 ;
    wire signal_22443 ;
    wire signal_22444 ;
    wire signal_22445 ;
    wire signal_22446 ;
    wire signal_22447 ;
    wire signal_22448 ;
    wire signal_22449 ;
    wire signal_22450 ;
    wire signal_22451 ;
    wire signal_22452 ;
    wire signal_22453 ;
    wire signal_22454 ;
    wire signal_22455 ;
    wire signal_22456 ;
    wire signal_22457 ;
    wire signal_22458 ;
    wire signal_22459 ;
    wire signal_22460 ;
    wire signal_22461 ;
    wire signal_22462 ;
    wire signal_22463 ;
    wire signal_22464 ;
    wire signal_22465 ;
    wire signal_22466 ;
    wire signal_22467 ;
    wire signal_22468 ;
    wire signal_22469 ;
    wire signal_22470 ;
    wire signal_22471 ;
    wire signal_22472 ;
    wire signal_22473 ;
    wire signal_22474 ;
    wire signal_22475 ;
    wire signal_22476 ;
    wire signal_22477 ;
    wire signal_22478 ;
    wire signal_22479 ;
    wire signal_22480 ;
    wire signal_22481 ;
    wire signal_22482 ;
    wire signal_22483 ;
    wire signal_22484 ;
    wire signal_22485 ;
    wire signal_22486 ;
    wire signal_22487 ;
    wire signal_22488 ;
    wire signal_22489 ;
    wire signal_22490 ;
    wire signal_22491 ;
    wire signal_22492 ;
    wire signal_22493 ;
    wire signal_22494 ;
    wire signal_22495 ;
    wire signal_22496 ;
    wire signal_22497 ;
    wire signal_22498 ;
    wire signal_22499 ;
    wire signal_22500 ;
    wire signal_22501 ;
    wire signal_22502 ;
    wire signal_22503 ;
    wire signal_22504 ;
    wire signal_22505 ;
    wire signal_22506 ;
    wire signal_22507 ;
    wire signal_22508 ;
    wire signal_22509 ;
    wire signal_22510 ;
    wire signal_22511 ;
    wire signal_22512 ;
    wire signal_22513 ;
    wire signal_22514 ;
    wire signal_22515 ;
    wire signal_22516 ;
    wire signal_22517 ;
    wire signal_22518 ;
    wire signal_22519 ;
    wire signal_22520 ;
    wire signal_22521 ;
    wire signal_22522 ;
    wire signal_22523 ;
    wire signal_22524 ;
    wire signal_22525 ;
    wire signal_22526 ;
    wire signal_22527 ;
    wire signal_22528 ;
    wire signal_22529 ;
    wire signal_22530 ;
    wire signal_22531 ;
    wire signal_22532 ;
    wire signal_22533 ;
    wire signal_22534 ;
    wire signal_22535 ;
    wire signal_22536 ;
    wire signal_22537 ;
    wire signal_22538 ;
    wire signal_22539 ;
    wire signal_22540 ;
    wire signal_22541 ;
    wire signal_22542 ;
    wire signal_22543 ;
    wire signal_22544 ;
    wire signal_22545 ;
    wire signal_22546 ;
    wire signal_22547 ;
    wire signal_22548 ;
    wire signal_22549 ;
    wire signal_22550 ;
    wire signal_22551 ;
    wire signal_22552 ;
    wire signal_22553 ;
    wire signal_22554 ;
    wire signal_22555 ;
    wire signal_22556 ;
    wire signal_22557 ;
    wire signal_22558 ;
    wire signal_22559 ;
    wire signal_22560 ;
    wire signal_22561 ;
    wire signal_22562 ;
    wire signal_22563 ;
    wire signal_22564 ;
    wire signal_22565 ;
    wire signal_22566 ;
    wire signal_22567 ;
    wire signal_22568 ;
    wire signal_22569 ;
    wire signal_22570 ;
    wire signal_22571 ;
    wire signal_22572 ;
    wire signal_22573 ;
    wire signal_22574 ;
    wire signal_22575 ;
    wire signal_22576 ;
    wire signal_22577 ;
    wire signal_22578 ;
    wire signal_22579 ;
    wire signal_22580 ;
    wire signal_22581 ;
    wire signal_22582 ;
    wire signal_22583 ;
    wire signal_22584 ;
    wire signal_22585 ;
    wire signal_22586 ;
    wire signal_22587 ;
    wire signal_22588 ;
    wire signal_22589 ;
    wire signal_22590 ;
    wire signal_22591 ;
    wire signal_22592 ;
    wire signal_22593 ;
    wire signal_22594 ;
    wire signal_22595 ;
    wire signal_22596 ;
    wire signal_22597 ;
    wire signal_22598 ;
    wire signal_22599 ;
    wire signal_22600 ;
    wire signal_22601 ;
    wire signal_22602 ;
    wire signal_22603 ;
    wire signal_22604 ;
    wire signal_22605 ;
    wire signal_22606 ;
    wire signal_22607 ;
    wire signal_22608 ;
    wire signal_22609 ;
    wire signal_22610 ;
    wire signal_22611 ;
    wire signal_22612 ;
    wire signal_22613 ;
    wire signal_22614 ;
    wire signal_22615 ;
    wire signal_22616 ;
    wire signal_22617 ;
    wire signal_22618 ;
    wire signal_22619 ;
    wire signal_22620 ;
    wire signal_22621 ;
    wire signal_22622 ;
    wire signal_22623 ;
    wire signal_22624 ;
    wire signal_22625 ;
    wire signal_22626 ;
    wire signal_22627 ;
    wire signal_22628 ;
    wire signal_22629 ;
    wire signal_22630 ;
    wire signal_22631 ;
    wire signal_22632 ;
    wire signal_22633 ;
    wire signal_22634 ;
    wire signal_22635 ;
    wire signal_22636 ;
    wire signal_22637 ;
    wire signal_22638 ;
    wire signal_22639 ;
    wire signal_22640 ;
    wire signal_22641 ;
    wire signal_22642 ;
    wire signal_22643 ;
    wire signal_22644 ;
    wire signal_22645 ;
    wire signal_22646 ;
    wire signal_22647 ;
    wire signal_22648 ;
    wire signal_22649 ;
    wire signal_22650 ;
    wire signal_22651 ;
    wire signal_22652 ;
    wire signal_22653 ;
    wire signal_22654 ;
    wire signal_22655 ;
    wire signal_22656 ;
    wire signal_22657 ;
    wire signal_22658 ;
    wire signal_22659 ;
    wire signal_22660 ;
    wire signal_22661 ;
    wire signal_22662 ;
    wire signal_22663 ;
    wire signal_22664 ;
    wire signal_22665 ;
    wire signal_22666 ;
    wire signal_22667 ;
    wire signal_22668 ;
    wire signal_22669 ;
    wire signal_22670 ;
    wire signal_22671 ;
    wire signal_22672 ;
    wire signal_22673 ;
    wire signal_22674 ;
    wire signal_22675 ;
    wire signal_22676 ;
    wire signal_22677 ;
    wire signal_22678 ;
    wire signal_22679 ;
    wire signal_22680 ;
    wire signal_22681 ;
    wire signal_22682 ;
    wire signal_22683 ;
    wire signal_22684 ;
    wire signal_22685 ;
    wire signal_22686 ;
    wire signal_22687 ;
    wire signal_22688 ;
    wire signal_22689 ;
    wire signal_22690 ;
    wire signal_22691 ;
    wire signal_22692 ;
    wire signal_22693 ;
    wire signal_22694 ;
    wire signal_22695 ;
    wire signal_22696 ;
    wire signal_22697 ;
    wire signal_22698 ;
    wire signal_22699 ;
    wire signal_22700 ;
    wire signal_22701 ;
    wire signal_22702 ;
    wire signal_22703 ;
    wire signal_22704 ;
    wire signal_22705 ;
    wire signal_22706 ;
    wire signal_22707 ;
    wire signal_22708 ;
    wire signal_22709 ;
    wire signal_22710 ;
    wire signal_22711 ;
    wire signal_22712 ;
    wire signal_22713 ;
    wire signal_22714 ;
    wire signal_22715 ;
    wire signal_22716 ;
    wire signal_22717 ;
    wire signal_22718 ;
    wire signal_22719 ;
    wire signal_22720 ;
    wire signal_22721 ;
    wire signal_22722 ;
    wire signal_22723 ;
    wire signal_22724 ;
    wire signal_22725 ;
    wire signal_22726 ;
    wire signal_22727 ;
    wire signal_22728 ;
    wire signal_22729 ;
    wire signal_22730 ;
    wire signal_22731 ;
    wire signal_22732 ;
    wire signal_22733 ;
    wire signal_22734 ;
    wire signal_22735 ;
    wire signal_22736 ;
    wire signal_22737 ;
    wire signal_22738 ;
    wire signal_22739 ;
    wire signal_22740 ;
    wire signal_22741 ;
    wire signal_22742 ;
    wire signal_22743 ;
    wire signal_22744 ;
    wire signal_22745 ;
    wire signal_22746 ;
    wire signal_22747 ;
    wire signal_22748 ;
    wire signal_22749 ;
    wire signal_22750 ;
    wire signal_22751 ;
    wire signal_22752 ;
    wire signal_22753 ;
    wire signal_22754 ;
    wire signal_22755 ;
    wire signal_22756 ;
    wire signal_22757 ;
    wire signal_22758 ;
    wire signal_22759 ;
    wire signal_22760 ;
    wire signal_22761 ;
    wire signal_22762 ;
    wire signal_22763 ;
    wire signal_22764 ;
    wire signal_22765 ;
    wire signal_22766 ;
    wire signal_22767 ;
    wire signal_22768 ;
    wire signal_22769 ;
    wire signal_22770 ;
    wire signal_22771 ;
    wire signal_22772 ;
    wire signal_22773 ;
    wire signal_22774 ;
    wire signal_22775 ;
    wire signal_22776 ;
    wire signal_22777 ;
    wire signal_22778 ;
    wire signal_22779 ;
    wire signal_22780 ;
    wire signal_22781 ;
    wire signal_22782 ;
    wire signal_22783 ;
    wire signal_22784 ;
    wire signal_22785 ;
    wire signal_22786 ;
    wire signal_22787 ;
    wire signal_22788 ;
    wire signal_22789 ;
    wire signal_22790 ;
    wire signal_22791 ;
    wire signal_22792 ;
    wire signal_22793 ;
    wire signal_22794 ;
    wire signal_22795 ;
    wire signal_22796 ;
    wire signal_22797 ;
    wire signal_22798 ;
    wire signal_22799 ;
    wire signal_22800 ;
    wire signal_22801 ;
    wire signal_22802 ;
    wire signal_22803 ;
    wire signal_22804 ;
    wire signal_22805 ;
    wire signal_22806 ;
    wire signal_22807 ;
    wire signal_22808 ;
    wire signal_22809 ;
    wire signal_22810 ;
    wire signal_22811 ;
    wire signal_22812 ;
    wire signal_22813 ;
    wire signal_22814 ;
    wire signal_22815 ;
    wire signal_22816 ;
    wire signal_22817 ;
    wire signal_22818 ;
    wire signal_22819 ;
    wire signal_22820 ;
    wire signal_22821 ;
    wire signal_22822 ;
    wire signal_22823 ;
    wire signal_22824 ;
    wire signal_22825 ;
    wire signal_22826 ;
    wire signal_22827 ;
    wire signal_22828 ;
    wire signal_22829 ;
    wire signal_22830 ;
    wire signal_22831 ;
    wire signal_22832 ;
    wire signal_22833 ;
    wire signal_22834 ;
    wire signal_22835 ;
    wire signal_22836 ;
    wire signal_22837 ;
    wire signal_22838 ;
    wire signal_22839 ;
    wire signal_22840 ;
    wire signal_22841 ;
    wire signal_22842 ;
    wire signal_22843 ;
    wire signal_22844 ;
    wire signal_22845 ;
    wire signal_22846 ;
    wire signal_22847 ;
    wire signal_22848 ;
    wire signal_22849 ;
    wire signal_22850 ;
    wire signal_22851 ;
    wire signal_22852 ;
    wire signal_22853 ;
    wire signal_22854 ;
    wire signal_22855 ;
    wire signal_22856 ;
    wire signal_22857 ;
    wire signal_22858 ;
    wire signal_22859 ;
    wire signal_22860 ;
    wire signal_22861 ;
    wire signal_22862 ;
    wire signal_22863 ;
    wire signal_22864 ;
    wire signal_22865 ;
    wire signal_22866 ;
    wire signal_22867 ;
    wire signal_22868 ;
    wire signal_22869 ;
    wire signal_22870 ;
    wire signal_22871 ;
    wire signal_22872 ;
    wire signal_22873 ;
    wire signal_22874 ;
    wire signal_22875 ;
    wire signal_22876 ;
    wire signal_22877 ;
    wire signal_22878 ;
    wire signal_22879 ;
    wire signal_22880 ;
    wire signal_22881 ;
    wire signal_22882 ;
    wire signal_22883 ;
    wire signal_22884 ;
    wire signal_22885 ;
    wire signal_22886 ;
    wire signal_22887 ;
    wire signal_22888 ;
    wire signal_22889 ;
    wire signal_22890 ;
    wire signal_22891 ;
    wire signal_22892 ;
    wire signal_22893 ;
    wire signal_22894 ;
    wire signal_22895 ;
    wire signal_22896 ;
    wire signal_22897 ;
    wire signal_22898 ;
    wire signal_22899 ;
    wire signal_22900 ;
    wire signal_22901 ;
    wire signal_22902 ;
    wire signal_22903 ;
    wire signal_22904 ;
    wire signal_22905 ;
    wire signal_22906 ;
    wire signal_22907 ;
    wire signal_22908 ;
    wire signal_22909 ;
    wire signal_22910 ;
    wire signal_22911 ;
    wire signal_22912 ;
    wire signal_22913 ;
    wire signal_22914 ;
    wire signal_22915 ;
    wire signal_22916 ;
    wire signal_22917 ;
    wire signal_22918 ;
    wire signal_22919 ;
    wire signal_22920 ;
    wire signal_22921 ;
    wire signal_22922 ;
    wire signal_22923 ;
    wire signal_22924 ;
    wire signal_22925 ;
    wire signal_22926 ;
    wire signal_22927 ;
    wire signal_22928 ;
    wire signal_22929 ;
    wire signal_22930 ;
    wire signal_22931 ;
    wire signal_22932 ;
    wire signal_22933 ;
    wire signal_22934 ;
    wire signal_22935 ;
    wire signal_22936 ;
    wire signal_22937 ;
    wire signal_22938 ;
    wire signal_22939 ;
    wire signal_22940 ;
    wire signal_22941 ;
    wire signal_22942 ;
    wire signal_22943 ;
    wire signal_22944 ;
    wire signal_22945 ;
    wire signal_22946 ;
    wire signal_22947 ;
    wire signal_22948 ;
    wire signal_22949 ;
    wire signal_22950 ;
    wire signal_22951 ;
    wire signal_22952 ;
    wire signal_22953 ;
    wire signal_22954 ;
    wire signal_22955 ;
    wire signal_22956 ;
    wire signal_22957 ;
    wire signal_22958 ;
    wire signal_22959 ;
    wire signal_22960 ;
    wire signal_22961 ;
    wire signal_22962 ;
    wire signal_22963 ;
    wire signal_22964 ;
    wire signal_22965 ;
    wire signal_22966 ;
    wire signal_22967 ;
    wire signal_22968 ;
    wire signal_22969 ;
    wire signal_22970 ;
    wire signal_22971 ;
    wire signal_22972 ;
    wire signal_22973 ;
    wire signal_22974 ;
    wire signal_22975 ;
    wire signal_22976 ;
    wire signal_22977 ;
    wire signal_22978 ;
    wire signal_22979 ;
    wire signal_22980 ;
    wire signal_22981 ;
    wire signal_22982 ;
    wire signal_22983 ;
    wire signal_22984 ;
    wire signal_22985 ;
    wire signal_22986 ;
    wire signal_22987 ;
    wire signal_22988 ;
    wire signal_22989 ;
    wire signal_22990 ;
    wire signal_22991 ;
    wire signal_22992 ;
    wire signal_22993 ;
    wire signal_22994 ;
    wire signal_22995 ;
    wire signal_22996 ;
    wire signal_22997 ;
    wire signal_22998 ;
    wire signal_22999 ;
    wire signal_23000 ;
    wire signal_23001 ;
    wire signal_23002 ;
    wire signal_23003 ;
    wire signal_23004 ;
    wire signal_23005 ;
    wire signal_23006 ;
    wire signal_23007 ;
    wire signal_23008 ;
    wire signal_23009 ;
    wire signal_23010 ;
    wire signal_23011 ;
    wire signal_23012 ;
    wire signal_23013 ;
    wire signal_23014 ;
    wire signal_23015 ;
    wire signal_23016 ;
    wire signal_23017 ;
    wire signal_23018 ;
    wire signal_23019 ;
    wire signal_23020 ;
    wire signal_23021 ;
    wire signal_23022 ;
    wire signal_23023 ;
    wire signal_23024 ;
    wire signal_23025 ;
    wire signal_23026 ;
    wire signal_23027 ;
    wire signal_23028 ;
    wire signal_23029 ;
    wire signal_23030 ;
    wire signal_23031 ;
    wire signal_23032 ;
    wire signal_23033 ;
    wire signal_23034 ;
    wire signal_23035 ;
    wire signal_23036 ;
    wire signal_23037 ;
    wire signal_23038 ;
    wire signal_23039 ;
    wire signal_23040 ;
    wire signal_23041 ;
    wire signal_23042 ;
    wire signal_23043 ;
    wire signal_23044 ;
    wire signal_23045 ;
    wire signal_23046 ;
    wire signal_23047 ;
    wire signal_23048 ;
    wire signal_23049 ;
    wire signal_23050 ;
    wire signal_23051 ;
    wire signal_23052 ;
    wire signal_23053 ;
    wire signal_23054 ;
    wire signal_23055 ;
    wire signal_23056 ;
    wire signal_23057 ;
    wire signal_23058 ;
    wire signal_23059 ;
    wire signal_23060 ;
    wire signal_23061 ;
    wire signal_23062 ;
    wire signal_23063 ;
    wire signal_23064 ;
    wire signal_23065 ;
    wire signal_23066 ;
    wire signal_23067 ;
    wire signal_23068 ;
    wire signal_23069 ;
    wire signal_23070 ;
    wire signal_23071 ;
    wire signal_23072 ;
    wire signal_23073 ;
    wire signal_23074 ;
    wire signal_23075 ;
    wire signal_23076 ;
    wire signal_23077 ;
    wire signal_23078 ;
    wire signal_23079 ;
    wire signal_23080 ;
    wire signal_23081 ;
    wire signal_23082 ;
    wire signal_23083 ;
    wire signal_23084 ;
    wire signal_23085 ;
    wire signal_23086 ;
    wire signal_23087 ;
    wire signal_23088 ;
    wire signal_23089 ;
    wire signal_23090 ;
    wire signal_23091 ;
    wire signal_23092 ;
    wire signal_23093 ;
    wire signal_23094 ;
    wire signal_23095 ;
    wire signal_23096 ;
    wire signal_23097 ;
    wire signal_23098 ;
    wire signal_23099 ;
    wire signal_23100 ;
    wire signal_23101 ;
    wire signal_23102 ;
    wire signal_23103 ;
    wire signal_23104 ;
    wire signal_23105 ;
    wire signal_23106 ;
    wire signal_23107 ;
    wire signal_23108 ;
    wire signal_23109 ;
    wire signal_23110 ;
    wire signal_23111 ;
    wire signal_23112 ;
    wire signal_23113 ;
    wire signal_23114 ;
    wire signal_23115 ;
    wire signal_23116 ;
    wire signal_23117 ;
    wire signal_23118 ;
    wire signal_23119 ;
    wire signal_23120 ;
    wire signal_23121 ;
    wire signal_23122 ;
    wire signal_23123 ;
    wire signal_23124 ;
    wire signal_23125 ;
    wire signal_23126 ;
    wire signal_23127 ;
    wire signal_23128 ;
    wire signal_23129 ;
    wire signal_23130 ;
    wire signal_23131 ;
    wire signal_23132 ;
    wire signal_23133 ;
    wire signal_23134 ;
    wire signal_23135 ;
    wire signal_23136 ;
    wire signal_23137 ;
    wire signal_23138 ;
    wire signal_23139 ;
    wire signal_23140 ;
    wire signal_23141 ;
    wire signal_23142 ;
    wire signal_23143 ;
    wire signal_23144 ;
    wire signal_23145 ;
    wire signal_23146 ;
    wire signal_23147 ;
    wire signal_23148 ;
    wire signal_23149 ;
    wire signal_23150 ;
    wire signal_23151 ;
    wire signal_23152 ;
    wire signal_23153 ;
    wire signal_23154 ;
    wire signal_23155 ;
    wire signal_23156 ;
    wire signal_23157 ;
    wire signal_23158 ;
    wire signal_23159 ;
    wire signal_23160 ;
    wire signal_23161 ;
    wire signal_23162 ;
    wire signal_23163 ;
    wire signal_23164 ;
    wire signal_23165 ;
    wire signal_23166 ;
    wire signal_23167 ;
    wire signal_23168 ;
    wire signal_23169 ;
    wire signal_23170 ;
    wire signal_23171 ;
    wire signal_23172 ;
    wire signal_23173 ;
    wire signal_23174 ;
    wire signal_23175 ;
    wire signal_23176 ;
    wire signal_23177 ;
    wire signal_23178 ;
    wire signal_23179 ;
    wire signal_23180 ;
    wire signal_23181 ;
    wire signal_23182 ;
    wire signal_23183 ;
    wire signal_23184 ;
    wire signal_23185 ;
    wire signal_23186 ;
    wire signal_23187 ;
    wire signal_23188 ;
    wire signal_23189 ;
    wire signal_23190 ;
    wire signal_23191 ;
    wire signal_23192 ;
    wire signal_23193 ;
    wire signal_23194 ;
    wire signal_23195 ;
    wire signal_23196 ;
    wire signal_23197 ;
    wire signal_23198 ;
    wire signal_23199 ;
    wire signal_23200 ;
    wire signal_23201 ;
    wire signal_23202 ;
    wire signal_23203 ;
    wire signal_23204 ;
    wire signal_23205 ;
    wire signal_23206 ;
    wire signal_23207 ;
    wire signal_23208 ;
    wire signal_23209 ;
    wire signal_23210 ;
    wire signal_23211 ;
    wire signal_23212 ;
    wire signal_23213 ;
    wire signal_23214 ;
    wire signal_23215 ;
    wire signal_23216 ;
    wire signal_23217 ;
    wire signal_23218 ;
    wire signal_23219 ;
    wire signal_23220 ;
    wire signal_23221 ;
    wire signal_23222 ;
    wire signal_23223 ;
    wire signal_23224 ;
    wire signal_23225 ;
    wire signal_23226 ;
    wire signal_23227 ;
    wire signal_23228 ;
    wire signal_23229 ;
    wire signal_23230 ;
    wire signal_23231 ;
    wire signal_23232 ;
    wire signal_23233 ;
    wire signal_23234 ;
    wire signal_23235 ;
    wire signal_23236 ;
    wire signal_23237 ;
    wire signal_23238 ;
    wire signal_23239 ;
    wire signal_23240 ;
    wire signal_23241 ;
    wire signal_23242 ;
    wire signal_23243 ;
    wire signal_23244 ;
    wire signal_23245 ;
    wire signal_23246 ;
    wire signal_23247 ;
    wire signal_23248 ;
    wire signal_23249 ;
    wire signal_23250 ;
    wire signal_23251 ;
    wire signal_23252 ;
    wire signal_23253 ;
    wire signal_23254 ;
    wire signal_23255 ;
    wire signal_23256 ;
    wire signal_23257 ;
    wire signal_23258 ;
    wire signal_23259 ;
    wire signal_23260 ;
    wire signal_23261 ;
    wire signal_23262 ;
    wire signal_23263 ;
    wire signal_23264 ;
    wire signal_23265 ;
    wire signal_23266 ;
    wire signal_23267 ;
    wire signal_23268 ;
    wire signal_23269 ;
    wire signal_23270 ;
    wire signal_23271 ;
    wire signal_23272 ;
    wire signal_23273 ;
    wire signal_23274 ;
    wire signal_23275 ;
    wire signal_23276 ;
    wire signal_23277 ;
    wire signal_23278 ;
    wire signal_23279 ;
    wire signal_23280 ;
    wire signal_23281 ;
    wire signal_23282 ;
    wire signal_23283 ;
    wire signal_23284 ;
    wire signal_23285 ;
    wire signal_23286 ;
    wire signal_23287 ;
    wire signal_23288 ;
    wire signal_23289 ;
    wire signal_23290 ;
    wire signal_23291 ;
    wire signal_23292 ;
    wire signal_23293 ;
    wire signal_23294 ;
    wire signal_23295 ;
    wire signal_23296 ;
    wire signal_23297 ;
    wire signal_23298 ;
    wire signal_23299 ;
    wire signal_23300 ;
    wire signal_23301 ;
    wire signal_23302 ;
    wire signal_23303 ;
    wire signal_23304 ;
    wire signal_23305 ;
    wire signal_23306 ;
    wire signal_23307 ;
    wire signal_23308 ;
    wire signal_23309 ;
    wire signal_23310 ;
    wire signal_23311 ;
    wire signal_23312 ;
    wire signal_23313 ;
    wire signal_23314 ;
    wire signal_23315 ;
    wire signal_23316 ;
    wire signal_23317 ;
    wire signal_23318 ;
    wire signal_23319 ;
    wire signal_23320 ;
    wire signal_23321 ;
    wire signal_23322 ;
    wire signal_23323 ;
    wire signal_23324 ;
    wire signal_23325 ;
    wire signal_23326 ;
    wire signal_23327 ;
    wire signal_23328 ;
    wire signal_23329 ;
    wire signal_23330 ;
    wire signal_23331 ;
    wire signal_23332 ;
    wire signal_23333 ;
    wire signal_23334 ;
    wire signal_23335 ;
    wire signal_23336 ;
    wire signal_23337 ;
    wire signal_23338 ;
    wire signal_23339 ;
    wire signal_23340 ;
    wire signal_23341 ;
    wire signal_23342 ;
    wire signal_23343 ;
    wire signal_23344 ;
    wire signal_23345 ;
    wire signal_23346 ;
    wire signal_23347 ;
    wire signal_23348 ;
    wire signal_23349 ;
    wire signal_23350 ;
    wire signal_23351 ;
    wire signal_23352 ;
    wire signal_23353 ;
    wire signal_23354 ;
    wire signal_23355 ;
    wire signal_23356 ;
    wire signal_23357 ;
    wire signal_23358 ;
    wire signal_23359 ;
    wire signal_23360 ;
    wire signal_23361 ;
    wire signal_23362 ;
    wire signal_23363 ;
    wire signal_23364 ;
    wire signal_23365 ;
    wire signal_23366 ;
    wire signal_23367 ;
    wire signal_23368 ;
    wire signal_23369 ;
    wire signal_23370 ;
    wire signal_23371 ;
    wire signal_23372 ;
    wire signal_23373 ;
    wire signal_23374 ;
    wire signal_23375 ;
    wire signal_23376 ;
    wire signal_23377 ;
    wire signal_23378 ;
    wire signal_23379 ;
    wire signal_23380 ;
    wire signal_23381 ;
    wire signal_23382 ;
    wire signal_23383 ;
    wire signal_23384 ;
    wire signal_23385 ;
    wire signal_23386 ;
    wire signal_23387 ;
    wire signal_23388 ;
    wire signal_23389 ;
    wire signal_23390 ;
    wire signal_23391 ;
    wire signal_23392 ;
    wire signal_23393 ;
    wire signal_23394 ;
    wire signal_23395 ;
    wire signal_23396 ;
    wire signal_23397 ;
    wire signal_23398 ;
    wire signal_23399 ;
    wire signal_23400 ;
    wire signal_23401 ;
    wire signal_23402 ;
    wire signal_23403 ;
    wire signal_23404 ;
    wire signal_23405 ;
    wire signal_23406 ;
    wire signal_23407 ;
    wire signal_23408 ;
    wire signal_23409 ;
    wire signal_23410 ;
    wire signal_23411 ;
    wire signal_23412 ;
    wire signal_23413 ;
    wire signal_23414 ;
    wire signal_23415 ;
    wire signal_23416 ;
    wire signal_23417 ;
    wire signal_23418 ;
    wire signal_23419 ;
    wire signal_23420 ;
    wire signal_23421 ;
    wire signal_23422 ;
    wire signal_23423 ;
    wire signal_23424 ;
    wire signal_23425 ;
    wire signal_23426 ;
    wire signal_23427 ;
    wire signal_23428 ;
    wire signal_23429 ;
    wire signal_23430 ;
    wire signal_23431 ;
    wire signal_23432 ;
    wire signal_23433 ;
    wire signal_23434 ;
    wire signal_23435 ;
    wire signal_23436 ;
    wire signal_23437 ;
    wire signal_23438 ;
    wire signal_23439 ;
    wire signal_23440 ;
    wire signal_23441 ;
    wire signal_23442 ;
    wire signal_23443 ;
    wire signal_23444 ;
    wire signal_23445 ;
    wire signal_23446 ;
    wire signal_23447 ;
    wire signal_23448 ;
    wire signal_23449 ;
    wire signal_23450 ;
    wire signal_23451 ;
    wire signal_23452 ;
    wire signal_23453 ;
    wire signal_23454 ;
    wire signal_23455 ;
    wire signal_23456 ;
    wire signal_23457 ;
    wire signal_23458 ;
    wire signal_23459 ;
    wire signal_23460 ;
    wire signal_23461 ;
    wire signal_23462 ;
    wire signal_23463 ;
    wire signal_23464 ;
    wire signal_23465 ;
    wire signal_23466 ;
    wire signal_23467 ;
    wire signal_23468 ;
    wire signal_23469 ;
    wire signal_23470 ;
    wire signal_23471 ;
    wire signal_23472 ;
    wire signal_23473 ;
    wire signal_23474 ;
    wire signal_23475 ;
    wire signal_23476 ;
    wire signal_23477 ;
    wire signal_23478 ;
    wire signal_23479 ;
    wire signal_23480 ;
    wire signal_23481 ;
    wire signal_23482 ;
    wire signal_23483 ;
    wire signal_23484 ;
    wire signal_23485 ;
    wire signal_23486 ;
    wire signal_23487 ;
    wire signal_23488 ;
    wire signal_23489 ;
    wire signal_23490 ;
    wire signal_23491 ;
    wire signal_23492 ;
    wire signal_23493 ;
    wire signal_23494 ;
    wire signal_23495 ;
    wire signal_23496 ;
    wire signal_23497 ;
    wire signal_23498 ;
    wire signal_23499 ;
    wire signal_23500 ;
    wire signal_23501 ;
    wire signal_23502 ;
    wire signal_23503 ;
    wire signal_23504 ;
    wire signal_23505 ;
    wire signal_23506 ;
    wire signal_23507 ;
    wire signal_23508 ;
    wire signal_23509 ;
    wire signal_23510 ;
    wire signal_23511 ;
    wire signal_23512 ;
    wire signal_23513 ;
    wire signal_23514 ;
    wire signal_23515 ;
    wire signal_23516 ;
    wire signal_23517 ;
    wire signal_23518 ;
    wire signal_23519 ;
    wire signal_23520 ;
    wire signal_23521 ;
    wire signal_23522 ;
    wire signal_23523 ;
    wire signal_23524 ;
    wire signal_23525 ;
    wire signal_23526 ;
    wire signal_23527 ;
    wire signal_23528 ;
    wire signal_23529 ;
    wire signal_23530 ;
    wire signal_23531 ;
    wire signal_23532 ;
    wire signal_23533 ;
    wire signal_23534 ;
    wire signal_23535 ;
    wire signal_23536 ;
    wire signal_23537 ;
    wire signal_23538 ;
    wire signal_23539 ;
    wire signal_23540 ;
    wire signal_23541 ;
    wire signal_23542 ;
    wire signal_23543 ;
    wire signal_23544 ;
    wire signal_23545 ;
    wire signal_23546 ;
    wire signal_23547 ;
    wire signal_23548 ;
    wire signal_23549 ;
    wire signal_23550 ;
    wire signal_23551 ;
    wire signal_23552 ;
    wire signal_23553 ;
    wire signal_23554 ;
    wire signal_23555 ;
    wire signal_23556 ;
    wire signal_23557 ;
    wire signal_23558 ;
    wire signal_23559 ;
    wire signal_23560 ;
    wire signal_23561 ;
    wire signal_23562 ;
    wire signal_23563 ;
    wire signal_23564 ;
    wire signal_23565 ;
    wire signal_23566 ;
    wire signal_23567 ;
    wire signal_23568 ;
    wire signal_23569 ;
    wire signal_23570 ;
    wire signal_23571 ;
    wire signal_23572 ;
    wire signal_23573 ;
    wire signal_23574 ;
    wire signal_23575 ;
    wire signal_23576 ;
    wire signal_23577 ;
    wire signal_23578 ;
    wire signal_23579 ;
    wire signal_23580 ;
    wire signal_23581 ;
    wire signal_23582 ;
    wire signal_23583 ;
    wire signal_23584 ;
    wire signal_23585 ;
    wire signal_23586 ;
    wire signal_23587 ;
    wire signal_23588 ;
    wire signal_23589 ;
    wire signal_23590 ;
    wire signal_23591 ;
    wire signal_23592 ;
    wire signal_23593 ;
    wire signal_23594 ;
    wire signal_23595 ;
    wire signal_23596 ;
    wire signal_23597 ;
    wire signal_23598 ;
    wire signal_23599 ;
    wire signal_23600 ;
    wire signal_23601 ;
    wire signal_23602 ;
    wire signal_23603 ;
    wire signal_23604 ;
    wire signal_23605 ;
    wire signal_23606 ;
    wire signal_23607 ;
    wire signal_23608 ;
    wire signal_23609 ;
    wire signal_23610 ;
    wire signal_23611 ;
    wire signal_23612 ;
    wire signal_23613 ;
    wire signal_23614 ;
    wire signal_23615 ;
    wire signal_23616 ;
    wire signal_23617 ;
    wire signal_23618 ;
    wire signal_23619 ;
    wire signal_23620 ;
    wire signal_23621 ;
    wire signal_23622 ;
    wire signal_23623 ;
    wire signal_23624 ;
    wire signal_23625 ;
    wire signal_23626 ;
    wire signal_23627 ;
    wire signal_23628 ;
    wire signal_23629 ;
    wire signal_23630 ;
    wire signal_23631 ;
    wire signal_23632 ;
    wire signal_23633 ;
    wire signal_23634 ;
    wire signal_23635 ;
    wire signal_23636 ;
    wire signal_23637 ;
    wire signal_23638 ;
    wire signal_23639 ;
    wire signal_23640 ;
    wire signal_23641 ;
    wire signal_23642 ;
    wire signal_23643 ;
    wire signal_23644 ;
    wire signal_23645 ;
    wire signal_23646 ;
    wire signal_23647 ;
    wire signal_23648 ;
    wire signal_23649 ;
    wire signal_23650 ;
    wire signal_23651 ;
    wire signal_23652 ;
    wire signal_23653 ;
    wire signal_23654 ;
    wire signal_23655 ;
    wire signal_23656 ;
    wire signal_23657 ;
    wire signal_23658 ;
    wire signal_23659 ;
    wire signal_23660 ;
    wire signal_23661 ;
    wire signal_23662 ;
    wire signal_23663 ;
    wire signal_23664 ;
    wire signal_23665 ;
    wire signal_23666 ;
    wire signal_23667 ;
    wire signal_23668 ;
    wire signal_23669 ;
    wire signal_23670 ;
    wire signal_23671 ;
    wire signal_23672 ;
    wire signal_23673 ;
    wire signal_23674 ;
    wire signal_23675 ;
    wire signal_23676 ;
    wire signal_23677 ;
    wire signal_23678 ;
    wire signal_23679 ;
    wire signal_23680 ;
    wire signal_23681 ;
    wire signal_23682 ;
    wire signal_23683 ;
    wire signal_23684 ;
    wire signal_23685 ;
    wire signal_23686 ;
    wire signal_23687 ;
    wire signal_23688 ;
    wire signal_23689 ;
    wire signal_23690 ;
    wire signal_23691 ;
    wire signal_23692 ;
    wire signal_23693 ;
    wire signal_23694 ;
    wire signal_23695 ;
    wire signal_23696 ;
    wire signal_23697 ;
    wire signal_23698 ;
    wire signal_23699 ;
    wire signal_23700 ;
    wire signal_23701 ;
    wire signal_23702 ;
    wire signal_23703 ;
    wire signal_23704 ;
    wire signal_23705 ;
    wire signal_23706 ;
    wire signal_23707 ;
    wire signal_23708 ;
    wire signal_23709 ;
    wire signal_23710 ;
    wire signal_23711 ;
    wire signal_23712 ;
    wire signal_23713 ;
    wire signal_23714 ;
    wire signal_23715 ;
    wire signal_23716 ;
    wire signal_23717 ;
    wire signal_23718 ;
    wire signal_23719 ;
    wire signal_23720 ;
    wire signal_23721 ;
    wire signal_23722 ;
    wire signal_23723 ;
    wire signal_23724 ;
    wire signal_23725 ;
    wire signal_23726 ;
    wire signal_23727 ;
    wire signal_23728 ;
    wire signal_23729 ;
    wire signal_23730 ;
    wire signal_23731 ;
    wire signal_23732 ;
    wire signal_23733 ;
    wire signal_23734 ;
    wire signal_23735 ;
    wire signal_23736 ;
    wire signal_23737 ;
    wire signal_23738 ;
    wire signal_23739 ;
    wire signal_23740 ;
    wire signal_23741 ;
    wire signal_23742 ;
    wire signal_23743 ;
    wire signal_23744 ;
    wire signal_23745 ;
    wire signal_23746 ;
    wire signal_23747 ;
    wire signal_23748 ;
    wire signal_23749 ;
    wire signal_23750 ;
    wire signal_23751 ;
    wire signal_23752 ;
    wire signal_23753 ;
    wire signal_23754 ;
    wire signal_23755 ;
    wire signal_23756 ;
    wire signal_23757 ;
    wire signal_23758 ;
    wire signal_23759 ;
    wire signal_23760 ;
    wire signal_23761 ;
    wire signal_23762 ;
    wire signal_23763 ;
    wire signal_23764 ;
    wire signal_23765 ;
    wire signal_23766 ;
    wire signal_23767 ;
    wire signal_23768 ;
    wire signal_23769 ;
    wire signal_23770 ;
    wire signal_23771 ;
    wire signal_23772 ;
    wire signal_23773 ;
    wire signal_23774 ;
    wire signal_23775 ;
    wire signal_23776 ;
    wire signal_23777 ;
    wire signal_23778 ;
    wire signal_23779 ;
    wire signal_23780 ;
    wire signal_23781 ;
    wire signal_23782 ;
    wire signal_23783 ;
    wire signal_23784 ;
    wire signal_23785 ;
    wire signal_23786 ;
    wire signal_23787 ;
    wire signal_23788 ;
    wire signal_23789 ;
    wire signal_23790 ;
    wire signal_23791 ;
    wire signal_23792 ;
    wire signal_23793 ;
    wire signal_23794 ;
    wire signal_23795 ;
    wire signal_23796 ;
    wire signal_23797 ;
    wire signal_23798 ;
    wire signal_23799 ;
    wire signal_23800 ;
    wire signal_23801 ;
    wire signal_23802 ;
    wire signal_23803 ;
    wire signal_23804 ;
    wire signal_23805 ;
    wire signal_23806 ;
    wire signal_23807 ;
    wire signal_23808 ;
    wire signal_23809 ;
    wire signal_23810 ;
    wire signal_23811 ;
    wire signal_23812 ;
    wire signal_23813 ;
    wire signal_23814 ;
    wire signal_23815 ;
    wire signal_23816 ;
    wire signal_23817 ;
    wire signal_23818 ;
    wire signal_23819 ;
    wire signal_23820 ;
    wire signal_23821 ;
    wire signal_23822 ;
    wire signal_23823 ;
    wire signal_23824 ;
    wire signal_23825 ;
    wire signal_23826 ;
    wire signal_23827 ;
    wire signal_23828 ;
    wire signal_23829 ;
    wire signal_23830 ;
    wire signal_23831 ;
    wire signal_23832 ;
    wire signal_23833 ;
    wire signal_23834 ;
    wire signal_23835 ;
    wire signal_23836 ;
    wire signal_23837 ;
    wire signal_23838 ;
    wire signal_23839 ;
    wire signal_23840 ;
    wire signal_23841 ;
    wire signal_23842 ;
    wire signal_23843 ;
    wire signal_23844 ;
    wire signal_23845 ;
    wire signal_23846 ;
    wire signal_23847 ;
    wire signal_23848 ;
    wire signal_23849 ;
    wire signal_23850 ;
    wire signal_23851 ;
    wire signal_23852 ;
    wire signal_23853 ;
    wire signal_23854 ;
    wire signal_23855 ;
    wire signal_23856 ;
    wire signal_23857 ;
    wire signal_23858 ;
    wire signal_23859 ;
    wire signal_23860 ;
    wire signal_23861 ;
    wire signal_23862 ;
    wire signal_23863 ;
    wire signal_23864 ;
    wire signal_23865 ;
    wire signal_23866 ;
    wire signal_23867 ;
    wire signal_23868 ;
    wire signal_23869 ;
    wire signal_23870 ;
    wire signal_23871 ;
    wire signal_23872 ;
    wire signal_23873 ;
    wire signal_23874 ;
    wire signal_23875 ;
    wire signal_23876 ;
    wire signal_23877 ;
    wire signal_23878 ;
    wire signal_23879 ;
    wire signal_23880 ;
    wire signal_23881 ;
    wire signal_23882 ;
    wire signal_23883 ;
    wire signal_23884 ;
    wire signal_23885 ;
    wire signal_23886 ;
    wire signal_23887 ;
    wire signal_23888 ;
    wire signal_23889 ;
    wire signal_23890 ;
    wire signal_23891 ;
    wire signal_23892 ;
    wire signal_23893 ;
    wire signal_23894 ;
    wire signal_23895 ;
    wire signal_23896 ;
    wire signal_23897 ;
    wire signal_23898 ;
    wire signal_23899 ;
    wire signal_23900 ;
    wire signal_23901 ;
    wire signal_23902 ;
    wire signal_23903 ;
    wire signal_23904 ;
    wire signal_23905 ;
    wire signal_23906 ;
    wire signal_23907 ;
    wire signal_23908 ;
    wire signal_23909 ;
    wire signal_23910 ;
    wire signal_23911 ;
    wire signal_23912 ;
    wire signal_23913 ;
    wire signal_23914 ;
    wire signal_23915 ;
    wire signal_23916 ;
    wire signal_23917 ;
    wire signal_23918 ;
    wire signal_23919 ;
    wire signal_23920 ;
    wire signal_23921 ;
    wire signal_23922 ;
    wire signal_23923 ;
    wire signal_23924 ;
    wire signal_23925 ;
    wire signal_23926 ;
    wire signal_23927 ;
    wire signal_23928 ;
    wire signal_23929 ;
    wire signal_23930 ;
    wire signal_23931 ;
    wire signal_23932 ;
    wire signal_23933 ;
    wire signal_23934 ;
    wire signal_23935 ;
    wire signal_23936 ;
    wire signal_23937 ;
    wire signal_23938 ;
    wire signal_23939 ;
    wire signal_23940 ;
    wire signal_23941 ;
    wire signal_23942 ;
    wire signal_23943 ;
    wire signal_23944 ;
    wire signal_23945 ;
    wire signal_23946 ;
    wire signal_23947 ;
    wire signal_23948 ;
    wire signal_23949 ;
    wire signal_23950 ;
    wire signal_23951 ;
    wire signal_23952 ;
    wire signal_23953 ;
    wire signal_23954 ;
    wire signal_23955 ;
    wire signal_23956 ;
    wire signal_23957 ;
    wire signal_23958 ;
    wire signal_23959 ;
    wire signal_23960 ;
    wire signal_23961 ;
    wire signal_23962 ;
    wire signal_23963 ;
    wire signal_23964 ;
    wire signal_23965 ;
    wire signal_23966 ;
    wire signal_23967 ;
    wire signal_23968 ;
    wire signal_23969 ;
    wire signal_23970 ;
    wire signal_23971 ;
    wire signal_23972 ;
    wire signal_23973 ;
    wire signal_23974 ;
    wire signal_23975 ;
    wire signal_23976 ;
    wire signal_23977 ;
    wire signal_23978 ;
    wire signal_23979 ;
    wire signal_23980 ;
    wire signal_23981 ;
    wire signal_23982 ;
    wire signal_23983 ;
    wire signal_23984 ;
    wire signal_23985 ;
    wire signal_23986 ;
    wire signal_23987 ;
    wire signal_23988 ;
    wire signal_23989 ;
    wire signal_23990 ;
    wire signal_23991 ;
    wire signal_23992 ;
    wire signal_23993 ;
    wire signal_23994 ;
    wire signal_23995 ;
    wire signal_23996 ;
    wire signal_23997 ;
    wire signal_23998 ;
    wire signal_23999 ;
    wire signal_24000 ;
    wire signal_24001 ;
    wire signal_24002 ;
    wire signal_24003 ;
    wire signal_24004 ;
    wire signal_24005 ;
    wire signal_24006 ;
    wire signal_24007 ;
    wire signal_24008 ;
    wire signal_24009 ;
    wire signal_24010 ;
    wire signal_24011 ;
    wire signal_24012 ;
    wire signal_24013 ;
    wire signal_24014 ;
    wire signal_24015 ;
    wire signal_24016 ;
    wire signal_24017 ;
    wire signal_24018 ;
    wire signal_24019 ;
    wire signal_24020 ;
    wire signal_24021 ;
    wire signal_24022 ;
    wire signal_24023 ;
    wire signal_24024 ;
    wire signal_24025 ;
    wire signal_24026 ;
    wire signal_24027 ;
    wire signal_24028 ;
    wire signal_24029 ;
    wire signal_24030 ;
    wire signal_24031 ;
    wire signal_24032 ;
    wire signal_24033 ;
    wire signal_24034 ;
    wire signal_24035 ;
    wire signal_24036 ;
    wire signal_24037 ;
    wire signal_24038 ;
    wire signal_24039 ;
    wire signal_24040 ;
    wire signal_24041 ;
    wire signal_24042 ;
    wire signal_24043 ;
    wire signal_24044 ;
    wire signal_24045 ;
    wire signal_24046 ;
    wire signal_24047 ;
    wire signal_24048 ;
    wire signal_24049 ;
    wire signal_24050 ;
    wire signal_24051 ;
    wire signal_24052 ;
    wire signal_24053 ;
    wire signal_24054 ;
    wire signal_24055 ;
    wire signal_24056 ;
    wire signal_24057 ;
    wire signal_24058 ;
    wire signal_24059 ;
    wire signal_24060 ;
    wire signal_24061 ;
    wire signal_24062 ;
    wire signal_24063 ;
    wire signal_24064 ;
    wire signal_24065 ;
    wire signal_24066 ;
    wire signal_24067 ;
    wire signal_24068 ;
    wire signal_24069 ;
    wire signal_24070 ;
    wire signal_24071 ;
    wire signal_24072 ;
    wire signal_24073 ;
    wire signal_24074 ;
    wire signal_24075 ;
    wire signal_24076 ;
    wire signal_24077 ;
    wire signal_24078 ;
    wire signal_24079 ;
    wire signal_24080 ;
    wire signal_24081 ;
    wire signal_24082 ;
    wire signal_24083 ;
    wire signal_24084 ;
    wire signal_24085 ;
    wire signal_24086 ;
    wire signal_24087 ;
    wire signal_24088 ;
    wire signal_24089 ;
    wire signal_24090 ;
    wire signal_24091 ;
    wire signal_24092 ;
    wire signal_24093 ;
    wire signal_24094 ;
    wire signal_24095 ;
    wire signal_24096 ;
    wire signal_24097 ;
    wire signal_24098 ;
    wire signal_24099 ;
    wire signal_24100 ;
    wire signal_24101 ;
    wire signal_24102 ;
    wire signal_24103 ;
    wire signal_24104 ;
    wire signal_24105 ;
    wire signal_24106 ;
    wire signal_24107 ;
    wire signal_24108 ;
    wire signal_24109 ;
    wire signal_24110 ;
    wire signal_24111 ;
    wire signal_24112 ;
    wire signal_24113 ;
    wire signal_24114 ;
    wire signal_24115 ;
    wire signal_24116 ;
    wire signal_24117 ;
    wire signal_24118 ;
    wire signal_24119 ;
    wire signal_24120 ;
    wire signal_24121 ;
    wire signal_24122 ;
    wire signal_24123 ;
    wire signal_24124 ;
    wire signal_24125 ;
    wire signal_24126 ;
    wire signal_24127 ;
    wire signal_24128 ;
    wire signal_24129 ;
    wire signal_24130 ;
    wire signal_24131 ;
    wire signal_24132 ;
    wire signal_24133 ;
    wire signal_24134 ;
    wire signal_24135 ;
    wire signal_24136 ;
    wire signal_24137 ;
    wire signal_24138 ;
    wire signal_24139 ;
    wire signal_24140 ;
    wire signal_24141 ;
    wire signal_24142 ;
    wire signal_24143 ;
    wire signal_24144 ;
    wire signal_24145 ;
    wire signal_24146 ;
    wire signal_24147 ;
    wire signal_24148 ;
    wire signal_24149 ;
    wire signal_24150 ;
    wire signal_24151 ;
    wire signal_24152 ;
    wire signal_24153 ;
    wire signal_24154 ;
    wire signal_24155 ;
    wire signal_24156 ;
    wire signal_24157 ;
    wire signal_24158 ;
    wire signal_24159 ;
    wire signal_24160 ;
    wire signal_24161 ;
    wire signal_24162 ;
    wire signal_24163 ;
    wire signal_24164 ;
    wire signal_24165 ;
    wire signal_24166 ;
    wire signal_24167 ;
    wire signal_24168 ;
    wire signal_24169 ;
    wire signal_24170 ;
    wire signal_24171 ;
    wire signal_24172 ;
    wire signal_24173 ;
    wire signal_24174 ;
    wire signal_24175 ;
    wire signal_24176 ;
    wire signal_24177 ;
    wire signal_24178 ;
    wire signal_24179 ;
    wire signal_24180 ;
    wire signal_24181 ;
    wire signal_24182 ;
    wire signal_24183 ;
    wire signal_24184 ;
    wire signal_24185 ;
    wire signal_24186 ;
    wire signal_24187 ;
    wire signal_24188 ;
    wire signal_24189 ;
    wire signal_24190 ;
    wire signal_24191 ;
    wire signal_24192 ;
    wire signal_24193 ;
    wire signal_24194 ;
    wire signal_24195 ;
    wire signal_24196 ;
    wire signal_24197 ;
    wire signal_24198 ;
    wire signal_24199 ;
    wire signal_24200 ;
    wire signal_24201 ;
    wire signal_24202 ;
    wire signal_24203 ;
    wire signal_24204 ;
    wire signal_24205 ;
    wire signal_24206 ;
    wire signal_24207 ;
    wire signal_24208 ;
    wire signal_24209 ;
    wire signal_24210 ;
    wire signal_24211 ;
    wire signal_24212 ;
    wire signal_24213 ;
    wire signal_24214 ;
    wire signal_24215 ;
    wire signal_24216 ;
    wire signal_24217 ;
    wire signal_24218 ;
    wire signal_24219 ;
    wire signal_24220 ;
    wire signal_24221 ;
    wire signal_24222 ;
    wire signal_24223 ;
    wire signal_24224 ;
    wire signal_24225 ;
    wire signal_24226 ;
    wire signal_24227 ;
    wire signal_24228 ;
    wire signal_24229 ;
    wire signal_24230 ;
    wire signal_24231 ;
    wire signal_24232 ;
    wire signal_24233 ;
    wire signal_24234 ;
    wire signal_24235 ;
    wire signal_24236 ;
    wire signal_24237 ;
    wire signal_24238 ;
    wire signal_24239 ;
    wire signal_24240 ;
    wire signal_24241 ;
    wire signal_24242 ;
    wire signal_24243 ;
    wire signal_24244 ;
    wire signal_24245 ;
    wire signal_24246 ;
    wire signal_24247 ;
    wire signal_24248 ;
    wire signal_24249 ;
    wire signal_24250 ;
    wire signal_24251 ;
    wire signal_24252 ;
    wire signal_24253 ;
    wire signal_24254 ;
    wire signal_24255 ;
    wire signal_24256 ;
    wire signal_24257 ;
    wire signal_24258 ;
    wire signal_24259 ;
    wire signal_24260 ;
    wire signal_24261 ;
    wire signal_24262 ;
    wire signal_24263 ;
    wire signal_24264 ;
    wire signal_24265 ;
    wire signal_24266 ;
    wire signal_24267 ;
    wire signal_24268 ;
    wire signal_24269 ;
    wire signal_24270 ;
    wire signal_24271 ;
    wire signal_24272 ;
    wire signal_24273 ;
    wire signal_24274 ;
    wire signal_24275 ;
    wire signal_24276 ;
    wire signal_24277 ;
    wire signal_24278 ;
    wire signal_24279 ;
    wire signal_24280 ;
    wire signal_24281 ;
    wire signal_24282 ;
    wire signal_24283 ;
    wire signal_24284 ;
    wire signal_24285 ;
    wire signal_24286 ;
    wire signal_24287 ;
    wire signal_24288 ;
    wire signal_24289 ;
    wire signal_24290 ;
    wire signal_24291 ;
    wire signal_24292 ;
    wire signal_24293 ;
    wire signal_24294 ;
    wire signal_24295 ;
    wire signal_24296 ;
    wire signal_24297 ;
    wire signal_24298 ;
    wire signal_24299 ;
    wire signal_24300 ;
    wire signal_24301 ;
    wire signal_24302 ;
    wire signal_24303 ;
    wire signal_24304 ;
    wire signal_24305 ;
    wire signal_24306 ;
    wire signal_24307 ;
    wire signal_24308 ;
    wire signal_24309 ;
    wire signal_24310 ;
    wire signal_24311 ;
    wire signal_24312 ;
    wire signal_24313 ;
    wire signal_24314 ;
    wire signal_24315 ;
    wire signal_24316 ;
    wire signal_24317 ;
    wire signal_24318 ;
    wire signal_24319 ;
    wire signal_24320 ;
    wire signal_24321 ;
    wire signal_24322 ;
    wire signal_24323 ;
    wire signal_24324 ;
    wire signal_24325 ;
    wire signal_24326 ;
    wire signal_24327 ;
    wire signal_24328 ;
    wire signal_24329 ;
    wire signal_24330 ;
    wire signal_24331 ;
    wire signal_24332 ;
    wire signal_24333 ;
    wire signal_24334 ;
    wire signal_24335 ;
    wire signal_24336 ;
    wire signal_24337 ;
    wire signal_24338 ;
    wire signal_24339 ;
    wire signal_24340 ;
    wire signal_24341 ;
    wire signal_24342 ;
    wire signal_24343 ;
    wire signal_24344 ;
    wire signal_24345 ;
    wire signal_24346 ;
    wire signal_24347 ;
    wire signal_24348 ;
    wire signal_24349 ;
    wire signal_24350 ;
    wire signal_24351 ;
    wire signal_24352 ;
    wire signal_24353 ;
    wire signal_24354 ;
    wire signal_24355 ;
    wire signal_24356 ;
    wire signal_24357 ;
    wire signal_24358 ;
    wire signal_24359 ;
    wire signal_24360 ;
    wire signal_24361 ;
    wire signal_24362 ;
    wire signal_24363 ;
    wire signal_24364 ;
    wire signal_24365 ;
    wire signal_24366 ;
    wire signal_24367 ;
    wire signal_24368 ;
    wire signal_24369 ;
    wire signal_24370 ;
    wire signal_24371 ;
    wire signal_24372 ;
    wire signal_24373 ;
    wire signal_24374 ;
    wire signal_24375 ;
    wire signal_24376 ;
    wire signal_24377 ;
    wire signal_24378 ;
    wire signal_24379 ;
    wire signal_24380 ;
    wire signal_24381 ;
    wire signal_24382 ;
    wire signal_24383 ;
    wire signal_24384 ;
    wire signal_24385 ;
    wire signal_24386 ;
    wire signal_24387 ;
    wire signal_24388 ;
    wire signal_24389 ;
    wire signal_24390 ;
    wire signal_24391 ;
    wire signal_24392 ;
    wire signal_24393 ;
    wire signal_24394 ;
    wire signal_24395 ;
    wire signal_24396 ;
    wire signal_24397 ;
    wire signal_24398 ;
    wire signal_24399 ;
    wire signal_24400 ;
    wire signal_24401 ;
    wire signal_24402 ;
    wire signal_24403 ;
    wire signal_24404 ;
    wire signal_24405 ;
    wire signal_24406 ;
    wire signal_24407 ;
    wire signal_24408 ;
    wire signal_24409 ;
    wire signal_24410 ;
    wire signal_24411 ;
    wire signal_24412 ;
    wire signal_24413 ;
    wire signal_24414 ;
    wire signal_24415 ;
    wire signal_24416 ;
    wire signal_24417 ;
    wire signal_24418 ;
    wire signal_24419 ;
    wire signal_24420 ;
    wire signal_24421 ;
    wire signal_24422 ;
    wire signal_24423 ;
    wire signal_24424 ;
    wire signal_24425 ;
    wire signal_24426 ;
    wire signal_24427 ;
    wire signal_24428 ;
    wire signal_24429 ;
    wire signal_24430 ;
    wire signal_24431 ;
    wire signal_24432 ;
    wire signal_24433 ;
    wire signal_24434 ;
    wire signal_24435 ;
    wire signal_24436 ;
    wire signal_24437 ;
    wire signal_24438 ;
    wire signal_24439 ;
    wire signal_24440 ;
    wire signal_24441 ;
    wire signal_24442 ;
    wire signal_24443 ;
    wire signal_24444 ;
    wire signal_24445 ;
    wire signal_24446 ;
    wire signal_24447 ;
    wire signal_24448 ;
    wire signal_24449 ;
    wire signal_24450 ;
    wire signal_24451 ;
    wire signal_24452 ;
    wire signal_24453 ;
    wire signal_24454 ;
    wire signal_24455 ;
    wire signal_24456 ;
    wire signal_24457 ;
    wire signal_24458 ;
    wire signal_24459 ;
    wire signal_24460 ;
    wire signal_24461 ;
    wire signal_24462 ;
    wire signal_24463 ;
    wire signal_24464 ;
    wire signal_24465 ;
    wire signal_24466 ;
    wire signal_24467 ;
    wire signal_24468 ;
    wire signal_24469 ;
    wire signal_24470 ;
    wire signal_24471 ;
    wire signal_24472 ;
    wire signal_24473 ;
    wire signal_24474 ;
    wire signal_24475 ;
    wire signal_24476 ;
    wire signal_24477 ;
    wire signal_24478 ;
    wire signal_24479 ;
    wire signal_24480 ;
    wire signal_24481 ;
    wire signal_24482 ;
    wire signal_24483 ;
    wire signal_24484 ;
    wire signal_24485 ;
    wire signal_24486 ;
    wire signal_24487 ;
    wire signal_24488 ;
    wire signal_24489 ;
    wire signal_24490 ;
    wire signal_24491 ;
    wire signal_24492 ;
    wire signal_24493 ;
    wire signal_24494 ;
    wire signal_24495 ;
    wire signal_24496 ;
    wire signal_24497 ;
    wire signal_24498 ;
    wire signal_24499 ;
    wire signal_24500 ;
    wire signal_24501 ;
    wire signal_24502 ;
    wire signal_24503 ;
    wire signal_24504 ;
    wire signal_24505 ;
    wire signal_24506 ;
    wire signal_24507 ;
    wire signal_24508 ;
    wire signal_24509 ;
    wire signal_24510 ;
    wire signal_24511 ;
    wire signal_24512 ;
    wire signal_24513 ;
    wire signal_24514 ;
    wire signal_24515 ;
    wire signal_24516 ;
    wire signal_24517 ;
    wire signal_24518 ;
    wire signal_24519 ;
    wire signal_24520 ;
    wire signal_24521 ;
    wire signal_24522 ;
    wire signal_24523 ;
    wire signal_24524 ;
    wire signal_24525 ;
    wire signal_24526 ;
    wire signal_24527 ;
    wire signal_24528 ;
    wire signal_24529 ;
    wire signal_24530 ;
    wire signal_24531 ;
    wire signal_24532 ;
    wire signal_24533 ;
    wire signal_24534 ;
    wire signal_24535 ;
    wire signal_24536 ;
    wire signal_24537 ;
    wire signal_24538 ;
    wire signal_24539 ;
    wire signal_24540 ;
    wire signal_24541 ;
    wire signal_24542 ;
    wire signal_24543 ;
    wire signal_24544 ;
    wire signal_24545 ;
    wire signal_24546 ;
    wire signal_24547 ;
    wire signal_24548 ;
    wire signal_24549 ;
    wire signal_24550 ;
    wire signal_24551 ;
    wire signal_24552 ;
    wire signal_24553 ;
    wire signal_24554 ;
    wire signal_24555 ;
    wire signal_24556 ;
    wire signal_24557 ;
    wire signal_24558 ;
    wire signal_24559 ;
    wire signal_24560 ;
    wire signal_24561 ;
    wire signal_24562 ;
    wire signal_24563 ;
    wire signal_24564 ;
    wire signal_24565 ;
    wire signal_24566 ;
    wire signal_24567 ;
    wire signal_24568 ;
    wire signal_24569 ;
    wire signal_24570 ;
    wire signal_24571 ;
    wire signal_24572 ;
    wire signal_24573 ;
    wire signal_24574 ;
    wire signal_24575 ;
    wire signal_24576 ;
    wire signal_24577 ;
    wire signal_24578 ;
    wire signal_24579 ;
    wire signal_24580 ;
    wire signal_24581 ;
    wire signal_24582 ;
    wire signal_24583 ;
    wire signal_24584 ;
    wire signal_24585 ;
    wire signal_24586 ;
    wire signal_24587 ;
    wire signal_24588 ;
    wire signal_24589 ;
    wire signal_24590 ;
    wire signal_24591 ;
    wire signal_24592 ;
    wire signal_24593 ;
    wire signal_24594 ;
    wire signal_24595 ;
    wire signal_24596 ;
    wire signal_24597 ;
    wire signal_24598 ;
    wire signal_24599 ;
    wire signal_24600 ;
    wire signal_24601 ;
    wire signal_24602 ;
    wire signal_24603 ;
    wire signal_24604 ;
    wire signal_24605 ;
    wire signal_24606 ;
    wire signal_24607 ;
    wire signal_24608 ;
    wire signal_24609 ;
    wire signal_24610 ;
    wire signal_24611 ;
    wire signal_24612 ;
    wire signal_24613 ;
    wire signal_24614 ;
    wire signal_24615 ;
    wire signal_24616 ;
    wire signal_24617 ;
    wire signal_24618 ;
    wire signal_24619 ;
    wire signal_24620 ;
    wire signal_24621 ;
    wire signal_24622 ;
    wire signal_24623 ;
    wire signal_24624 ;
    wire signal_24625 ;
    wire signal_24626 ;
    wire signal_24627 ;
    wire signal_24628 ;
    wire signal_24629 ;
    wire signal_24630 ;
    wire signal_24631 ;
    wire signal_24632 ;
    wire signal_24633 ;
    wire signal_24634 ;
    wire signal_24635 ;
    wire signal_24636 ;
    wire signal_24637 ;
    wire signal_24638 ;
    wire signal_24639 ;
    wire signal_24640 ;
    wire signal_24641 ;
    wire signal_24642 ;
    wire signal_24643 ;
    wire signal_24644 ;
    wire signal_24645 ;
    wire signal_24646 ;
    wire signal_24647 ;
    wire signal_24648 ;
    wire signal_24649 ;
    wire signal_24650 ;
    wire signal_24651 ;
    wire signal_24652 ;
    wire signal_24653 ;
    wire signal_24654 ;
    wire signal_24655 ;
    wire signal_24656 ;
    wire signal_24657 ;
    wire signal_24658 ;
    wire signal_24659 ;
    wire signal_24660 ;
    wire signal_24661 ;
    wire signal_24662 ;
    wire signal_24663 ;
    wire signal_24664 ;
    wire signal_24665 ;
    wire signal_24666 ;
    wire signal_24667 ;
    wire signal_24668 ;
    wire signal_24669 ;
    wire signal_24670 ;
    wire signal_24671 ;
    wire signal_24672 ;
    wire signal_24673 ;
    wire signal_24674 ;
    wire signal_24675 ;
    wire signal_24676 ;
    wire signal_24677 ;
    wire signal_24678 ;
    wire signal_24679 ;
    wire signal_24680 ;
    wire signal_24681 ;
    wire signal_24682 ;
    wire signal_24683 ;
    wire signal_24684 ;
    wire signal_24685 ;
    wire signal_24686 ;
    wire signal_24687 ;
    wire signal_24688 ;
    wire signal_24689 ;
    wire signal_24690 ;
    wire signal_24691 ;
    wire signal_24692 ;
    wire signal_24693 ;
    wire signal_24694 ;
    wire signal_24695 ;
    wire signal_24696 ;
    wire signal_24697 ;
    wire signal_24698 ;
    wire signal_24699 ;
    wire signal_24700 ;
    wire signal_24701 ;
    wire signal_24702 ;
    wire signal_24703 ;
    wire signal_24704 ;
    wire signal_24705 ;
    wire signal_24706 ;
    wire signal_24707 ;
    wire signal_24708 ;
    wire signal_24709 ;
    wire signal_24710 ;
    wire signal_24711 ;
    wire signal_24712 ;
    wire signal_24713 ;
    wire signal_24714 ;
    wire signal_24715 ;
    wire signal_24716 ;
    wire signal_24717 ;
    wire signal_24718 ;
    wire signal_24719 ;
    wire signal_24720 ;
    wire signal_24721 ;
    wire signal_24722 ;
    wire signal_24723 ;
    wire signal_24724 ;
    wire signal_24725 ;
    wire signal_24726 ;
    wire signal_24727 ;
    wire signal_24728 ;
    wire signal_24729 ;
    wire signal_24730 ;
    wire signal_24731 ;
    wire signal_24732 ;
    wire signal_24733 ;
    wire signal_24734 ;
    wire signal_24735 ;
    wire signal_24736 ;
    wire signal_24737 ;
    wire signal_24738 ;
    wire signal_24739 ;
    wire signal_24740 ;
    wire signal_24741 ;
    wire signal_24742 ;
    wire signal_24743 ;
    wire signal_24744 ;
    wire signal_24745 ;
    wire signal_24746 ;
    wire signal_24747 ;
    wire signal_24748 ;
    wire signal_24749 ;
    wire signal_24750 ;
    wire signal_24751 ;
    wire signal_24752 ;
    wire signal_24753 ;
    wire signal_24754 ;
    wire signal_24755 ;
    wire signal_24756 ;
    wire signal_24757 ;
    wire signal_24758 ;
    wire signal_24759 ;
    wire signal_24760 ;
    wire signal_24761 ;
    wire signal_24762 ;
    wire signal_24763 ;
    wire signal_24764 ;
    wire signal_24765 ;
    wire signal_24766 ;
    wire signal_24767 ;
    wire signal_24768 ;
    wire signal_24769 ;
    wire signal_24770 ;
    wire signal_24771 ;
    wire signal_24772 ;
    wire signal_24773 ;
    wire signal_24774 ;
    wire signal_24775 ;
    wire signal_24776 ;
    wire signal_24777 ;
    wire signal_24778 ;
    wire signal_24779 ;
    wire signal_24780 ;
    wire signal_24781 ;
    wire signal_24782 ;
    wire signal_24783 ;
    wire signal_24784 ;
    wire signal_24785 ;
    wire signal_24786 ;
    wire signal_24787 ;
    wire signal_24788 ;
    wire signal_24789 ;
    wire signal_24790 ;
    wire signal_24791 ;
    wire signal_24792 ;
    wire signal_24793 ;
    wire signal_24794 ;
    wire signal_24795 ;
    wire signal_24796 ;
    wire signal_24797 ;
    wire signal_24798 ;
    wire signal_24799 ;
    wire signal_24800 ;
    wire signal_24801 ;
    wire signal_24802 ;
    wire signal_24803 ;
    wire signal_24804 ;
    wire signal_24805 ;
    wire signal_24806 ;
    wire signal_24807 ;
    wire signal_24808 ;
    wire signal_24809 ;
    wire signal_24810 ;
    wire signal_24811 ;
    wire signal_24812 ;
    wire signal_24813 ;
    wire signal_24814 ;
    wire signal_24815 ;
    wire signal_24816 ;
    wire signal_24817 ;
    wire signal_24818 ;
    wire signal_24819 ;
    wire signal_24820 ;
    wire signal_24821 ;
    wire signal_24822 ;
    wire signal_24823 ;
    wire signal_24824 ;
    wire signal_24825 ;
    wire signal_24826 ;
    wire signal_24827 ;
    wire signal_24828 ;
    wire signal_24829 ;
    wire signal_24830 ;
    wire signal_24831 ;
    wire signal_24832 ;
    wire signal_24833 ;
    wire signal_24834 ;
    wire signal_24835 ;
    wire signal_24836 ;
    wire signal_24837 ;
    wire signal_24838 ;
    wire signal_24839 ;
    wire signal_24840 ;
    wire signal_24841 ;
    wire signal_24842 ;
    wire signal_24843 ;
    wire signal_24844 ;
    wire signal_24845 ;
    wire signal_24846 ;
    wire signal_24847 ;
    wire signal_24848 ;
    wire signal_24849 ;
    wire signal_24850 ;
    wire signal_24851 ;
    wire signal_24852 ;
    wire signal_24853 ;
    wire signal_24854 ;
    wire signal_24855 ;
    wire signal_24856 ;
    wire signal_24857 ;
    wire signal_24858 ;
    wire signal_24859 ;
    wire signal_24860 ;
    wire signal_24861 ;
    wire signal_24862 ;
    wire signal_24863 ;
    wire signal_24864 ;
    wire signal_24865 ;
    wire signal_24866 ;
    wire signal_24867 ;
    wire signal_24868 ;
    wire signal_24869 ;
    wire signal_24870 ;
    wire signal_24871 ;
    wire signal_24872 ;
    wire signal_24873 ;
    wire signal_24874 ;
    wire signal_24875 ;
    wire signal_24876 ;
    wire signal_24877 ;
    wire signal_24878 ;
    wire signal_24879 ;
    wire signal_24880 ;
    wire signal_24881 ;
    wire signal_24882 ;
    wire signal_24883 ;
    wire signal_24884 ;
    wire signal_24885 ;
    wire signal_24886 ;
    wire signal_24887 ;
    wire signal_24888 ;
    wire signal_24889 ;
    wire signal_24890 ;
    wire signal_24891 ;
    wire signal_24892 ;
    wire signal_24893 ;
    wire signal_24894 ;
    wire signal_24895 ;
    wire signal_24896 ;
    wire signal_24897 ;
    wire signal_24898 ;
    wire signal_24899 ;
    wire signal_24900 ;
    wire signal_24901 ;
    wire signal_24902 ;
    wire signal_24903 ;
    wire signal_24904 ;
    wire signal_24905 ;
    wire signal_24906 ;
    wire signal_24907 ;
    wire signal_24908 ;
    wire signal_24909 ;
    wire signal_24910 ;
    wire signal_24911 ;
    wire signal_24912 ;
    wire signal_24913 ;
    wire signal_24914 ;
    wire signal_24915 ;
    wire signal_24916 ;
    wire signal_24917 ;
    wire signal_24918 ;
    wire signal_24919 ;
    wire signal_24920 ;
    wire signal_24921 ;
    wire signal_24922 ;
    wire signal_24923 ;
    wire signal_24924 ;
    wire signal_24925 ;
    wire signal_24926 ;
    wire signal_24927 ;
    wire signal_24928 ;
    wire signal_24929 ;
    wire signal_24930 ;
    wire signal_24931 ;
    wire signal_24932 ;
    wire signal_24933 ;
    wire signal_24934 ;
    wire signal_24935 ;
    wire signal_24936 ;
    wire signal_24937 ;
    wire signal_24938 ;
    wire signal_24939 ;
    wire signal_24940 ;
    wire signal_24941 ;
    wire signal_24942 ;
    wire signal_24943 ;
    wire signal_24944 ;
    wire signal_24945 ;
    wire signal_24946 ;
    wire signal_24947 ;
    wire signal_24948 ;
    wire signal_24949 ;
    wire signal_24950 ;
    wire signal_24951 ;
    wire signal_24952 ;
    wire signal_24953 ;
    wire signal_24954 ;
    wire signal_24955 ;
    wire signal_24956 ;
    wire signal_24957 ;
    wire signal_24958 ;
    wire signal_24959 ;
    wire signal_24960 ;
    wire signal_24961 ;
    wire signal_24962 ;
    wire signal_24963 ;
    wire signal_24964 ;
    wire signal_24965 ;
    wire signal_24966 ;
    wire signal_24967 ;
    wire signal_24968 ;
    wire signal_24969 ;
    wire signal_24970 ;
    wire signal_24971 ;
    wire signal_24972 ;
    wire signal_24973 ;
    wire signal_24974 ;
    wire signal_24975 ;
    wire signal_24976 ;
    wire signal_24977 ;
    wire signal_24978 ;
    wire signal_24979 ;
    wire signal_24980 ;
    wire signal_24981 ;
    wire signal_24982 ;
    wire signal_24983 ;
    wire signal_24984 ;
    wire signal_24985 ;
    wire signal_24986 ;
    wire signal_24987 ;
    wire signal_24988 ;
    wire signal_24989 ;
    wire signal_24990 ;
    wire signal_24991 ;
    wire signal_24992 ;
    wire signal_24993 ;
    wire signal_24994 ;
    wire signal_24995 ;
    wire signal_24996 ;
    wire signal_24997 ;
    wire signal_24998 ;
    wire signal_24999 ;
    wire signal_25000 ;
    wire signal_25001 ;
    wire signal_25002 ;
    wire signal_25003 ;
    wire signal_25004 ;
    wire signal_25005 ;
    wire signal_25006 ;
    wire signal_25007 ;
    wire signal_25008 ;
    wire signal_25009 ;
    wire signal_25010 ;
    wire signal_25011 ;
    wire signal_25012 ;
    wire signal_25013 ;
    wire signal_25014 ;
    wire signal_25015 ;
    wire signal_25016 ;
    wire signal_25017 ;
    wire signal_25018 ;
    wire signal_25019 ;
    wire signal_25020 ;
    wire signal_25021 ;
    wire signal_25022 ;
    wire signal_25023 ;
    wire signal_25024 ;
    wire signal_25025 ;
    wire signal_25026 ;
    wire signal_25027 ;
    wire signal_25028 ;
    wire signal_25029 ;
    wire signal_25030 ;
    wire signal_25031 ;
    wire signal_25032 ;
    wire signal_25033 ;
    wire signal_25034 ;
    wire signal_25035 ;
    wire signal_25036 ;
    wire signal_25037 ;
    wire signal_25038 ;
    wire signal_25039 ;
    wire signal_25040 ;
    wire signal_25041 ;
    wire signal_25042 ;
    wire signal_25043 ;
    wire signal_25044 ;
    wire signal_25045 ;
    wire signal_25046 ;
    wire signal_25047 ;
    wire signal_25048 ;
    wire signal_25049 ;
    wire signal_25050 ;
    wire signal_25051 ;
    wire signal_25052 ;
    wire signal_25053 ;
    wire signal_25054 ;
    wire signal_25055 ;
    wire signal_25056 ;
    wire signal_25057 ;
    wire signal_25058 ;
    wire signal_25059 ;
    wire signal_25060 ;
    wire signal_25061 ;
    wire signal_25062 ;
    wire signal_25063 ;
    wire signal_25064 ;
    wire signal_25065 ;
    wire signal_25066 ;
    wire signal_25067 ;
    wire signal_25068 ;
    wire signal_25069 ;
    wire signal_25070 ;
    wire signal_25071 ;
    wire signal_25072 ;
    wire signal_25073 ;
    wire signal_25074 ;
    wire signal_25075 ;
    wire signal_25076 ;
    wire signal_25077 ;
    wire signal_25078 ;
    wire signal_25079 ;
    wire signal_25080 ;
    wire signal_25081 ;
    wire signal_25082 ;
    wire signal_25083 ;
    wire signal_25084 ;
    wire signal_25085 ;
    wire signal_25086 ;
    wire signal_25087 ;
    wire signal_25088 ;
    wire signal_25089 ;
    wire signal_25090 ;
    wire signal_25091 ;
    wire signal_25092 ;
    wire signal_25093 ;
    wire signal_25094 ;
    wire signal_25095 ;
    wire signal_25096 ;
    wire signal_25097 ;
    wire signal_25098 ;
    wire signal_25099 ;
    wire signal_25100 ;
    wire signal_25101 ;
    wire signal_25102 ;
    wire signal_25103 ;
    wire signal_25104 ;
    wire signal_25105 ;
    wire signal_25106 ;
    wire signal_25107 ;
    wire signal_25108 ;
    wire signal_25109 ;
    wire signal_25110 ;
    wire signal_25111 ;
    wire signal_25112 ;
    wire signal_25113 ;
    wire signal_25114 ;
    wire signal_25115 ;
    wire signal_25116 ;
    wire signal_25117 ;
    wire signal_25118 ;
    wire signal_25119 ;
    wire signal_25120 ;
    wire signal_25121 ;
    wire signal_25122 ;
    wire signal_25123 ;
    wire signal_25124 ;
    wire signal_25125 ;
    wire signal_25126 ;
    wire signal_25127 ;
    wire signal_25128 ;
    wire signal_25129 ;
    wire signal_25130 ;
    wire signal_25131 ;
    wire signal_25132 ;
    wire signal_25133 ;
    wire signal_25134 ;
    wire signal_25135 ;
    wire signal_25136 ;
    wire signal_25137 ;
    wire signal_25138 ;
    wire signal_25139 ;
    wire signal_25140 ;
    wire signal_25141 ;
    wire signal_25142 ;
    wire signal_25143 ;
    wire signal_25144 ;
    wire signal_25145 ;
    wire signal_25146 ;
    wire signal_25147 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) cell_927 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2399, signal_2398, signal_2397, signal_2396, signal_942}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_928 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2407, signal_2406, signal_2405, signal_2404, signal_943}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_929 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_930 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_931 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_932 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_933 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_934 ( .a ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2455, signal_2454, signal_2453, signal_2452, signal_949}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_949 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .c ({signal_2515, signal_2514, signal_2513, signal_2512, signal_964}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_950 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .c ({signal_2519, signal_2518, signal_2517, signal_2516, signal_965}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_962 ( .a ({signal_2515, signal_2514, signal_2513, signal_2512, signal_964}), .b ({signal_2567, signal_2566, signal_2565, signal_2564, signal_977}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_963 ( .a ({signal_2519, signal_2518, signal_2517, signal_2516, signal_965}), .b ({signal_2571, signal_2570, signal_2569, signal_2568, signal_978}) ) ;

    /* cells in depth 1 */
    buf_clk cell_2385 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( signal_17078 ) ) ;
    buf_clk cell_2387 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( signal_17080 ) ) ;
    buf_clk cell_2389 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( signal_17082 ) ) ;
    buf_clk cell_2391 ( .C ( clk ), .D ( SI_s3[6] ), .Q ( signal_17084 ) ) ;
    buf_clk cell_2393 ( .C ( clk ), .D ( SI_s4[6] ), .Q ( signal_17086 ) ) ;
    buf_clk cell_2395 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_17088 ) ) ;
    buf_clk cell_2397 ( .C ( clk ), .D ( signal_2452 ), .Q ( signal_17090 ) ) ;
    buf_clk cell_2399 ( .C ( clk ), .D ( signal_2453 ), .Q ( signal_17092 ) ) ;
    buf_clk cell_2401 ( .C ( clk ), .D ( signal_2454 ), .Q ( signal_17094 ) ) ;
    buf_clk cell_2403 ( .C ( clk ), .D ( signal_2455 ), .Q ( signal_17096 ) ) ;
    buf_clk cell_2405 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_17098 ) ) ;
    buf_clk cell_2407 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_17100 ) ) ;
    buf_clk cell_2409 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_17102 ) ) ;
    buf_clk cell_2411 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( signal_17104 ) ) ;
    buf_clk cell_2413 ( .C ( clk ), .D ( SI_s4[0] ), .Q ( signal_17106 ) ) ;
    buf_clk cell_2415 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_17108 ) ) ;
    buf_clk cell_2417 ( .C ( clk ), .D ( signal_2412 ), .Q ( signal_17110 ) ) ;
    buf_clk cell_2419 ( .C ( clk ), .D ( signal_2413 ), .Q ( signal_17112 ) ) ;
    buf_clk cell_2421 ( .C ( clk ), .D ( signal_2414 ), .Q ( signal_17114 ) ) ;
    buf_clk cell_2423 ( .C ( clk ), .D ( signal_2415 ), .Q ( signal_17116 ) ) ;
    buf_clk cell_2425 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_17118 ) ) ;
    buf_clk cell_2427 ( .C ( clk ), .D ( signal_2396 ), .Q ( signal_17120 ) ) ;
    buf_clk cell_2429 ( .C ( clk ), .D ( signal_2397 ), .Q ( signal_17122 ) ) ;
    buf_clk cell_2431 ( .C ( clk ), .D ( signal_2398 ), .Q ( signal_17124 ) ) ;
    buf_clk cell_2433 ( .C ( clk ), .D ( signal_2399 ), .Q ( signal_17126 ) ) ;
    buf_clk cell_2435 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_17128 ) ) ;
    buf_clk cell_2437 ( .C ( clk ), .D ( signal_2428 ), .Q ( signal_17130 ) ) ;
    buf_clk cell_2439 ( .C ( clk ), .D ( signal_2429 ), .Q ( signal_17132 ) ) ;
    buf_clk cell_2441 ( .C ( clk ), .D ( signal_2430 ), .Q ( signal_17134 ) ) ;
    buf_clk cell_2443 ( .C ( clk ), .D ( signal_2431 ), .Q ( signal_17136 ) ) ;
    buf_clk cell_2445 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_17138 ) ) ;
    buf_clk cell_2447 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_17140 ) ) ;
    buf_clk cell_2449 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_17142 ) ) ;
    buf_clk cell_2451 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( signal_17144 ) ) ;
    buf_clk cell_2453 ( .C ( clk ), .D ( SI_s4[1] ), .Q ( signal_17146 ) ) ;
    buf_clk cell_2455 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( signal_17148 ) ) ;
    buf_clk cell_2457 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( signal_17150 ) ) ;
    buf_clk cell_2459 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( signal_17152 ) ) ;
    buf_clk cell_2461 ( .C ( clk ), .D ( SI_s3[4] ), .Q ( signal_17154 ) ) ;
    buf_clk cell_2463 ( .C ( clk ), .D ( SI_s4[4] ), .Q ( signal_17156 ) ) ;
    buf_clk cell_2465 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_17158 ) ) ;
    buf_clk cell_2467 ( .C ( clk ), .D ( signal_2420 ), .Q ( signal_17160 ) ) ;
    buf_clk cell_2469 ( .C ( clk ), .D ( signal_2421 ), .Q ( signal_17162 ) ) ;
    buf_clk cell_2471 ( .C ( clk ), .D ( signal_2422 ), .Q ( signal_17164 ) ) ;
    buf_clk cell_2473 ( .C ( clk ), .D ( signal_2423 ), .Q ( signal_17166 ) ) ;
    buf_clk cell_2475 ( .C ( clk ), .D ( signal_948 ), .Q ( signal_17168 ) ) ;
    buf_clk cell_2477 ( .C ( clk ), .D ( signal_2444 ), .Q ( signal_17170 ) ) ;
    buf_clk cell_2479 ( .C ( clk ), .D ( signal_2445 ), .Q ( signal_17172 ) ) ;
    buf_clk cell_2481 ( .C ( clk ), .D ( signal_2446 ), .Q ( signal_17174 ) ) ;
    buf_clk cell_2483 ( .C ( clk ), .D ( signal_2447 ), .Q ( signal_17176 ) ) ;
    buf_clk cell_2485 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( signal_17178 ) ) ;
    buf_clk cell_2487 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( signal_17180 ) ) ;
    buf_clk cell_2489 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( signal_17182 ) ) ;
    buf_clk cell_2491 ( .C ( clk ), .D ( SI_s3[5] ), .Q ( signal_17184 ) ) ;
    buf_clk cell_2493 ( .C ( clk ), .D ( SI_s4[5] ), .Q ( signal_17186 ) ) ;
    buf_clk cell_2495 ( .C ( clk ), .D ( signal_978 ), .Q ( signal_17188 ) ) ;
    buf_clk cell_2497 ( .C ( clk ), .D ( signal_2568 ), .Q ( signal_17190 ) ) ;
    buf_clk cell_2499 ( .C ( clk ), .D ( signal_2569 ), .Q ( signal_17192 ) ) ;
    buf_clk cell_2501 ( .C ( clk ), .D ( signal_2570 ), .Q ( signal_17194 ) ) ;
    buf_clk cell_2503 ( .C ( clk ), .D ( signal_2571 ), .Q ( signal_17196 ) ) ;
    buf_clk cell_2505 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_17198 ) ) ;
    buf_clk cell_2507 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_17200 ) ) ;
    buf_clk cell_2509 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_17202 ) ) ;
    buf_clk cell_2511 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( signal_17204 ) ) ;
    buf_clk cell_2513 ( .C ( clk ), .D ( SI_s4[2] ), .Q ( signal_17206 ) ) ;
    buf_clk cell_2515 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_17208 ) ) ;
    buf_clk cell_2519 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_17212 ) ) ;
    buf_clk cell_2523 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_17216 ) ) ;
    buf_clk cell_2527 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( signal_17220 ) ) ;
    buf_clk cell_2531 ( .C ( clk ), .D ( SI_s4[3] ), .Q ( signal_17224 ) ) ;
    buf_clk cell_2875 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_17568 ) ) ;
    buf_clk cell_2879 ( .C ( clk ), .D ( signal_2404 ), .Q ( signal_17572 ) ) ;
    buf_clk cell_2883 ( .C ( clk ), .D ( signal_2405 ), .Q ( signal_17576 ) ) ;
    buf_clk cell_2887 ( .C ( clk ), .D ( signal_2406 ), .Q ( signal_17580 ) ) ;
    buf_clk cell_2891 ( .C ( clk ), .D ( signal_2407 ), .Q ( signal_17584 ) ) ;
    buf_clk cell_3225 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( signal_17918 ) ) ;
    buf_clk cell_3231 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( signal_17924 ) ) ;
    buf_clk cell_3237 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( signal_17930 ) ) ;
    buf_clk cell_3243 ( .C ( clk ), .D ( SI_s3[7] ), .Q ( signal_17936 ) ) ;
    buf_clk cell_3249 ( .C ( clk ), .D ( SI_s4[7] ), .Q ( signal_17942 ) ) ;
    buf_clk cell_3705 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_18398 ) ) ;
    buf_clk cell_3711 ( .C ( clk ), .D ( signal_2436 ), .Q ( signal_18404 ) ) ;
    buf_clk cell_3717 ( .C ( clk ), .D ( signal_2437 ), .Q ( signal_18410 ) ) ;
    buf_clk cell_3723 ( .C ( clk ), .D ( signal_2438 ), .Q ( signal_18416 ) ) ;
    buf_clk cell_3729 ( .C ( clk ), .D ( signal_2439 ), .Q ( signal_18422 ) ) ;
    buf_clk cell_4075 ( .C ( clk ), .D ( signal_977 ), .Q ( signal_18768 ) ) ;
    buf_clk cell_4083 ( .C ( clk ), .D ( signal_2564 ), .Q ( signal_18776 ) ) ;
    buf_clk cell_4091 ( .C ( clk ), .D ( signal_2565 ), .Q ( signal_18784 ) ) ;
    buf_clk cell_4099 ( .C ( clk ), .D ( signal_2566 ), .Q ( signal_18792 ) ) ;
    buf_clk cell_4107 ( .C ( clk ), .D ( signal_2567 ), .Q ( signal_18800 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_935 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_2459, signal_2458, signal_2457, signal_2456, signal_950}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_936 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_937 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_938 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_939 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_2475, signal_2474, signal_2473, signal_2472, signal_954}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_940 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_2479, signal_2478, signal_2477, signal_2476, signal_955}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_941 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_2483, signal_2482, signal_2481, signal_2480, signal_956}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_942 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_943 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_2491, signal_2490, signal_2489, signal_2488, signal_958}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_944 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_2495, signal_2494, signal_2493, signal_2492, signal_959}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_945 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_946 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_947 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_948 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_2511, signal_2510, signal_2509, signal_2508, signal_963}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_951 ( .a ({signal_2459, signal_2458, signal_2457, signal_2456, signal_950}), .b ({signal_2523, signal_2522, signal_2521, signal_2520, signal_966}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_952 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2527, signal_2526, signal_2525, signal_2524, signal_967}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_953 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2531, signal_2530, signal_2529, signal_2528, signal_968}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_954 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2535, signal_2534, signal_2533, signal_2532, signal_969}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_955 ( .a ({signal_2475, signal_2474, signal_2473, signal_2472, signal_954}), .b ({signal_2539, signal_2538, signal_2537, signal_2536, signal_970}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_956 ( .a ({signal_2483, signal_2482, signal_2481, signal_2480, signal_956}), .b ({signal_2543, signal_2542, signal_2541, signal_2540, signal_971}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_957 ( .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .b ({signal_2547, signal_2546, signal_2545, signal_2544, signal_972}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_958 ( .a ({signal_2495, signal_2494, signal_2493, signal_2492, signal_959}), .b ({signal_2551, signal_2550, signal_2549, signal_2548, signal_973}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_959 ( .a ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}), .b ({signal_2555, signal_2554, signal_2553, signal_2552, signal_974}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_960 ( .a ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .b ({signal_2559, signal_2558, signal_2557, signal_2556, signal_975}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_961 ( .a ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .b ({signal_2563, signal_2562, signal_2561, signal_2560, signal_976}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_964 ( .a ({signal_2407, signal_2406, signal_2405, signal_2404, signal_943}), .b ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_965 ( .a ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}), .b ({signal_2455, signal_2454, signal_2453, signal_2452, signal_949}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_966 ( .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .clk ( clk ), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_967 ( .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_2587, signal_2586, signal_2585, signal_2584, signal_982}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_968 ( .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .b ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .clk ( clk ), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_969 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2407, signal_2406, signal_2405, signal_2404, signal_943}), .clk ( clk ), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_970 ( .a ({signal_2399, signal_2398, signal_2397, signal_2396, signal_942}), .b ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_971 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .clk ( clk ), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_972 ( .a ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .b ({signal_2455, signal_2454, signal_2453, signal_2452, signal_949}), .clk ( clk ), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_2607, signal_2606, signal_2605, signal_2604, signal_987}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_973 ( .a ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .b ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_974 ( .a ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .b ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_975 ( .a ({signal_2407, signal_2406, signal_2405, signal_2404, signal_943}), .b ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_976 ( .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .b ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_977 ( .a ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_978 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .clk ( clk ), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_979 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_980 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .clk ( clk ), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_981 ( .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .b ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_982 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_983 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2455, signal_2454, signal_2453, signal_2452, signal_949}), .clk ( clk ), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_984 ( .a ({signal_2399, signal_2398, signal_2397, signal_2396, signal_942}), .b ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({signal_2655, signal_2654, signal_2653, signal_2652, signal_999}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_985 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .c ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_986 ( .a ({signal_2399, signal_2398, signal_2397, signal_2396, signal_942}), .b ({signal_2407, signal_2406, signal_2405, signal_2404, signal_943}), .clk ( clk ), .r ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_987 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .clk ( clk ), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .c ({signal_2667, signal_2666, signal_2665, signal_2664, signal_1002}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_989 ( .a ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_990 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .clk ( clk ), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_991 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .clk ( clk ), .r ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .c ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1006}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_992 ( .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .b ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .c ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_993 ( .a ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_994 ( .a ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .b ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .clk ( clk ), .r ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .c ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_995 ( .a ({signal_2399, signal_2398, signal_2397, signal_2396, signal_942}), .b ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .c ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1010}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_996 ( .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_944}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_2703, signal_2702, signal_2701, signal_2700, signal_1011}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_997 ( .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .b ({signal_2439, signal_2438, signal_2437, signal_2436, signal_947}), .clk ( clk ), .r ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .c ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1012}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_998 ( .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .c ({signal_2711, signal_2710, signal_2709, signal_2708, signal_1013}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1000 ( .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_945}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1015}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1001 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2447, signal_2446, signal_2445, signal_2444, signal_948}), .clk ( clk ), .r ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .c ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1016}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1002 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2431, signal_2430, signal_2429, signal_2428, signal_946}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .c ({signal_2727, signal_2726, signal_2725, signal_2724, signal_1017}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1003 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2455, signal_2454, signal_2453, signal_2452, signal_949}), .clk ( clk ), .r ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_2731, signal_2730, signal_2729, signal_2728, signal_1018}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1016 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_2783, signal_2782, signal_2781, signal_2780, signal_1031}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1017 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2787, signal_2786, signal_2785, signal_2784, signal_1032}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1018 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2791, signal_2790, signal_2789, signal_2788, signal_1033}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1019 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2795, signal_2794, signal_2793, signal_2792, signal_1034}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1020 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2799, signal_2798, signal_2797, signal_2796, signal_1035}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1021 ( .a ({signal_2607, signal_2606, signal_2605, signal_2604, signal_987}), .b ({signal_2803, signal_2802, signal_2801, signal_2800, signal_1036}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1022 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2807, signal_2806, signal_2805, signal_2804, signal_1037}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1023 ( .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .b ({signal_2811, signal_2810, signal_2809, signal_2808, signal_1038}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1024 ( .a ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}), .b ({signal_2815, signal_2814, signal_2813, signal_2812, signal_1039}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1025 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2819, signal_2818, signal_2817, signal_2816, signal_1040}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1026 ( .a ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .b ({signal_2823, signal_2822, signal_2821, signal_2820, signal_1041}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1027 ( .a ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .b ({signal_2827, signal_2826, signal_2825, signal_2824, signal_1042}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1028 ( .a ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}), .b ({signal_2831, signal_2830, signal_2829, signal_2828, signal_1043}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1029 ( .a ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .b ({signal_2835, signal_2834, signal_2833, signal_2832, signal_1044}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1030 ( .a ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .b ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1031 ( .a ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}), .b ({signal_2843, signal_2842, signal_2841, signal_2840, signal_1046}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1032 ( .a ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .b ({signal_2847, signal_2846, signal_2845, signal_2844, signal_1047}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1034 ( .a ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .b ({signal_2855, signal_2854, signal_2853, signal_2852, signal_1049}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1035 ( .a ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .b ({signal_2859, signal_2858, signal_2857, signal_2856, signal_1050}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1036 ( .a ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1006}), .b ({signal_2863, signal_2862, signal_2861, signal_2860, signal_1051}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1037 ( .a ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}), .b ({signal_2867, signal_2866, signal_2865, signal_2864, signal_1052}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1038 ( .a ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .b ({signal_2871, signal_2870, signal_2869, signal_2868, signal_1053}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1039 ( .a ({signal_2711, signal_2710, signal_2709, signal_2708, signal_1013}), .b ({signal_2875, signal_2874, signal_2873, signal_2872, signal_1054}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1041 ( .a ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1015}), .b ({signal_2883, signal_2882, signal_2881, signal_2880, signal_1056}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1042 ( .a ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1016}), .b ({signal_2887, signal_2886, signal_2885, signal_2884, signal_1057}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1043 ( .a ({signal_2727, signal_2726, signal_2725, signal_2724, signal_1017}), .b ({signal_2891, signal_2890, signal_2889, signal_2888, signal_1058}) ) ;
    buf_clk cell_2386 ( .C ( clk ), .D ( signal_17078 ), .Q ( signal_17079 ) ) ;
    buf_clk cell_2388 ( .C ( clk ), .D ( signal_17080 ), .Q ( signal_17081 ) ) ;
    buf_clk cell_2390 ( .C ( clk ), .D ( signal_17082 ), .Q ( signal_17083 ) ) ;
    buf_clk cell_2392 ( .C ( clk ), .D ( signal_17084 ), .Q ( signal_17085 ) ) ;
    buf_clk cell_2394 ( .C ( clk ), .D ( signal_17086 ), .Q ( signal_17087 ) ) ;
    buf_clk cell_2396 ( .C ( clk ), .D ( signal_17088 ), .Q ( signal_17089 ) ) ;
    buf_clk cell_2398 ( .C ( clk ), .D ( signal_17090 ), .Q ( signal_17091 ) ) ;
    buf_clk cell_2400 ( .C ( clk ), .D ( signal_17092 ), .Q ( signal_17093 ) ) ;
    buf_clk cell_2402 ( .C ( clk ), .D ( signal_17094 ), .Q ( signal_17095 ) ) ;
    buf_clk cell_2404 ( .C ( clk ), .D ( signal_17096 ), .Q ( signal_17097 ) ) ;
    buf_clk cell_2406 ( .C ( clk ), .D ( signal_17098 ), .Q ( signal_17099 ) ) ;
    buf_clk cell_2408 ( .C ( clk ), .D ( signal_17100 ), .Q ( signal_17101 ) ) ;
    buf_clk cell_2410 ( .C ( clk ), .D ( signal_17102 ), .Q ( signal_17103 ) ) ;
    buf_clk cell_2412 ( .C ( clk ), .D ( signal_17104 ), .Q ( signal_17105 ) ) ;
    buf_clk cell_2414 ( .C ( clk ), .D ( signal_17106 ), .Q ( signal_17107 ) ) ;
    buf_clk cell_2416 ( .C ( clk ), .D ( signal_17108 ), .Q ( signal_17109 ) ) ;
    buf_clk cell_2418 ( .C ( clk ), .D ( signal_17110 ), .Q ( signal_17111 ) ) ;
    buf_clk cell_2420 ( .C ( clk ), .D ( signal_17112 ), .Q ( signal_17113 ) ) ;
    buf_clk cell_2422 ( .C ( clk ), .D ( signal_17114 ), .Q ( signal_17115 ) ) ;
    buf_clk cell_2424 ( .C ( clk ), .D ( signal_17116 ), .Q ( signal_17117 ) ) ;
    buf_clk cell_2426 ( .C ( clk ), .D ( signal_17118 ), .Q ( signal_17119 ) ) ;
    buf_clk cell_2428 ( .C ( clk ), .D ( signal_17120 ), .Q ( signal_17121 ) ) ;
    buf_clk cell_2430 ( .C ( clk ), .D ( signal_17122 ), .Q ( signal_17123 ) ) ;
    buf_clk cell_2432 ( .C ( clk ), .D ( signal_17124 ), .Q ( signal_17125 ) ) ;
    buf_clk cell_2434 ( .C ( clk ), .D ( signal_17126 ), .Q ( signal_17127 ) ) ;
    buf_clk cell_2436 ( .C ( clk ), .D ( signal_17128 ), .Q ( signal_17129 ) ) ;
    buf_clk cell_2438 ( .C ( clk ), .D ( signal_17130 ), .Q ( signal_17131 ) ) ;
    buf_clk cell_2440 ( .C ( clk ), .D ( signal_17132 ), .Q ( signal_17133 ) ) ;
    buf_clk cell_2442 ( .C ( clk ), .D ( signal_17134 ), .Q ( signal_17135 ) ) ;
    buf_clk cell_2444 ( .C ( clk ), .D ( signal_17136 ), .Q ( signal_17137 ) ) ;
    buf_clk cell_2446 ( .C ( clk ), .D ( signal_17138 ), .Q ( signal_17139 ) ) ;
    buf_clk cell_2448 ( .C ( clk ), .D ( signal_17140 ), .Q ( signal_17141 ) ) ;
    buf_clk cell_2450 ( .C ( clk ), .D ( signal_17142 ), .Q ( signal_17143 ) ) ;
    buf_clk cell_2452 ( .C ( clk ), .D ( signal_17144 ), .Q ( signal_17145 ) ) ;
    buf_clk cell_2454 ( .C ( clk ), .D ( signal_17146 ), .Q ( signal_17147 ) ) ;
    buf_clk cell_2456 ( .C ( clk ), .D ( signal_17148 ), .Q ( signal_17149 ) ) ;
    buf_clk cell_2458 ( .C ( clk ), .D ( signal_17150 ), .Q ( signal_17151 ) ) ;
    buf_clk cell_2460 ( .C ( clk ), .D ( signal_17152 ), .Q ( signal_17153 ) ) ;
    buf_clk cell_2462 ( .C ( clk ), .D ( signal_17154 ), .Q ( signal_17155 ) ) ;
    buf_clk cell_2464 ( .C ( clk ), .D ( signal_17156 ), .Q ( signal_17157 ) ) ;
    buf_clk cell_2466 ( .C ( clk ), .D ( signal_17158 ), .Q ( signal_17159 ) ) ;
    buf_clk cell_2468 ( .C ( clk ), .D ( signal_17160 ), .Q ( signal_17161 ) ) ;
    buf_clk cell_2470 ( .C ( clk ), .D ( signal_17162 ), .Q ( signal_17163 ) ) ;
    buf_clk cell_2472 ( .C ( clk ), .D ( signal_17164 ), .Q ( signal_17165 ) ) ;
    buf_clk cell_2474 ( .C ( clk ), .D ( signal_17166 ), .Q ( signal_17167 ) ) ;
    buf_clk cell_2476 ( .C ( clk ), .D ( signal_17168 ), .Q ( signal_17169 ) ) ;
    buf_clk cell_2478 ( .C ( clk ), .D ( signal_17170 ), .Q ( signal_17171 ) ) ;
    buf_clk cell_2480 ( .C ( clk ), .D ( signal_17172 ), .Q ( signal_17173 ) ) ;
    buf_clk cell_2482 ( .C ( clk ), .D ( signal_17174 ), .Q ( signal_17175 ) ) ;
    buf_clk cell_2484 ( .C ( clk ), .D ( signal_17176 ), .Q ( signal_17177 ) ) ;
    buf_clk cell_2486 ( .C ( clk ), .D ( signal_17178 ), .Q ( signal_17179 ) ) ;
    buf_clk cell_2488 ( .C ( clk ), .D ( signal_17180 ), .Q ( signal_17181 ) ) ;
    buf_clk cell_2490 ( .C ( clk ), .D ( signal_17182 ), .Q ( signal_17183 ) ) ;
    buf_clk cell_2492 ( .C ( clk ), .D ( signal_17184 ), .Q ( signal_17185 ) ) ;
    buf_clk cell_2494 ( .C ( clk ), .D ( signal_17186 ), .Q ( signal_17187 ) ) ;
    buf_clk cell_2496 ( .C ( clk ), .D ( signal_17188 ), .Q ( signal_17189 ) ) ;
    buf_clk cell_2498 ( .C ( clk ), .D ( signal_17190 ), .Q ( signal_17191 ) ) ;
    buf_clk cell_2500 ( .C ( clk ), .D ( signal_17192 ), .Q ( signal_17193 ) ) ;
    buf_clk cell_2502 ( .C ( clk ), .D ( signal_17194 ), .Q ( signal_17195 ) ) ;
    buf_clk cell_2504 ( .C ( clk ), .D ( signal_17196 ), .Q ( signal_17197 ) ) ;
    buf_clk cell_2506 ( .C ( clk ), .D ( signal_17198 ), .Q ( signal_17199 ) ) ;
    buf_clk cell_2508 ( .C ( clk ), .D ( signal_17200 ), .Q ( signal_17201 ) ) ;
    buf_clk cell_2510 ( .C ( clk ), .D ( signal_17202 ), .Q ( signal_17203 ) ) ;
    buf_clk cell_2512 ( .C ( clk ), .D ( signal_17204 ), .Q ( signal_17205 ) ) ;
    buf_clk cell_2514 ( .C ( clk ), .D ( signal_17206 ), .Q ( signal_17207 ) ) ;
    buf_clk cell_2516 ( .C ( clk ), .D ( signal_17208 ), .Q ( signal_17209 ) ) ;
    buf_clk cell_2520 ( .C ( clk ), .D ( signal_17212 ), .Q ( signal_17213 ) ) ;
    buf_clk cell_2524 ( .C ( clk ), .D ( signal_17216 ), .Q ( signal_17217 ) ) ;
    buf_clk cell_2528 ( .C ( clk ), .D ( signal_17220 ), .Q ( signal_17221 ) ) ;
    buf_clk cell_2532 ( .C ( clk ), .D ( signal_17224 ), .Q ( signal_17225 ) ) ;
    buf_clk cell_2876 ( .C ( clk ), .D ( signal_17568 ), .Q ( signal_17569 ) ) ;
    buf_clk cell_2880 ( .C ( clk ), .D ( signal_17572 ), .Q ( signal_17573 ) ) ;
    buf_clk cell_2884 ( .C ( clk ), .D ( signal_17576 ), .Q ( signal_17577 ) ) ;
    buf_clk cell_2888 ( .C ( clk ), .D ( signal_17580 ), .Q ( signal_17581 ) ) ;
    buf_clk cell_2892 ( .C ( clk ), .D ( signal_17584 ), .Q ( signal_17585 ) ) ;
    buf_clk cell_3226 ( .C ( clk ), .D ( signal_17918 ), .Q ( signal_17919 ) ) ;
    buf_clk cell_3232 ( .C ( clk ), .D ( signal_17924 ), .Q ( signal_17925 ) ) ;
    buf_clk cell_3238 ( .C ( clk ), .D ( signal_17930 ), .Q ( signal_17931 ) ) ;
    buf_clk cell_3244 ( .C ( clk ), .D ( signal_17936 ), .Q ( signal_17937 ) ) ;
    buf_clk cell_3250 ( .C ( clk ), .D ( signal_17942 ), .Q ( signal_17943 ) ) ;
    buf_clk cell_3706 ( .C ( clk ), .D ( signal_18398 ), .Q ( signal_18399 ) ) ;
    buf_clk cell_3712 ( .C ( clk ), .D ( signal_18404 ), .Q ( signal_18405 ) ) ;
    buf_clk cell_3718 ( .C ( clk ), .D ( signal_18410 ), .Q ( signal_18411 ) ) ;
    buf_clk cell_3724 ( .C ( clk ), .D ( signal_18416 ), .Q ( signal_18417 ) ) ;
    buf_clk cell_3730 ( .C ( clk ), .D ( signal_18422 ), .Q ( signal_18423 ) ) ;
    buf_clk cell_4076 ( .C ( clk ), .D ( signal_18768 ), .Q ( signal_18769 ) ) ;
    buf_clk cell_4084 ( .C ( clk ), .D ( signal_18776 ), .Q ( signal_18777 ) ) ;
    buf_clk cell_4092 ( .C ( clk ), .D ( signal_18784 ), .Q ( signal_18785 ) ) ;
    buf_clk cell_4100 ( .C ( clk ), .D ( signal_18792 ), .Q ( signal_18793 ) ) ;
    buf_clk cell_4108 ( .C ( clk ), .D ( signal_18800 ), .Q ( signal_18801 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_2517 ( .C ( clk ), .D ( signal_17209 ), .Q ( signal_17210 ) ) ;
    buf_clk cell_2521 ( .C ( clk ), .D ( signal_17213 ), .Q ( signal_17214 ) ) ;
    buf_clk cell_2525 ( .C ( clk ), .D ( signal_17217 ), .Q ( signal_17218 ) ) ;
    buf_clk cell_2529 ( .C ( clk ), .D ( signal_17221 ), .Q ( signal_17222 ) ) ;
    buf_clk cell_2533 ( .C ( clk ), .D ( signal_17225 ), .Q ( signal_17226 ) ) ;
    buf_clk cell_2535 ( .C ( clk ), .D ( signal_17159 ), .Q ( signal_17228 ) ) ;
    buf_clk cell_2537 ( .C ( clk ), .D ( signal_17161 ), .Q ( signal_17230 ) ) ;
    buf_clk cell_2539 ( .C ( clk ), .D ( signal_17163 ), .Q ( signal_17232 ) ) ;
    buf_clk cell_2541 ( .C ( clk ), .D ( signal_17165 ), .Q ( signal_17234 ) ) ;
    buf_clk cell_2543 ( .C ( clk ), .D ( signal_17167 ), .Q ( signal_17236 ) ) ;
    buf_clk cell_2545 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_17238 ) ) ;
    buf_clk cell_2547 ( .C ( clk ), .D ( signal_2636 ), .Q ( signal_17240 ) ) ;
    buf_clk cell_2549 ( .C ( clk ), .D ( signal_2637 ), .Q ( signal_17242 ) ) ;
    buf_clk cell_2551 ( .C ( clk ), .D ( signal_2638 ), .Q ( signal_17244 ) ) ;
    buf_clk cell_2553 ( .C ( clk ), .D ( signal_2639 ), .Q ( signal_17246 ) ) ;
    buf_clk cell_2555 ( .C ( clk ), .D ( signal_1010 ), .Q ( signal_17248 ) ) ;
    buf_clk cell_2557 ( .C ( clk ), .D ( signal_2696 ), .Q ( signal_17250 ) ) ;
    buf_clk cell_2559 ( .C ( clk ), .D ( signal_2697 ), .Q ( signal_17252 ) ) ;
    buf_clk cell_2561 ( .C ( clk ), .D ( signal_2698 ), .Q ( signal_17254 ) ) ;
    buf_clk cell_2563 ( .C ( clk ), .D ( signal_2699 ), .Q ( signal_17256 ) ) ;
    buf_clk cell_2565 ( .C ( clk ), .D ( signal_992 ), .Q ( signal_17258 ) ) ;
    buf_clk cell_2567 ( .C ( clk ), .D ( signal_2624 ), .Q ( signal_17260 ) ) ;
    buf_clk cell_2569 ( .C ( clk ), .D ( signal_2625 ), .Q ( signal_17262 ) ) ;
    buf_clk cell_2571 ( .C ( clk ), .D ( signal_2626 ), .Q ( signal_17264 ) ) ;
    buf_clk cell_2573 ( .C ( clk ), .D ( signal_2627 ), .Q ( signal_17266 ) ) ;
    buf_clk cell_2575 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_17268 ) ) ;
    buf_clk cell_2577 ( .C ( clk ), .D ( signal_2628 ), .Q ( signal_17270 ) ) ;
    buf_clk cell_2579 ( .C ( clk ), .D ( signal_2629 ), .Q ( signal_17272 ) ) ;
    buf_clk cell_2581 ( .C ( clk ), .D ( signal_2630 ), .Q ( signal_17274 ) ) ;
    buf_clk cell_2583 ( .C ( clk ), .D ( signal_2631 ), .Q ( signal_17276 ) ) ;
    buf_clk cell_2585 ( .C ( clk ), .D ( signal_1008 ), .Q ( signal_17278 ) ) ;
    buf_clk cell_2587 ( .C ( clk ), .D ( signal_2688 ), .Q ( signal_17280 ) ) ;
    buf_clk cell_2589 ( .C ( clk ), .D ( signal_2689 ), .Q ( signal_17282 ) ) ;
    buf_clk cell_2591 ( .C ( clk ), .D ( signal_2690 ), .Q ( signal_17284 ) ) ;
    buf_clk cell_2593 ( .C ( clk ), .D ( signal_2691 ), .Q ( signal_17286 ) ) ;
    buf_clk cell_2595 ( .C ( clk ), .D ( signal_991 ), .Q ( signal_17288 ) ) ;
    buf_clk cell_2597 ( .C ( clk ), .D ( signal_2620 ), .Q ( signal_17290 ) ) ;
    buf_clk cell_2599 ( .C ( clk ), .D ( signal_2621 ), .Q ( signal_17292 ) ) ;
    buf_clk cell_2601 ( .C ( clk ), .D ( signal_2622 ), .Q ( signal_17294 ) ) ;
    buf_clk cell_2603 ( .C ( clk ), .D ( signal_2623 ), .Q ( signal_17296 ) ) ;
    buf_clk cell_2605 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_17298 ) ) ;
    buf_clk cell_2607 ( .C ( clk ), .D ( signal_2492 ), .Q ( signal_17300 ) ) ;
    buf_clk cell_2609 ( .C ( clk ), .D ( signal_2493 ), .Q ( signal_17302 ) ) ;
    buf_clk cell_2611 ( .C ( clk ), .D ( signal_2494 ), .Q ( signal_17304 ) ) ;
    buf_clk cell_2613 ( .C ( clk ), .D ( signal_2495 ), .Q ( signal_17306 ) ) ;
    buf_clk cell_2615 ( .C ( clk ), .D ( signal_987 ), .Q ( signal_17308 ) ) ;
    buf_clk cell_2617 ( .C ( clk ), .D ( signal_2604 ), .Q ( signal_17310 ) ) ;
    buf_clk cell_2619 ( .C ( clk ), .D ( signal_2605 ), .Q ( signal_17312 ) ) ;
    buf_clk cell_2621 ( .C ( clk ), .D ( signal_2606 ), .Q ( signal_17314 ) ) ;
    buf_clk cell_2623 ( .C ( clk ), .D ( signal_2607 ), .Q ( signal_17316 ) ) ;
    buf_clk cell_2625 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_17318 ) ) ;
    buf_clk cell_2627 ( .C ( clk ), .D ( signal_2500 ), .Q ( signal_17320 ) ) ;
    buf_clk cell_2629 ( .C ( clk ), .D ( signal_2501 ), .Q ( signal_17322 ) ) ;
    buf_clk cell_2631 ( .C ( clk ), .D ( signal_2502 ), .Q ( signal_17324 ) ) ;
    buf_clk cell_2633 ( .C ( clk ), .D ( signal_2503 ), .Q ( signal_17326 ) ) ;
    buf_clk cell_2635 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_17328 ) ) ;
    buf_clk cell_2637 ( .C ( clk ), .D ( signal_2572 ), .Q ( signal_17330 ) ) ;
    buf_clk cell_2639 ( .C ( clk ), .D ( signal_2573 ), .Q ( signal_17332 ) ) ;
    buf_clk cell_2641 ( .C ( clk ), .D ( signal_2574 ), .Q ( signal_17334 ) ) ;
    buf_clk cell_2643 ( .C ( clk ), .D ( signal_2575 ), .Q ( signal_17336 ) ) ;
    buf_clk cell_2645 ( .C ( clk ), .D ( signal_17139 ), .Q ( signal_17338 ) ) ;
    buf_clk cell_2647 ( .C ( clk ), .D ( signal_17141 ), .Q ( signal_17340 ) ) ;
    buf_clk cell_2649 ( .C ( clk ), .D ( signal_17143 ), .Q ( signal_17342 ) ) ;
    buf_clk cell_2651 ( .C ( clk ), .D ( signal_17145 ), .Q ( signal_17344 ) ) ;
    buf_clk cell_2653 ( .C ( clk ), .D ( signal_17147 ), .Q ( signal_17346 ) ) ;
    buf_clk cell_2655 ( .C ( clk ), .D ( signal_960 ), .Q ( signal_17348 ) ) ;
    buf_clk cell_2657 ( .C ( clk ), .D ( signal_2496 ), .Q ( signal_17350 ) ) ;
    buf_clk cell_2659 ( .C ( clk ), .D ( signal_2497 ), .Q ( signal_17352 ) ) ;
    buf_clk cell_2661 ( .C ( clk ), .D ( signal_2498 ), .Q ( signal_17354 ) ) ;
    buf_clk cell_2663 ( .C ( clk ), .D ( signal_2499 ), .Q ( signal_17356 ) ) ;
    buf_clk cell_2665 ( .C ( clk ), .D ( signal_17199 ), .Q ( signal_17358 ) ) ;
    buf_clk cell_2667 ( .C ( clk ), .D ( signal_17201 ), .Q ( signal_17360 ) ) ;
    buf_clk cell_2669 ( .C ( clk ), .D ( signal_17203 ), .Q ( signal_17362 ) ) ;
    buf_clk cell_2671 ( .C ( clk ), .D ( signal_17205 ), .Q ( signal_17364 ) ) ;
    buf_clk cell_2673 ( .C ( clk ), .D ( signal_17207 ), .Q ( signal_17366 ) ) ;
    buf_clk cell_2675 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_17368 ) ) ;
    buf_clk cell_2677 ( .C ( clk ), .D ( signal_2456 ), .Q ( signal_17370 ) ) ;
    buf_clk cell_2679 ( .C ( clk ), .D ( signal_2457 ), .Q ( signal_17372 ) ) ;
    buf_clk cell_2681 ( .C ( clk ), .D ( signal_2458 ), .Q ( signal_17374 ) ) ;
    buf_clk cell_2683 ( .C ( clk ), .D ( signal_2459 ), .Q ( signal_17376 ) ) ;
    buf_clk cell_2685 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_17378 ) ) ;
    buf_clk cell_2687 ( .C ( clk ), .D ( signal_2656 ), .Q ( signal_17380 ) ) ;
    buf_clk cell_2689 ( .C ( clk ), .D ( signal_2657 ), .Q ( signal_17382 ) ) ;
    buf_clk cell_2691 ( .C ( clk ), .D ( signal_2658 ), .Q ( signal_17384 ) ) ;
    buf_clk cell_2693 ( .C ( clk ), .D ( signal_2659 ), .Q ( signal_17386 ) ) ;
    buf_clk cell_2695 ( .C ( clk ), .D ( signal_17089 ), .Q ( signal_17388 ) ) ;
    buf_clk cell_2697 ( .C ( clk ), .D ( signal_17091 ), .Q ( signal_17390 ) ) ;
    buf_clk cell_2699 ( .C ( clk ), .D ( signal_17093 ), .Q ( signal_17392 ) ) ;
    buf_clk cell_2701 ( .C ( clk ), .D ( signal_17095 ), .Q ( signal_17394 ) ) ;
    buf_clk cell_2703 ( .C ( clk ), .D ( signal_17097 ), .Q ( signal_17396 ) ) ;
    buf_clk cell_2705 ( .C ( clk ), .D ( signal_17129 ), .Q ( signal_17398 ) ) ;
    buf_clk cell_2707 ( .C ( clk ), .D ( signal_17131 ), .Q ( signal_17400 ) ) ;
    buf_clk cell_2709 ( .C ( clk ), .D ( signal_17133 ), .Q ( signal_17402 ) ) ;
    buf_clk cell_2711 ( .C ( clk ), .D ( signal_17135 ), .Q ( signal_17404 ) ) ;
    buf_clk cell_2713 ( .C ( clk ), .D ( signal_17137 ), .Q ( signal_17406 ) ) ;
    buf_clk cell_2715 ( .C ( clk ), .D ( signal_989 ), .Q ( signal_17408 ) ) ;
    buf_clk cell_2717 ( .C ( clk ), .D ( signal_2612 ), .Q ( signal_17410 ) ) ;
    buf_clk cell_2719 ( .C ( clk ), .D ( signal_2613 ), .Q ( signal_17412 ) ) ;
    buf_clk cell_2721 ( .C ( clk ), .D ( signal_2614 ), .Q ( signal_17414 ) ) ;
    buf_clk cell_2723 ( .C ( clk ), .D ( signal_2615 ), .Q ( signal_17416 ) ) ;
    buf_clk cell_2725 ( .C ( clk ), .D ( signal_17169 ), .Q ( signal_17418 ) ) ;
    buf_clk cell_2727 ( .C ( clk ), .D ( signal_17171 ), .Q ( signal_17420 ) ) ;
    buf_clk cell_2729 ( .C ( clk ), .D ( signal_17173 ), .Q ( signal_17422 ) ) ;
    buf_clk cell_2731 ( .C ( clk ), .D ( signal_17175 ), .Q ( signal_17424 ) ) ;
    buf_clk cell_2733 ( .C ( clk ), .D ( signal_17177 ), .Q ( signal_17426 ) ) ;
    buf_clk cell_2735 ( .C ( clk ), .D ( signal_986 ), .Q ( signal_17428 ) ) ;
    buf_clk cell_2737 ( .C ( clk ), .D ( signal_2600 ), .Q ( signal_17430 ) ) ;
    buf_clk cell_2739 ( .C ( clk ), .D ( signal_2601 ), .Q ( signal_17432 ) ) ;
    buf_clk cell_2741 ( .C ( clk ), .D ( signal_2602 ), .Q ( signal_17434 ) ) ;
    buf_clk cell_2743 ( .C ( clk ), .D ( signal_2603 ), .Q ( signal_17436 ) ) ;
    buf_clk cell_2745 ( .C ( clk ), .D ( signal_1032 ), .Q ( signal_17438 ) ) ;
    buf_clk cell_2747 ( .C ( clk ), .D ( signal_2784 ), .Q ( signal_17440 ) ) ;
    buf_clk cell_2749 ( .C ( clk ), .D ( signal_2785 ), .Q ( signal_17442 ) ) ;
    buf_clk cell_2751 ( .C ( clk ), .D ( signal_2786 ), .Q ( signal_17444 ) ) ;
    buf_clk cell_2753 ( .C ( clk ), .D ( signal_2787 ), .Q ( signal_17446 ) ) ;
    buf_clk cell_2755 ( .C ( clk ), .D ( signal_1016 ), .Q ( signal_17448 ) ) ;
    buf_clk cell_2757 ( .C ( clk ), .D ( signal_2720 ), .Q ( signal_17450 ) ) ;
    buf_clk cell_2759 ( .C ( clk ), .D ( signal_2721 ), .Q ( signal_17452 ) ) ;
    buf_clk cell_2761 ( .C ( clk ), .D ( signal_2722 ), .Q ( signal_17454 ) ) ;
    buf_clk cell_2763 ( .C ( clk ), .D ( signal_2723 ), .Q ( signal_17456 ) ) ;
    buf_clk cell_2765 ( .C ( clk ), .D ( signal_17149 ), .Q ( signal_17458 ) ) ;
    buf_clk cell_2767 ( .C ( clk ), .D ( signal_17151 ), .Q ( signal_17460 ) ) ;
    buf_clk cell_2769 ( .C ( clk ), .D ( signal_17153 ), .Q ( signal_17462 ) ) ;
    buf_clk cell_2771 ( .C ( clk ), .D ( signal_17155 ), .Q ( signal_17464 ) ) ;
    buf_clk cell_2773 ( .C ( clk ), .D ( signal_17157 ), .Q ( signal_17466 ) ) ;
    buf_clk cell_2775 ( .C ( clk ), .D ( signal_17179 ), .Q ( signal_17468 ) ) ;
    buf_clk cell_2777 ( .C ( clk ), .D ( signal_17181 ), .Q ( signal_17470 ) ) ;
    buf_clk cell_2779 ( .C ( clk ), .D ( signal_17183 ), .Q ( signal_17472 ) ) ;
    buf_clk cell_2781 ( .C ( clk ), .D ( signal_17185 ), .Q ( signal_17474 ) ) ;
    buf_clk cell_2783 ( .C ( clk ), .D ( signal_17187 ), .Q ( signal_17476 ) ) ;
    buf_clk cell_2785 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_17478 ) ) ;
    buf_clk cell_2787 ( .C ( clk ), .D ( signal_2504 ), .Q ( signal_17480 ) ) ;
    buf_clk cell_2789 ( .C ( clk ), .D ( signal_2505 ), .Q ( signal_17482 ) ) ;
    buf_clk cell_2791 ( .C ( clk ), .D ( signal_2506 ), .Q ( signal_17484 ) ) ;
    buf_clk cell_2793 ( .C ( clk ), .D ( signal_2507 ), .Q ( signal_17486 ) ) ;
    buf_clk cell_2795 ( .C ( clk ), .D ( signal_998 ), .Q ( signal_17488 ) ) ;
    buf_clk cell_2797 ( .C ( clk ), .D ( signal_2648 ), .Q ( signal_17490 ) ) ;
    buf_clk cell_2799 ( .C ( clk ), .D ( signal_2649 ), .Q ( signal_17492 ) ) ;
    buf_clk cell_2801 ( .C ( clk ), .D ( signal_2650 ), .Q ( signal_17494 ) ) ;
    buf_clk cell_2803 ( .C ( clk ), .D ( signal_2651 ), .Q ( signal_17496 ) ) ;
    buf_clk cell_2805 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_17498 ) ) ;
    buf_clk cell_2807 ( .C ( clk ), .D ( signal_2660 ), .Q ( signal_17500 ) ) ;
    buf_clk cell_2809 ( .C ( clk ), .D ( signal_2661 ), .Q ( signal_17502 ) ) ;
    buf_clk cell_2811 ( .C ( clk ), .D ( signal_2662 ), .Q ( signal_17504 ) ) ;
    buf_clk cell_2813 ( .C ( clk ), .D ( signal_2663 ), .Q ( signal_17506 ) ) ;
    buf_clk cell_2815 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_17508 ) ) ;
    buf_clk cell_2817 ( .C ( clk ), .D ( signal_2692 ), .Q ( signal_17510 ) ) ;
    buf_clk cell_2819 ( .C ( clk ), .D ( signal_2693 ), .Q ( signal_17512 ) ) ;
    buf_clk cell_2821 ( .C ( clk ), .D ( signal_2694 ), .Q ( signal_17514 ) ) ;
    buf_clk cell_2823 ( .C ( clk ), .D ( signal_2695 ), .Q ( signal_17516 ) ) ;
    buf_clk cell_2825 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_17518 ) ) ;
    buf_clk cell_2827 ( .C ( clk ), .D ( signal_2468 ), .Q ( signal_17520 ) ) ;
    buf_clk cell_2829 ( .C ( clk ), .D ( signal_2469 ), .Q ( signal_17522 ) ) ;
    buf_clk cell_2831 ( .C ( clk ), .D ( signal_2470 ), .Q ( signal_17524 ) ) ;
    buf_clk cell_2833 ( .C ( clk ), .D ( signal_2471 ), .Q ( signal_17526 ) ) ;
    buf_clk cell_2835 ( .C ( clk ), .D ( signal_988 ), .Q ( signal_17528 ) ) ;
    buf_clk cell_2837 ( .C ( clk ), .D ( signal_2608 ), .Q ( signal_17530 ) ) ;
    buf_clk cell_2839 ( .C ( clk ), .D ( signal_2609 ), .Q ( signal_17532 ) ) ;
    buf_clk cell_2841 ( .C ( clk ), .D ( signal_2610 ), .Q ( signal_17534 ) ) ;
    buf_clk cell_2843 ( .C ( clk ), .D ( signal_2611 ), .Q ( signal_17536 ) ) ;
    buf_clk cell_2845 ( .C ( clk ), .D ( signal_17099 ), .Q ( signal_17538 ) ) ;
    buf_clk cell_2847 ( .C ( clk ), .D ( signal_17101 ), .Q ( signal_17540 ) ) ;
    buf_clk cell_2849 ( .C ( clk ), .D ( signal_17103 ), .Q ( signal_17542 ) ) ;
    buf_clk cell_2851 ( .C ( clk ), .D ( signal_17105 ), .Q ( signal_17544 ) ) ;
    buf_clk cell_2853 ( .C ( clk ), .D ( signal_17107 ), .Q ( signal_17546 ) ) ;
    buf_clk cell_2855 ( .C ( clk ), .D ( signal_1004 ), .Q ( signal_17548 ) ) ;
    buf_clk cell_2857 ( .C ( clk ), .D ( signal_2672 ), .Q ( signal_17550 ) ) ;
    buf_clk cell_2859 ( .C ( clk ), .D ( signal_2673 ), .Q ( signal_17552 ) ) ;
    buf_clk cell_2861 ( .C ( clk ), .D ( signal_2674 ), .Q ( signal_17554 ) ) ;
    buf_clk cell_2863 ( .C ( clk ), .D ( signal_2675 ), .Q ( signal_17556 ) ) ;
    buf_clk cell_2865 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_17558 ) ) ;
    buf_clk cell_2867 ( .C ( clk ), .D ( signal_2484 ), .Q ( signal_17560 ) ) ;
    buf_clk cell_2869 ( .C ( clk ), .D ( signal_2485 ), .Q ( signal_17562 ) ) ;
    buf_clk cell_2871 ( .C ( clk ), .D ( signal_2486 ), .Q ( signal_17564 ) ) ;
    buf_clk cell_2873 ( .C ( clk ), .D ( signal_2487 ), .Q ( signal_17566 ) ) ;
    buf_clk cell_2877 ( .C ( clk ), .D ( signal_17569 ), .Q ( signal_17570 ) ) ;
    buf_clk cell_2881 ( .C ( clk ), .D ( signal_17573 ), .Q ( signal_17574 ) ) ;
    buf_clk cell_2885 ( .C ( clk ), .D ( signal_17577 ), .Q ( signal_17578 ) ) ;
    buf_clk cell_2889 ( .C ( clk ), .D ( signal_17581 ), .Q ( signal_17582 ) ) ;
    buf_clk cell_2893 ( .C ( clk ), .D ( signal_17585 ), .Q ( signal_17586 ) ) ;
    buf_clk cell_2895 ( .C ( clk ), .D ( signal_984 ), .Q ( signal_17588 ) ) ;
    buf_clk cell_2897 ( .C ( clk ), .D ( signal_2592 ), .Q ( signal_17590 ) ) ;
    buf_clk cell_2899 ( .C ( clk ), .D ( signal_2593 ), .Q ( signal_17592 ) ) ;
    buf_clk cell_2901 ( .C ( clk ), .D ( signal_2594 ), .Q ( signal_17594 ) ) ;
    buf_clk cell_2903 ( .C ( clk ), .D ( signal_2595 ), .Q ( signal_17596 ) ) ;
    buf_clk cell_2905 ( .C ( clk ), .D ( signal_997 ), .Q ( signal_17598 ) ) ;
    buf_clk cell_2907 ( .C ( clk ), .D ( signal_2644 ), .Q ( signal_17600 ) ) ;
    buf_clk cell_2909 ( .C ( clk ), .D ( signal_2645 ), .Q ( signal_17602 ) ) ;
    buf_clk cell_2911 ( .C ( clk ), .D ( signal_2646 ), .Q ( signal_17604 ) ) ;
    buf_clk cell_2913 ( .C ( clk ), .D ( signal_2647 ), .Q ( signal_17606 ) ) ;
    buf_clk cell_2915 ( .C ( clk ), .D ( signal_1007 ), .Q ( signal_17608 ) ) ;
    buf_clk cell_2917 ( .C ( clk ), .D ( signal_2684 ), .Q ( signal_17610 ) ) ;
    buf_clk cell_2919 ( .C ( clk ), .D ( signal_2685 ), .Q ( signal_17612 ) ) ;
    buf_clk cell_2921 ( .C ( clk ), .D ( signal_2686 ), .Q ( signal_17614 ) ) ;
    buf_clk cell_2923 ( .C ( clk ), .D ( signal_2687 ), .Q ( signal_17616 ) ) ;
    buf_clk cell_2925 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_17618 ) ) ;
    buf_clk cell_2927 ( .C ( clk ), .D ( signal_2460 ), .Q ( signal_17620 ) ) ;
    buf_clk cell_2929 ( .C ( clk ), .D ( signal_2461 ), .Q ( signal_17622 ) ) ;
    buf_clk cell_2931 ( .C ( clk ), .D ( signal_2462 ), .Q ( signal_17624 ) ) ;
    buf_clk cell_2933 ( .C ( clk ), .D ( signal_2463 ), .Q ( signal_17626 ) ) ;
    buf_clk cell_2935 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_17628 ) ) ;
    buf_clk cell_2937 ( .C ( clk ), .D ( signal_2580 ), .Q ( signal_17630 ) ) ;
    buf_clk cell_2939 ( .C ( clk ), .D ( signal_2581 ), .Q ( signal_17632 ) ) ;
    buf_clk cell_2941 ( .C ( clk ), .D ( signal_2582 ), .Q ( signal_17634 ) ) ;
    buf_clk cell_2943 ( .C ( clk ), .D ( signal_2583 ), .Q ( signal_17636 ) ) ;
    buf_clk cell_2945 ( .C ( clk ), .D ( signal_17079 ), .Q ( signal_17638 ) ) ;
    buf_clk cell_2947 ( .C ( clk ), .D ( signal_17081 ), .Q ( signal_17640 ) ) ;
    buf_clk cell_2949 ( .C ( clk ), .D ( signal_17083 ), .Q ( signal_17642 ) ) ;
    buf_clk cell_2951 ( .C ( clk ), .D ( signal_17085 ), .Q ( signal_17644 ) ) ;
    buf_clk cell_2953 ( .C ( clk ), .D ( signal_17087 ), .Q ( signal_17646 ) ) ;
    buf_clk cell_2955 ( .C ( clk ), .D ( signal_990 ), .Q ( signal_17648 ) ) ;
    buf_clk cell_2957 ( .C ( clk ), .D ( signal_2616 ), .Q ( signal_17650 ) ) ;
    buf_clk cell_2959 ( .C ( clk ), .D ( signal_2617 ), .Q ( signal_17652 ) ) ;
    buf_clk cell_2961 ( .C ( clk ), .D ( signal_2618 ), .Q ( signal_17654 ) ) ;
    buf_clk cell_2963 ( .C ( clk ), .D ( signal_2619 ), .Q ( signal_17656 ) ) ;
    buf_clk cell_2965 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_17658 ) ) ;
    buf_clk cell_2967 ( .C ( clk ), .D ( signal_2680 ), .Q ( signal_17660 ) ) ;
    buf_clk cell_2969 ( .C ( clk ), .D ( signal_2681 ), .Q ( signal_17662 ) ) ;
    buf_clk cell_2971 ( .C ( clk ), .D ( signal_2682 ), .Q ( signal_17664 ) ) ;
    buf_clk cell_2973 ( .C ( clk ), .D ( signal_2683 ), .Q ( signal_17666 ) ) ;
    buf_clk cell_2975 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_17668 ) ) ;
    buf_clk cell_2977 ( .C ( clk ), .D ( signal_2588 ), .Q ( signal_17670 ) ) ;
    buf_clk cell_2979 ( .C ( clk ), .D ( signal_2589 ), .Q ( signal_17672 ) ) ;
    buf_clk cell_2981 ( .C ( clk ), .D ( signal_2590 ), .Q ( signal_17674 ) ) ;
    buf_clk cell_2983 ( .C ( clk ), .D ( signal_2591 ), .Q ( signal_17676 ) ) ;
    buf_clk cell_2985 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_17678 ) ) ;
    buf_clk cell_2987 ( .C ( clk ), .D ( signal_2576 ), .Q ( signal_17680 ) ) ;
    buf_clk cell_2989 ( .C ( clk ), .D ( signal_2577 ), .Q ( signal_17682 ) ) ;
    buf_clk cell_2991 ( .C ( clk ), .D ( signal_2578 ), .Q ( signal_17684 ) ) ;
    buf_clk cell_2993 ( .C ( clk ), .D ( signal_2579 ), .Q ( signal_17686 ) ) ;
    buf_clk cell_2995 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_17688 ) ) ;
    buf_clk cell_2997 ( .C ( clk ), .D ( signal_2652 ), .Q ( signal_17690 ) ) ;
    buf_clk cell_2999 ( .C ( clk ), .D ( signal_2653 ), .Q ( signal_17692 ) ) ;
    buf_clk cell_3001 ( .C ( clk ), .D ( signal_2654 ), .Q ( signal_17694 ) ) ;
    buf_clk cell_3003 ( .C ( clk ), .D ( signal_2655 ), .Q ( signal_17696 ) ) ;
    buf_clk cell_3005 ( .C ( clk ), .D ( signal_972 ), .Q ( signal_17698 ) ) ;
    buf_clk cell_3007 ( .C ( clk ), .D ( signal_2544 ), .Q ( signal_17700 ) ) ;
    buf_clk cell_3009 ( .C ( clk ), .D ( signal_2545 ), .Q ( signal_17702 ) ) ;
    buf_clk cell_3011 ( .C ( clk ), .D ( signal_2546 ), .Q ( signal_17704 ) ) ;
    buf_clk cell_3013 ( .C ( clk ), .D ( signal_2547 ), .Q ( signal_17706 ) ) ;
    buf_clk cell_3015 ( .C ( clk ), .D ( signal_976 ), .Q ( signal_17708 ) ) ;
    buf_clk cell_3017 ( .C ( clk ), .D ( signal_2560 ), .Q ( signal_17710 ) ) ;
    buf_clk cell_3019 ( .C ( clk ), .D ( signal_2561 ), .Q ( signal_17712 ) ) ;
    buf_clk cell_3021 ( .C ( clk ), .D ( signal_2562 ), .Q ( signal_17714 ) ) ;
    buf_clk cell_3023 ( .C ( clk ), .D ( signal_2563 ), .Q ( signal_17716 ) ) ;
    buf_clk cell_3025 ( .C ( clk ), .D ( signal_1057 ), .Q ( signal_17718 ) ) ;
    buf_clk cell_3027 ( .C ( clk ), .D ( signal_2884 ), .Q ( signal_17720 ) ) ;
    buf_clk cell_3029 ( .C ( clk ), .D ( signal_2885 ), .Q ( signal_17722 ) ) ;
    buf_clk cell_3031 ( .C ( clk ), .D ( signal_2886 ), .Q ( signal_17724 ) ) ;
    buf_clk cell_3033 ( .C ( clk ), .D ( signal_2887 ), .Q ( signal_17726 ) ) ;
    buf_clk cell_3035 ( .C ( clk ), .D ( signal_1039 ), .Q ( signal_17728 ) ) ;
    buf_clk cell_3037 ( .C ( clk ), .D ( signal_2812 ), .Q ( signal_17730 ) ) ;
    buf_clk cell_3039 ( .C ( clk ), .D ( signal_2813 ), .Q ( signal_17732 ) ) ;
    buf_clk cell_3041 ( .C ( clk ), .D ( signal_2814 ), .Q ( signal_17734 ) ) ;
    buf_clk cell_3043 ( .C ( clk ), .D ( signal_2815 ), .Q ( signal_17736 ) ) ;
    buf_clk cell_3045 ( .C ( clk ), .D ( signal_1046 ), .Q ( signal_17738 ) ) ;
    buf_clk cell_3047 ( .C ( clk ), .D ( signal_2840 ), .Q ( signal_17740 ) ) ;
    buf_clk cell_3049 ( .C ( clk ), .D ( signal_2841 ), .Q ( signal_17742 ) ) ;
    buf_clk cell_3051 ( .C ( clk ), .D ( signal_2842 ), .Q ( signal_17744 ) ) ;
    buf_clk cell_3053 ( .C ( clk ), .D ( signal_2843 ), .Q ( signal_17746 ) ) ;
    buf_clk cell_3055 ( .C ( clk ), .D ( signal_1005 ), .Q ( signal_17748 ) ) ;
    buf_clk cell_3057 ( .C ( clk ), .D ( signal_2676 ), .Q ( signal_17750 ) ) ;
    buf_clk cell_3059 ( .C ( clk ), .D ( signal_2677 ), .Q ( signal_17752 ) ) ;
    buf_clk cell_3061 ( .C ( clk ), .D ( signal_2678 ), .Q ( signal_17754 ) ) ;
    buf_clk cell_3063 ( .C ( clk ), .D ( signal_2679 ), .Q ( signal_17756 ) ) ;
    buf_clk cell_3065 ( .C ( clk ), .D ( signal_1041 ), .Q ( signal_17758 ) ) ;
    buf_clk cell_3067 ( .C ( clk ), .D ( signal_2820 ), .Q ( signal_17760 ) ) ;
    buf_clk cell_3069 ( .C ( clk ), .D ( signal_2821 ), .Q ( signal_17762 ) ) ;
    buf_clk cell_3071 ( .C ( clk ), .D ( signal_2822 ), .Q ( signal_17764 ) ) ;
    buf_clk cell_3073 ( .C ( clk ), .D ( signal_2823 ), .Q ( signal_17766 ) ) ;
    buf_clk cell_3075 ( .C ( clk ), .D ( signal_1034 ), .Q ( signal_17768 ) ) ;
    buf_clk cell_3077 ( .C ( clk ), .D ( signal_2792 ), .Q ( signal_17770 ) ) ;
    buf_clk cell_3079 ( .C ( clk ), .D ( signal_2793 ), .Q ( signal_17772 ) ) ;
    buf_clk cell_3081 ( .C ( clk ), .D ( signal_2794 ), .Q ( signal_17774 ) ) ;
    buf_clk cell_3083 ( .C ( clk ), .D ( signal_2795 ), .Q ( signal_17776 ) ) ;
    buf_clk cell_3085 ( .C ( clk ), .D ( signal_996 ), .Q ( signal_17778 ) ) ;
    buf_clk cell_3087 ( .C ( clk ), .D ( signal_2640 ), .Q ( signal_17780 ) ) ;
    buf_clk cell_3089 ( .C ( clk ), .D ( signal_2641 ), .Q ( signal_17782 ) ) ;
    buf_clk cell_3091 ( .C ( clk ), .D ( signal_2642 ), .Q ( signal_17784 ) ) ;
    buf_clk cell_3093 ( .C ( clk ), .D ( signal_2643 ), .Q ( signal_17786 ) ) ;
    buf_clk cell_3095 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_17788 ) ) ;
    buf_clk cell_3097 ( .C ( clk ), .D ( signal_2632 ), .Q ( signal_17790 ) ) ;
    buf_clk cell_3099 ( .C ( clk ), .D ( signal_2633 ), .Q ( signal_17792 ) ) ;
    buf_clk cell_3101 ( .C ( clk ), .D ( signal_2634 ), .Q ( signal_17794 ) ) ;
    buf_clk cell_3103 ( .C ( clk ), .D ( signal_2635 ), .Q ( signal_17796 ) ) ;
    buf_clk cell_3105 ( .C ( clk ), .D ( signal_985 ), .Q ( signal_17798 ) ) ;
    buf_clk cell_3107 ( .C ( clk ), .D ( signal_2596 ), .Q ( signal_17800 ) ) ;
    buf_clk cell_3109 ( .C ( clk ), .D ( signal_2597 ), .Q ( signal_17802 ) ) ;
    buf_clk cell_3111 ( .C ( clk ), .D ( signal_2598 ), .Q ( signal_17804 ) ) ;
    buf_clk cell_3113 ( .C ( clk ), .D ( signal_2599 ), .Q ( signal_17806 ) ) ;
    buf_clk cell_3227 ( .C ( clk ), .D ( signal_17919 ), .Q ( signal_17920 ) ) ;
    buf_clk cell_3233 ( .C ( clk ), .D ( signal_17925 ), .Q ( signal_17926 ) ) ;
    buf_clk cell_3239 ( .C ( clk ), .D ( signal_17931 ), .Q ( signal_17932 ) ) ;
    buf_clk cell_3245 ( .C ( clk ), .D ( signal_17937 ), .Q ( signal_17938 ) ) ;
    buf_clk cell_3251 ( .C ( clk ), .D ( signal_17943 ), .Q ( signal_17944 ) ) ;
    buf_clk cell_3455 ( .C ( clk ), .D ( signal_1054 ), .Q ( signal_18148 ) ) ;
    buf_clk cell_3459 ( .C ( clk ), .D ( signal_2872 ), .Q ( signal_18152 ) ) ;
    buf_clk cell_3463 ( .C ( clk ), .D ( signal_2873 ), .Q ( signal_18156 ) ) ;
    buf_clk cell_3467 ( .C ( clk ), .D ( signal_2874 ), .Q ( signal_18160 ) ) ;
    buf_clk cell_3471 ( .C ( clk ), .D ( signal_2875 ), .Q ( signal_18164 ) ) ;
    buf_clk cell_3495 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_18188 ) ) ;
    buf_clk cell_3499 ( .C ( clk ), .D ( signal_2464 ), .Q ( signal_18192 ) ) ;
    buf_clk cell_3503 ( .C ( clk ), .D ( signal_2465 ), .Q ( signal_18196 ) ) ;
    buf_clk cell_3507 ( .C ( clk ), .D ( signal_2466 ), .Q ( signal_18200 ) ) ;
    buf_clk cell_3511 ( .C ( clk ), .D ( signal_2467 ), .Q ( signal_18204 ) ) ;
    buf_clk cell_3625 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_18318 ) ) ;
    buf_clk cell_3629 ( .C ( clk ), .D ( signal_2488 ), .Q ( signal_18322 ) ) ;
    buf_clk cell_3633 ( .C ( clk ), .D ( signal_2489 ), .Q ( signal_18326 ) ) ;
    buf_clk cell_3637 ( .C ( clk ), .D ( signal_2490 ), .Q ( signal_18330 ) ) ;
    buf_clk cell_3641 ( .C ( clk ), .D ( signal_2491 ), .Q ( signal_18334 ) ) ;
    buf_clk cell_3655 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_18348 ) ) ;
    buf_clk cell_3659 ( .C ( clk ), .D ( signal_2472 ), .Q ( signal_18352 ) ) ;
    buf_clk cell_3663 ( .C ( clk ), .D ( signal_2473 ), .Q ( signal_18356 ) ) ;
    buf_clk cell_3667 ( .C ( clk ), .D ( signal_2474 ), .Q ( signal_18360 ) ) ;
    buf_clk cell_3671 ( .C ( clk ), .D ( signal_2475 ), .Q ( signal_18364 ) ) ;
    buf_clk cell_3707 ( .C ( clk ), .D ( signal_18399 ), .Q ( signal_18400 ) ) ;
    buf_clk cell_3713 ( .C ( clk ), .D ( signal_18405 ), .Q ( signal_18406 ) ) ;
    buf_clk cell_3719 ( .C ( clk ), .D ( signal_18411 ), .Q ( signal_18412 ) ) ;
    buf_clk cell_3725 ( .C ( clk ), .D ( signal_18417 ), .Q ( signal_18418 ) ) ;
    buf_clk cell_3731 ( .C ( clk ), .D ( signal_18423 ), .Q ( signal_18424 ) ) ;
    buf_clk cell_3775 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_18468 ) ) ;
    buf_clk cell_3779 ( .C ( clk ), .D ( signal_2508 ), .Q ( signal_18472 ) ) ;
    buf_clk cell_3783 ( .C ( clk ), .D ( signal_2509 ), .Q ( signal_18476 ) ) ;
    buf_clk cell_3787 ( .C ( clk ), .D ( signal_2510 ), .Q ( signal_18480 ) ) ;
    buf_clk cell_3791 ( .C ( clk ), .D ( signal_2511 ), .Q ( signal_18484 ) ) ;
    buf_clk cell_3885 ( .C ( clk ), .D ( signal_17119 ), .Q ( signal_18578 ) ) ;
    buf_clk cell_3889 ( .C ( clk ), .D ( signal_17121 ), .Q ( signal_18582 ) ) ;
    buf_clk cell_3893 ( .C ( clk ), .D ( signal_17123 ), .Q ( signal_18586 ) ) ;
    buf_clk cell_3897 ( .C ( clk ), .D ( signal_17125 ), .Q ( signal_18590 ) ) ;
    buf_clk cell_3901 ( .C ( clk ), .D ( signal_17127 ), .Q ( signal_18594 ) ) ;
    buf_clk cell_4077 ( .C ( clk ), .D ( signal_18769 ), .Q ( signal_18770 ) ) ;
    buf_clk cell_4085 ( .C ( clk ), .D ( signal_18777 ), .Q ( signal_18778 ) ) ;
    buf_clk cell_4093 ( .C ( clk ), .D ( signal_18785 ), .Q ( signal_18786 ) ) ;
    buf_clk cell_4101 ( .C ( clk ), .D ( signal_18793 ), .Q ( signal_18794 ) ) ;
    buf_clk cell_4109 ( .C ( clk ), .D ( signal_18801 ), .Q ( signal_18802 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_988 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .clk ( clk ), .r ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .c ({signal_2671, signal_2670, signal_2669, signal_2668, signal_1003}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_999 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2479, signal_2478, signal_2477, signal_2476, signal_955}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .c ({signal_2715, signal_2714, signal_2713, signal_2712, signal_1014}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1004 ( .a ({signal_17087, signal_17085, signal_17083, signal_17081, signal_17079}), .b ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .clk ( clk ), .r ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_2735, signal_2734, signal_2733, signal_2732, signal_1019}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1005 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2491, signal_2490, signal_2489, signal_2488, signal_958}), .clk ( clk ), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .c ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1020}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1006 ( .a ({signal_17097, signal_17095, signal_17093, signal_17091, signal_17089}), .b ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .c ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1007 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}), .clk ( clk ), .r ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_2747, signal_2746, signal_2745, signal_2744, signal_1022}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1008 ( .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .b ({signal_2495, signal_2494, signal_2493, signal_2492, signal_959}), .clk ( clk ), .r ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .c ({signal_2751, signal_2750, signal_2749, signal_2748, signal_1023}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1009 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .c ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1024}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1010 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_2759, signal_2758, signal_2757, signal_2756, signal_1025}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1011 ( .a ({signal_2479, signal_2478, signal_2477, signal_2476, signal_955}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .c ({signal_2763, signal_2762, signal_2761, signal_2760, signal_1026}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1012 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .c ({signal_2767, signal_2766, signal_2765, signal_2764, signal_1027}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1013 ( .a ({signal_2459, signal_2458, signal_2457, signal_2456, signal_950}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_2771, signal_2770, signal_2769, signal_2768, signal_1028}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1014 ( .a ({signal_17117, signal_17115, signal_17113, signal_17111, signal_17109}), .b ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}), .clk ( clk ), .r ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .c ({signal_2775, signal_2774, signal_2773, signal_2772, signal_1029}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1015 ( .a ({signal_2483, signal_2482, signal_2481, signal_2480, signal_956}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .c ({signal_2779, signal_2778, signal_2777, signal_2776, signal_1030}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1033 ( .a ({signal_2671, signal_2670, signal_2669, signal_2668, signal_1003}), .b ({signal_2851, signal_2850, signal_2849, signal_2848, signal_1048}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1040 ( .a ({signal_2715, signal_2714, signal_2713, signal_2712, signal_1014}), .b ({signal_2879, signal_2878, signal_2877, signal_2876, signal_1055}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1044 ( .a ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1020}), .b ({signal_2895, signal_2894, signal_2893, signal_2892, signal_1059}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1045 ( .a ({signal_2751, signal_2750, signal_2749, signal_2748, signal_1023}), .b ({signal_2899, signal_2898, signal_2897, signal_2896, signal_1060}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1046 ( .a ({signal_2759, signal_2758, signal_2757, signal_2756, signal_1025}), .b ({signal_2903, signal_2902, signal_2901, signal_2900, signal_1061}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1047 ( .a ({signal_2763, signal_2762, signal_2761, signal_2760, signal_1026}), .b ({signal_2907, signal_2906, signal_2905, signal_2904, signal_1062}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1048 ( .a ({signal_2767, signal_2766, signal_2765, signal_2764, signal_1027}), .b ({signal_2911, signal_2910, signal_2909, signal_2908, signal_1063}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1049 ( .a ({signal_2771, signal_2770, signal_2769, signal_2768, signal_1028}), .b ({signal_2915, signal_2914, signal_2913, signal_2912, signal_1064}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1050 ( .a ({signal_2775, signal_2774, signal_2773, signal_2772, signal_1029}), .b ({signal_2919, signal_2918, signal_2917, signal_2916, signal_1065}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1051 ( .a ({signal_2779, signal_2778, signal_2777, signal_2776, signal_1030}), .b ({signal_2923, signal_2922, signal_2921, signal_2920, signal_1066}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1052 ( .a ({signal_17097, signal_17095, signal_17093, signal_17091, signal_17089}), .b ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .clk ( clk ), .r ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_2927, signal_2926, signal_2925, signal_2924, signal_1067}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1053 ( .a ({signal_17127, signal_17125, signal_17123, signal_17121, signal_17119}), .b ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .clk ( clk ), .r ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .c ({signal_2931, signal_2930, signal_2929, signal_2928, signal_1068}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1054 ( .a ({signal_2527, signal_2526, signal_2525, signal_2524, signal_967}), .b ({signal_2531, signal_2530, signal_2529, signal_2528, signal_968}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .c ({signal_2935, signal_2934, signal_2933, signal_2932, signal_1069}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1055 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2523, signal_2522, signal_2521, signal_2520, signal_966}), .clk ( clk ), .r ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_2939, signal_2938, signal_2937, signal_2936, signal_1070}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1056 ( .a ({signal_17137, signal_17135, signal_17133, signal_17131, signal_17129}), .b ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .clk ( clk ), .r ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .c ({signal_2943, signal_2942, signal_2941, signal_2940, signal_1071}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1057 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .c ({signal_2947, signal_2946, signal_2945, signal_2944, signal_1072}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1058 ( .a ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .b ({signal_2491, signal_2490, signal_2489, signal_2488, signal_958}), .clk ( clk ), .r ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1059 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .clk ( clk ), .r ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .c ({signal_2955, signal_2954, signal_2953, signal_2952, signal_1074}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1060 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .c ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1061 ( .a ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .b ({signal_2655, signal_2654, signal_2653, signal_2652, signal_999}), .clk ( clk ), .r ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_2963, signal_2962, signal_2961, signal_2960, signal_1076}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1062 ( .a ({signal_17127, signal_17125, signal_17123, signal_17121, signal_17119}), .b ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .clk ( clk ), .r ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .c ({signal_2967, signal_2966, signal_2965, signal_2964, signal_1077}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1063 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .c ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1078}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1064 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2667, signal_2666, signal_2665, signal_2664, signal_1002}), .clk ( clk ), .r ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_2975, signal_2974, signal_2973, signal_2972, signal_1079}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1065 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .c ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1080}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1066 ( .a ({signal_17147, signal_17145, signal_17143, signal_17141, signal_17139}), .b ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .c ({signal_2983, signal_2982, signal_2981, signal_2980, signal_1081}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1067 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .clk ( clk ), .r ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1068 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .c ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1069 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .c ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1070 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}), .clk ( clk ), .r ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_2999, signal_2998, signal_2997, signal_2996, signal_1085}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1071 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .c ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1072 ( .a ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .c ({signal_3007, signal_3006, signal_3005, signal_3004, signal_1087}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1073 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .clk ( clk ), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_3011, signal_3010, signal_3009, signal_3008, signal_1088}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1074 ( .a ({signal_17087, signal_17085, signal_17083, signal_17081, signal_17079}), .b ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .clk ( clk ), .r ({Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .c ({signal_3015, signal_3014, signal_3013, signal_3012, signal_1089}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1075 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890]}), .c ({signal_3019, signal_3018, signal_3017, signal_3016, signal_1090}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1076 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_3023, signal_3022, signal_3021, signal_3020, signal_1091}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1077 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910]}), .c ({signal_3027, signal_3026, signal_3025, signal_3024, signal_1092}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1078 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .c ({signal_3031, signal_3030, signal_3029, signal_3028, signal_1093}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1079 ( .a ({signal_2459, signal_2458, signal_2457, signal_2456, signal_950}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .clk ( clk ), .r ({Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_3035, signal_3034, signal_3033, signal_3032, signal_1094}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1080 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2491, signal_2490, signal_2489, signal_2488, signal_958}), .clk ( clk ), .r ({Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .c ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1081 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1012}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950]}), .c ({signal_3043, signal_3042, signal_3041, signal_3040, signal_1096}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1082 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_3047, signal_3046, signal_3045, signal_3044, signal_1097}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1083 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .clk ( clk ), .r ({Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970]}), .c ({signal_3051, signal_3050, signal_3049, signal_3048, signal_1098}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1084 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .c ({signal_3055, signal_3054, signal_3053, signal_3052, signal_1099}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1086 ( .a ({signal_2587, signal_2586, signal_2585, signal_2584, signal_982}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_3063, signal_3062, signal_3061, signal_3060, signal_1101}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1087 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2587, signal_2586, signal_2585, signal_2584, signal_982}), .clk ( clk ), .r ({Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .c ({signal_3067, signal_3066, signal_3065, signal_3064, signal_1102}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1088 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010]}), .c ({signal_3071, signal_3070, signal_3069, signal_3068, signal_1103}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1089 ( .a ({signal_17097, signal_17095, signal_17093, signal_17091, signal_17089}), .b ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .clk ( clk ), .r ({Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_3075, signal_3074, signal_3073, signal_3072, signal_1104}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1090 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}), .clk ( clk ), .r ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030]}), .c ({signal_3079, signal_3078, signal_3077, signal_3076, signal_1105}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1091 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1016}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .c ({signal_3083, signal_3082, signal_3081, signal_3080, signal_1106}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1092 ( .a ({signal_17127, signal_17125, signal_17123, signal_17121, signal_17119}), .b ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .clk ( clk ), .r ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_3087, signal_3086, signal_3085, signal_3084, signal_1107}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1093 ( .a ({signal_17157, signal_17155, signal_17153, signal_17151, signal_17149}), .b ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .clk ( clk ), .r ({Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .c ({signal_3091, signal_3090, signal_3089, signal_3088, signal_1108}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1094 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1012}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070]}), .c ({signal_3095, signal_3094, signal_3093, signal_3092, signal_1109}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1095 ( .a ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_3099, signal_3098, signal_3097, signal_3096, signal_1110}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1096 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .clk ( clk ), .r ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090]}), .c ({signal_3103, signal_3102, signal_3101, signal_3100, signal_1111}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1097 ( .a ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .b ({signal_2711, signal_2710, signal_2709, signal_2708, signal_1013}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .c ({signal_3107, signal_3106, signal_3105, signal_3104, signal_1112}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1098 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_3111, signal_3110, signal_3109, signal_3108, signal_1113}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1099 ( .a ({signal_17167, signal_17165, signal_17163, signal_17161, signal_17159}), .b ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1010}), .clk ( clk ), .r ({Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .c ({signal_3115, signal_3114, signal_3113, signal_3112, signal_1114}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1100 ( .a ({signal_17137, signal_17135, signal_17133, signal_17131, signal_17129}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130]}), .c ({signal_3119, signal_3118, signal_3117, signal_3116, signal_1115}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1101 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1010}), .clk ( clk ), .r ({Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_3123, signal_3122, signal_3121, signal_3120, signal_1116}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1102 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150]}), .c ({signal_3127, signal_3126, signal_3125, signal_3124, signal_1117}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1103 ( .a ({signal_17147, signal_17145, signal_17143, signal_17141, signal_17139}), .b ({signal_2667, signal_2666, signal_2665, signal_2664, signal_1002}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .c ({signal_3131, signal_3130, signal_3129, signal_3128, signal_1118}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1104 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .clk ( clk ), .r ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_3135, signal_3134, signal_3133, signal_3132, signal_1119}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1105 ( .a ({signal_17177, signal_17175, signal_17173, signal_17171, signal_17169}), .b ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .clk ( clk ), .r ({Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .c ({signal_3139, signal_3138, signal_3137, signal_3136, signal_1120}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1106 ( .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190]}), .c ({signal_3143, signal_3142, signal_3141, signal_3140, signal_1121}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1107 ( .a ({signal_2499, signal_2498, signal_2497, signal_2496, signal_960}), .b ({signal_2731, signal_2730, signal_2729, signal_2728, signal_1018}), .clk ( clk ), .r ({Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_3147, signal_3146, signal_3145, signal_3144, signal_1122}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1108 ( .a ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .b ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}), .clk ( clk ), .r ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210]}), .c ({signal_3151, signal_3150, signal_3149, signal_3148, signal_1123}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1109 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2655, signal_2654, signal_2653, signal_2652, signal_999}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .c ({signal_3155, signal_3154, signal_3153, signal_3152, signal_1124}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1110 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_3159, signal_3158, signal_3157, signal_3156, signal_1125}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1111 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}), .clk ( clk ), .r ({Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .c ({signal_3163, signal_3162, signal_3161, signal_3160, signal_1126}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1112 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2483, signal_2482, signal_2481, signal_2480, signal_956}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250]}), .c ({signal_3167, signal_3166, signal_3165, signal_3164, signal_1127}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1113 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_2511, signal_2510, signal_2509, signal_2508, signal_963}), .clk ( clk ), .r ({Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_3171, signal_3170, signal_3169, signal_3168, signal_1128}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1114 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1016}), .clk ( clk ), .r ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270]}), .c ({signal_3175, signal_3174, signal_3173, signal_3172, signal_1129}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1115 ( .a ({signal_2475, signal_2474, signal_2473, signal_2472, signal_954}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .c ({signal_3179, signal_3178, signal_3177, signal_3176, signal_1130}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1116 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_3183, signal_3182, signal_3181, signal_3180, signal_1131}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1117 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .clk ( clk ), .r ({Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .c ({signal_3187, signal_3186, signal_3185, signal_3184, signal_1132}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1118 ( .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .b ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310]}), .c ({signal_3191, signal_3190, signal_3189, signal_3188, signal_1133}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1119 ( .a ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .clk ( clk ), .r ({Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_3195, signal_3194, signal_3193, signal_3192, signal_1134}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1120 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .clk ( clk ), .r ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330]}), .c ({signal_3199, signal_3198, signal_3197, signal_3196, signal_1135}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1121 ( .a ({signal_2619, signal_2618, signal_2617, signal_2616, signal_990}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .c ({signal_3203, signal_3202, signal_3201, signal_3200, signal_1136}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1122 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}), .clk ( clk ), .r ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_3207, signal_3206, signal_3205, signal_3204, signal_1137}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1123 ( .a ({signal_17157, signal_17155, signal_17153, signal_17151, signal_17149}), .b ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .clk ( clk ), .r ({Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .c ({signal_3211, signal_3210, signal_3209, signal_3208, signal_1138}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1125 ( .a ({signal_2587, signal_2586, signal_2585, signal_2584, signal_982}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370]}), .c ({signal_3219, signal_3218, signal_3217, signal_3216, signal_1140}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1126 ( .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .b ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .clk ( clk ), .r ({Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_3223, signal_3222, signal_3221, signal_3220, signal_1141}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1127 ( .a ({signal_2491, signal_2490, signal_2489, signal_2488, signal_958}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390]}), .c ({signal_3227, signal_3226, signal_3225, signal_3224, signal_1142}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1128 ( .a ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .c ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1129 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .clk ( clk ), .r ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_3235, signal_3234, signal_3233, signal_3232, signal_1144}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1130 ( .a ({signal_17147, signal_17145, signal_17143, signal_17141, signal_17139}), .b ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .clk ( clk ), .r ({Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .c ({signal_3239, signal_3238, signal_3237, signal_3236, signal_1145}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1131 ( .a ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .b ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1006}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430]}), .c ({signal_3243, signal_3242, signal_3241, signal_3240, signal_1146}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1133 ( .a ({signal_2475, signal_2474, signal_2473, signal_2472, signal_954}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_3251, signal_3250, signal_3249, signal_3248, signal_1148}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1134 ( .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450]}), .c ({signal_3255, signal_3254, signal_3253, signal_3252, signal_1149}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1135 ( .a ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .c ({signal_3259, signal_3258, signal_3257, signal_3256, signal_1150}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1136 ( .a ({signal_17187, signal_17185, signal_17183, signal_17181, signal_17179}), .b ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}), .clk ( clk ), .r ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_3263, signal_3262, signal_3261, signal_3260, signal_1151}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1137 ( .a ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .b ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .clk ( clk ), .r ({Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .c ({signal_3267, signal_3266, signal_3265, signal_3264, signal_1152}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1138 ( .a ({signal_17097, signal_17095, signal_17093, signal_17091, signal_17089}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490]}), .c ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1139 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_3275, signal_3274, signal_3273, signal_3272, signal_1154}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1141 ( .a ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510]}), .c ({signal_3283, signal_3282, signal_3281, signal_3280, signal_1156}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1142 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .c ({signal_3287, signal_3286, signal_3285, signal_3284, signal_1157}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1143 ( .a ({signal_17107, signal_17105, signal_17103, signal_17101, signal_17099}), .b ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .clk ( clk ), .r ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1144 ( .a ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .b ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .clk ( clk ), .r ({Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .c ({signal_3295, signal_3294, signal_3293, signal_3292, signal_1159}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1145 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550]}), .c ({signal_3299, signal_3298, signal_3297, signal_3296, signal_1160}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1146 ( .a ({signal_2467, signal_2466, signal_2465, signal_2464, signal_952}), .b ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .clk ( clk ), .r ({Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_3303, signal_3302, signal_3301, signal_3300, signal_1161}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1147 ( .a ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .clk ( clk ), .r ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570]}), .c ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1148 ( .a ({signal_2523, signal_2522, signal_2521, signal_2520, signal_966}), .b ({signal_2551, signal_2550, signal_2549, signal_2548, signal_973}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .c ({signal_3311, signal_3310, signal_3309, signal_3308, signal_1163}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1149 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_3315, signal_3314, signal_3313, signal_3312, signal_1164}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1150 ( .a ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .b ({signal_2703, signal_2702, signal_2701, signal_2700, signal_1011}), .clk ( clk ), .r ({Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .c ({signal_3319, signal_3318, signal_3317, signal_3316, signal_1165}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1151 ( .a ({signal_2587, signal_2586, signal_2585, signal_2584, signal_982}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610]}), .c ({signal_3323, signal_3322, signal_3321, signal_3320, signal_1166}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1152 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .clk ( clk ), .r ({Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_3327, signal_3326, signal_3325, signal_3324, signal_1167}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1153 ( .a ({signal_17187, signal_17185, signal_17183, signal_17181, signal_17179}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_994}), .clk ( clk ), .r ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630]}), .c ({signal_3331, signal_3330, signal_3329, signal_3328, signal_1168}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1154 ( .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .b ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1010}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .c ({signal_3335, signal_3334, signal_3333, signal_3332, signal_1169}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1156 ( .a ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1006}), .b ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1010}), .clk ( clk ), .r ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_3343, signal_3342, signal_3341, signal_3340, signal_1171}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1157 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .clk ( clk ), .r ({Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .c ({signal_3347, signal_3346, signal_3345, signal_3344, signal_1172}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1158 ( .a ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670]}), .c ({signal_3351, signal_3350, signal_3349, signal_3348, signal_1173}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1159 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1008}), .clk ( clk ), .r ({Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_3355, signal_3354, signal_3353, signal_3352, signal_1174}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1160 ( .a ({signal_17157, signal_17155, signal_17153, signal_17151, signal_17149}), .b ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .clk ( clk ), .r ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690]}), .c ({signal_3359, signal_3358, signal_3357, signal_3356, signal_1175}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1161 ( .a ({signal_17137, signal_17135, signal_17133, signal_17131, signal_17129}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .c ({signal_3363, signal_3362, signal_3361, signal_3360, signal_1176}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1162 ( .a ({signal_17127, signal_17125, signal_17123, signal_17121, signal_17119}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_3367, signal_3366, signal_3365, signal_3364, signal_1177}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1163 ( .a ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}), .b ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1015}), .clk ( clk ), .r ({Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .c ({signal_3371, signal_3370, signal_3369, signal_3368, signal_1178}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1164 ( .a ({signal_2523, signal_2522, signal_2521, signal_2520, signal_966}), .b ({signal_2547, signal_2546, signal_2545, signal_2544, signal_972}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730]}), .c ({signal_3375, signal_3374, signal_3373, signal_3372, signal_1179}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1165 ( .a ({signal_2543, signal_2542, signal_2541, signal_2540, signal_971}), .b ({signal_2547, signal_2546, signal_2545, signal_2544, signal_972}), .clk ( clk ), .r ({Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_3379, signal_3378, signal_3377, signal_3376, signal_1180}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1166 ( .a ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .b ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1012}), .clk ( clk ), .r ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750]}), .c ({signal_3383, signal_3382, signal_3381, signal_3380, signal_1181}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1167 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .c ({signal_3387, signal_3386, signal_3385, signal_3384, signal_1182}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1168 ( .a ({signal_2479, signal_2478, signal_2477, signal_2476, signal_955}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_3391, signal_3390, signal_3389, signal_3388, signal_1183}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1169 ( .a ({signal_17117, signal_17115, signal_17113, signal_17111, signal_17109}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .c ({signal_3395, signal_3394, signal_3393, signal_3392, signal_1184}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1170 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1000}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790]}), .c ({signal_3399, signal_3398, signal_3397, signal_3396, signal_1185}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1171 ( .a ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .b ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1015}), .clk ( clk ), .r ({Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_3403, signal_3402, signal_3401, signal_3400, signal_1186}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1172 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}), .clk ( clk ), .r ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810]}), .c ({signal_3407, signal_3406, signal_3405, signal_3404, signal_1187}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1174 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .c ({signal_3415, signal_3414, signal_3413, signal_3412, signal_1189}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1175 ( .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_983}), .b ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .clk ( clk ), .r ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_3419, signal_3418, signal_3417, signal_3416, signal_1190}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1176 ( .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_951}), .b ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .clk ( clk ), .r ({Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .c ({signal_3423, signal_3422, signal_3421, signal_3420, signal_1191}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1177 ( .a ({signal_2643, signal_2642, signal_2641, signal_2640, signal_996}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850]}), .c ({signal_3427, signal_3426, signal_3425, signal_3424, signal_1192}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1178 ( .a ({signal_2535, signal_2534, signal_2533, signal_2532, signal_969}), .b ({signal_2563, signal_2562, signal_2561, signal_2560, signal_976}), .clk ( clk ), .r ({Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_3431, signal_3430, signal_3429, signal_3428, signal_1193}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1179 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .clk ( clk ), .r ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870]}), .c ({signal_3435, signal_3434, signal_3433, signal_3432, signal_1194}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1180 ( .a ({signal_2607, signal_2606, signal_2605, signal_2604, signal_987}), .b ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .c ({signal_3439, signal_3438, signal_3437, signal_3436, signal_1195}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1181 ( .a ({signal_2507, signal_2506, signal_2505, signal_2504, signal_962}), .b ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .clk ( clk ), .r ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_3443, signal_3442, signal_3441, signal_3440, signal_1196}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1182 ( .a ({signal_17147, signal_17145, signal_17143, signal_17141, signal_17139}), .b ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .clk ( clk ), .r ({Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .c ({signal_3447, signal_3446, signal_3445, signal_3444, signal_1197}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1183 ( .a ({signal_2579, signal_2578, signal_2577, signal_2576, signal_980}), .b ({signal_2503, signal_2502, signal_2501, signal_2500, signal_961}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910]}), .c ({signal_3451, signal_3450, signal_3449, signal_3448, signal_1198}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1185 ( .a ({signal_2595, signal_2594, signal_2593, signal_2592, signal_984}), .b ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1015}), .clk ( clk ), .r ({Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_3459, signal_3458, signal_3457, signal_3456, signal_1200}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1186 ( .a ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930]}), .c ({signal_3463, signal_3462, signal_3461, signal_3460, signal_1201}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1187 ( .a ({signal_17187, signal_17185, signal_17183, signal_17181, signal_17179}), .b ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .c ({signal_3467, signal_3466, signal_3465, signal_3464, signal_1202}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1188 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2495, signal_2494, signal_2493, signal_2492, signal_959}), .clk ( clk ), .r ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_3471, signal_3470, signal_3469, signal_3468, signal_1203}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1191 ( .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_981}), .b ({signal_2607, signal_2606, signal_2605, signal_2604, signal_987}), .clk ( clk ), .r ({Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .c ({signal_3483, signal_3482, signal_3481, signal_3480, signal_1206}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1192 ( .a ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}), .b ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970]}), .c ({signal_3487, signal_3486, signal_3485, signal_3484, signal_1207}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1193 ( .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_957}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .clk ( clk ), .r ({Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_3491, signal_3490, signal_3489, signal_3488, signal_1208}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1194 ( .a ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990]}), .c ({signal_3495, signal_3494, signal_3493, signal_3492, signal_1209}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1195 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .c ({signal_3499, signal_3498, signal_3497, signal_3496, signal_1210}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1196 ( .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_3503, signal_3502, signal_3501, signal_3500, signal_1211}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1197 ( .a ({signal_2599, signal_2598, signal_2597, signal_2596, signal_985}), .b ({signal_2603, signal_2602, signal_2601, signal_2600, signal_986}), .clk ( clk ), .r ({Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .c ({signal_3507, signal_3506, signal_3505, signal_3504, signal_1212}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1199 ( .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_991}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_992}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030]}), .c ({signal_3515, signal_3514, signal_3513, signal_3512, signal_1214}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1200 ( .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_953}), .b ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1007}), .clk ( clk ), .r ({Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_3519, signal_3518, signal_3517, signal_3516, signal_1215}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1201 ( .a ({signal_2631, signal_2630, signal_2629, signal_2628, signal_993}), .b ({signal_2651, signal_2650, signal_2649, signal_2648, signal_998}), .clk ( clk ), .r ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050]}), .c ({signal_3523, signal_3522, signal_3521, signal_3520, signal_1216}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1202 ( .a ({signal_2611, signal_2610, signal_2609, signal_2608, signal_988}), .b ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1001}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .c ({signal_3527, signal_3526, signal_3525, signal_3524, signal_1217}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1203 ( .a ({signal_2639, signal_2638, signal_2637, signal_2636, signal_995}), .b ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .clk ( clk ), .r ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_3531, signal_3530, signal_3529, signal_3528, signal_1218}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1204 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_2615, signal_2614, signal_2613, signal_2612, signal_989}), .clk ( clk ), .r ({Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .c ({signal_3535, signal_3534, signal_3533, signal_3532, signal_1219}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1205 ( .a ({signal_17167, signal_17165, signal_17163, signal_17161, signal_17159}), .b ({signal_2647, signal_2646, signal_2645, signal_2644, signal_997}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090]}), .c ({signal_3539, signal_3538, signal_3537, signal_3536, signal_1220}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1206 ( .a ({signal_17117, signal_17115, signal_17113, signal_17111, signal_17109}), .b ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1009}), .clk ( clk ), .r ({Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_3543, signal_3542, signal_3541, signal_3540, signal_1221}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1208 ( .a ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1004}), .b ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1005}), .clk ( clk ), .r ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110]}), .c ({signal_3551, signal_3550, signal_3549, signal_3548, signal_1223}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1210 ( .a ({signal_17177, signal_17175, signal_17173, signal_17171, signal_17169}), .b ({signal_2539, signal_2538, signal_2537, signal_2536, signal_970}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .c ({signal_3559, signal_3558, signal_3557, signal_3556, signal_1225}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1213 ( .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_979}), .b ({signal_17197, signal_17195, signal_17193, signal_17191, signal_17189}), .clk ( clk ), .r ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_3571, signal_3570, signal_3569, signal_3568, signal_1228}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1214 ( .a ({signal_17177, signal_17175, signal_17173, signal_17171, signal_17169}), .b ({signal_2547, signal_2546, signal_2545, signal_2544, signal_972}), .clk ( clk ), .r ({Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .c ({signal_3575, signal_3574, signal_3573, signal_3572, signal_1229}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1215 ( .a ({signal_2935, signal_2934, signal_2933, signal_2932, signal_1069}), .b ({signal_3579, signal_3578, signal_3577, signal_3576, signal_1230}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1216 ( .a ({signal_2939, signal_2938, signal_2937, signal_2936, signal_1070}), .b ({signal_3583, signal_3582, signal_3581, signal_3580, signal_1231}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1217 ( .a ({signal_2947, signal_2946, signal_2945, signal_2944, signal_1072}), .b ({signal_3587, signal_3586, signal_3585, signal_3584, signal_1232}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1218 ( .a ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .b ({signal_3591, signal_3590, signal_3589, signal_3588, signal_1233}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1219 ( .a ({signal_2955, signal_2954, signal_2953, signal_2952, signal_1074}), .b ({signal_3595, signal_3594, signal_3593, signal_3592, signal_1234}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1220 ( .a ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .b ({signal_3599, signal_3598, signal_3597, signal_3596, signal_1235}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1221 ( .a ({signal_2963, signal_2962, signal_2961, signal_2960, signal_1076}), .b ({signal_3603, signal_3602, signal_3601, signal_3600, signal_1236}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1222 ( .a ({signal_2967, signal_2966, signal_2965, signal_2964, signal_1077}), .b ({signal_3607, signal_3606, signal_3605, signal_3604, signal_1237}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1223 ( .a ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1078}), .b ({signal_3611, signal_3610, signal_3609, signal_3608, signal_1238}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1224 ( .a ({signal_2975, signal_2974, signal_2973, signal_2972, signal_1079}), .b ({signal_3615, signal_3614, signal_3613, signal_3612, signal_1239}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1225 ( .a ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1080}), .b ({signal_3619, signal_3618, signal_3617, signal_3616, signal_1240}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1226 ( .a ({signal_2983, signal_2982, signal_2981, signal_2980, signal_1081}), .b ({signal_3623, signal_3622, signal_3621, signal_3620, signal_1241}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1227 ( .a ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}), .b ({signal_3627, signal_3626, signal_3625, signal_3624, signal_1242}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1228 ( .a ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .b ({signal_3631, signal_3630, signal_3629, signal_3628, signal_1243}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1229 ( .a ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}), .b ({signal_3635, signal_3634, signal_3633, signal_3632, signal_1244}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1230 ( .a ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}), .b ({signal_3639, signal_3638, signal_3637, signal_3636, signal_1245}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1231 ( .a ({signal_3007, signal_3006, signal_3005, signal_3004, signal_1087}), .b ({signal_3643, signal_3642, signal_3641, signal_3640, signal_1246}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1232 ( .a ({signal_3011, signal_3010, signal_3009, signal_3008, signal_1088}), .b ({signal_3647, signal_3646, signal_3645, signal_3644, signal_1247}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1233 ( .a ({signal_3019, signal_3018, signal_3017, signal_3016, signal_1090}), .b ({signal_3651, signal_3650, signal_3649, signal_3648, signal_1248}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1234 ( .a ({signal_3023, signal_3022, signal_3021, signal_3020, signal_1091}), .b ({signal_3655, signal_3654, signal_3653, signal_3652, signal_1249}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1235 ( .a ({signal_3027, signal_3026, signal_3025, signal_3024, signal_1092}), .b ({signal_3659, signal_3658, signal_3657, signal_3656, signal_1250}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1236 ( .a ({signal_3031, signal_3030, signal_3029, signal_3028, signal_1093}), .b ({signal_3663, signal_3662, signal_3661, signal_3660, signal_1251}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1237 ( .a ({signal_3035, signal_3034, signal_3033, signal_3032, signal_1094}), .b ({signal_3667, signal_3666, signal_3665, signal_3664, signal_1252}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1238 ( .a ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .b ({signal_3671, signal_3670, signal_3669, signal_3668, signal_1253}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1239 ( .a ({signal_3043, signal_3042, signal_3041, signal_3040, signal_1096}), .b ({signal_3675, signal_3674, signal_3673, signal_3672, signal_1254}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1240 ( .a ({signal_3047, signal_3046, signal_3045, signal_3044, signal_1097}), .b ({signal_3679, signal_3678, signal_3677, signal_3676, signal_1255}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1241 ( .a ({signal_3051, signal_3050, signal_3049, signal_3048, signal_1098}), .b ({signal_3683, signal_3682, signal_3681, signal_3680, signal_1256}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1242 ( .a ({signal_3055, signal_3054, signal_3053, signal_3052, signal_1099}), .b ({signal_3687, signal_3686, signal_3685, signal_3684, signal_1257}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1244 ( .a ({signal_3063, signal_3062, signal_3061, signal_3060, signal_1101}), .b ({signal_3695, signal_3694, signal_3693, signal_3692, signal_1259}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1245 ( .a ({signal_3071, signal_3070, signal_3069, signal_3068, signal_1103}), .b ({signal_3699, signal_3698, signal_3697, signal_3696, signal_1260}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1246 ( .a ({signal_3079, signal_3078, signal_3077, signal_3076, signal_1105}), .b ({signal_3703, signal_3702, signal_3701, signal_3700, signal_1261}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1247 ( .a ({signal_3083, signal_3082, signal_3081, signal_3080, signal_1106}), .b ({signal_3707, signal_3706, signal_3705, signal_3704, signal_1262}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1248 ( .a ({signal_3091, signal_3090, signal_3089, signal_3088, signal_1108}), .b ({signal_3711, signal_3710, signal_3709, signal_3708, signal_1263}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1249 ( .a ({signal_3095, signal_3094, signal_3093, signal_3092, signal_1109}), .b ({signal_3715, signal_3714, signal_3713, signal_3712, signal_1264}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1250 ( .a ({signal_3099, signal_3098, signal_3097, signal_3096, signal_1110}), .b ({signal_3719, signal_3718, signal_3717, signal_3716, signal_1265}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1251 ( .a ({signal_3103, signal_3102, signal_3101, signal_3100, signal_1111}), .b ({signal_3723, signal_3722, signal_3721, signal_3720, signal_1266}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1252 ( .a ({signal_3107, signal_3106, signal_3105, signal_3104, signal_1112}), .b ({signal_3727, signal_3726, signal_3725, signal_3724, signal_1267}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1253 ( .a ({signal_3111, signal_3110, signal_3109, signal_3108, signal_1113}), .b ({signal_3731, signal_3730, signal_3729, signal_3728, signal_1268}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1254 ( .a ({signal_3119, signal_3118, signal_3117, signal_3116, signal_1115}), .b ({signal_3735, signal_3734, signal_3733, signal_3732, signal_1269}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1255 ( .a ({signal_3123, signal_3122, signal_3121, signal_3120, signal_1116}), .b ({signal_3739, signal_3738, signal_3737, signal_3736, signal_1270}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1256 ( .a ({signal_3127, signal_3126, signal_3125, signal_3124, signal_1117}), .b ({signal_3743, signal_3742, signal_3741, signal_3740, signal_1271}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1257 ( .a ({signal_3131, signal_3130, signal_3129, signal_3128, signal_1118}), .b ({signal_3747, signal_3746, signal_3745, signal_3744, signal_1272}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1258 ( .a ({signal_3139, signal_3138, signal_3137, signal_3136, signal_1120}), .b ({signal_3751, signal_3750, signal_3749, signal_3748, signal_1273}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1259 ( .a ({signal_3143, signal_3142, signal_3141, signal_3140, signal_1121}), .b ({signal_3755, signal_3754, signal_3753, signal_3752, signal_1274}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1260 ( .a ({signal_3147, signal_3146, signal_3145, signal_3144, signal_1122}), .b ({signal_3759, signal_3758, signal_3757, signal_3756, signal_1275}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1261 ( .a ({signal_3155, signal_3154, signal_3153, signal_3152, signal_1124}), .b ({signal_3763, signal_3762, signal_3761, signal_3760, signal_1276}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1262 ( .a ({signal_3159, signal_3158, signal_3157, signal_3156, signal_1125}), .b ({signal_3767, signal_3766, signal_3765, signal_3764, signal_1277}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1263 ( .a ({signal_3163, signal_3162, signal_3161, signal_3160, signal_1126}), .b ({signal_3771, signal_3770, signal_3769, signal_3768, signal_1278}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1264 ( .a ({signal_3167, signal_3166, signal_3165, signal_3164, signal_1127}), .b ({signal_3775, signal_3774, signal_3773, signal_3772, signal_1279}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1265 ( .a ({signal_3175, signal_3174, signal_3173, signal_3172, signal_1129}), .b ({signal_3779, signal_3778, signal_3777, signal_3776, signal_1280}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1266 ( .a ({signal_3179, signal_3178, signal_3177, signal_3176, signal_1130}), .b ({signal_3783, signal_3782, signal_3781, signal_3780, signal_1281}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1267 ( .a ({signal_3183, signal_3182, signal_3181, signal_3180, signal_1131}), .b ({signal_3787, signal_3786, signal_3785, signal_3784, signal_1282}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1268 ( .a ({signal_3195, signal_3194, signal_3193, signal_3192, signal_1134}), .b ({signal_3791, signal_3790, signal_3789, signal_3788, signal_1283}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1269 ( .a ({signal_3199, signal_3198, signal_3197, signal_3196, signal_1135}), .b ({signal_3795, signal_3794, signal_3793, signal_3792, signal_1284}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1270 ( .a ({signal_3203, signal_3202, signal_3201, signal_3200, signal_1136}), .b ({signal_3799, signal_3798, signal_3797, signal_3796, signal_1285}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1271 ( .a ({signal_3207, signal_3206, signal_3205, signal_3204, signal_1137}), .b ({signal_3803, signal_3802, signal_3801, signal_3800, signal_1286}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1273 ( .a ({signal_3223, signal_3222, signal_3221, signal_3220, signal_1141}), .b ({signal_3811, signal_3810, signal_3809, signal_3808, signal_1288}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1274 ( .a ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .b ({signal_3815, signal_3814, signal_3813, signal_3812, signal_1289}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1275 ( .a ({signal_3235, signal_3234, signal_3233, signal_3232, signal_1144}), .b ({signal_3819, signal_3818, signal_3817, signal_3816, signal_1290}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1276 ( .a ({signal_3243, signal_3242, signal_3241, signal_3240, signal_1146}), .b ({signal_3823, signal_3822, signal_3821, signal_3820, signal_1291}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1278 ( .a ({signal_3251, signal_3250, signal_3249, signal_3248, signal_1148}), .b ({signal_3831, signal_3830, signal_3829, signal_3828, signal_1293}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1279 ( .a ({signal_3255, signal_3254, signal_3253, signal_3252, signal_1149}), .b ({signal_3835, signal_3834, signal_3833, signal_3832, signal_1294}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1280 ( .a ({signal_3259, signal_3258, signal_3257, signal_3256, signal_1150}), .b ({signal_3839, signal_3838, signal_3837, signal_3836, signal_1295}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1281 ( .a ({signal_3267, signal_3266, signal_3265, signal_3264, signal_1152}), .b ({signal_3843, signal_3842, signal_3841, signal_3840, signal_1296}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1282 ( .a ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .b ({signal_3847, signal_3846, signal_3845, signal_3844, signal_1297}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1283 ( .a ({signal_3275, signal_3274, signal_3273, signal_3272, signal_1154}), .b ({signal_3851, signal_3850, signal_3849, signal_3848, signal_1298}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1285 ( .a ({signal_3283, signal_3282, signal_3281, signal_3280, signal_1156}), .b ({signal_3859, signal_3858, signal_3857, signal_3856, signal_1300}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1286 ( .a ({signal_3287, signal_3286, signal_3285, signal_3284, signal_1157}), .b ({signal_3863, signal_3862, signal_3861, signal_3860, signal_1301}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1287 ( .a ({signal_3295, signal_3294, signal_3293, signal_3292, signal_1159}), .b ({signal_3867, signal_3866, signal_3865, signal_3864, signal_1302}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1288 ( .a ({signal_3299, signal_3298, signal_3297, signal_3296, signal_1160}), .b ({signal_3871, signal_3870, signal_3869, signal_3868, signal_1303}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1289 ( .a ({signal_3303, signal_3302, signal_3301, signal_3300, signal_1161}), .b ({signal_3875, signal_3874, signal_3873, signal_3872, signal_1304}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1290 ( .a ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .b ({signal_3879, signal_3878, signal_3877, signal_3876, signal_1305}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1291 ( .a ({signal_3311, signal_3310, signal_3309, signal_3308, signal_1163}), .b ({signal_3883, signal_3882, signal_3881, signal_3880, signal_1306}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1292 ( .a ({signal_3315, signal_3314, signal_3313, signal_3312, signal_1164}), .b ({signal_3887, signal_3886, signal_3885, signal_3884, signal_1307}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1293 ( .a ({signal_3319, signal_3318, signal_3317, signal_3316, signal_1165}), .b ({signal_3891, signal_3890, signal_3889, signal_3888, signal_1308}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1294 ( .a ({signal_3323, signal_3322, signal_3321, signal_3320, signal_1166}), .b ({signal_3895, signal_3894, signal_3893, signal_3892, signal_1309}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1295 ( .a ({signal_3327, signal_3326, signal_3325, signal_3324, signal_1167}), .b ({signal_3899, signal_3898, signal_3897, signal_3896, signal_1310}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1296 ( .a ({signal_3335, signal_3334, signal_3333, signal_3332, signal_1169}), .b ({signal_3903, signal_3902, signal_3901, signal_3900, signal_1311}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1298 ( .a ({signal_3343, signal_3342, signal_3341, signal_3340, signal_1171}), .b ({signal_3911, signal_3910, signal_3909, signal_3908, signal_1313}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1299 ( .a ({signal_3347, signal_3346, signal_3345, signal_3344, signal_1172}), .b ({signal_3915, signal_3914, signal_3913, signal_3912, signal_1314}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1300 ( .a ({signal_3351, signal_3350, signal_3349, signal_3348, signal_1173}), .b ({signal_3919, signal_3918, signal_3917, signal_3916, signal_1315}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1301 ( .a ({signal_3355, signal_3354, signal_3353, signal_3352, signal_1174}), .b ({signal_3923, signal_3922, signal_3921, signal_3920, signal_1316}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1302 ( .a ({signal_3359, signal_3358, signal_3357, signal_3356, signal_1175}), .b ({signal_3927, signal_3926, signal_3925, signal_3924, signal_1317}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1303 ( .a ({signal_3363, signal_3362, signal_3361, signal_3360, signal_1176}), .b ({signal_3931, signal_3930, signal_3929, signal_3928, signal_1318}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1304 ( .a ({signal_3367, signal_3366, signal_3365, signal_3364, signal_1177}), .b ({signal_3935, signal_3934, signal_3933, signal_3932, signal_1319}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1305 ( .a ({signal_3375, signal_3374, signal_3373, signal_3372, signal_1179}), .b ({signal_3939, signal_3938, signal_3937, signal_3936, signal_1320}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1306 ( .a ({signal_3379, signal_3378, signal_3377, signal_3376, signal_1180}), .b ({signal_3943, signal_3942, signal_3941, signal_3940, signal_1321}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1307 ( .a ({signal_3383, signal_3382, signal_3381, signal_3380, signal_1181}), .b ({signal_3947, signal_3946, signal_3945, signal_3944, signal_1322}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1308 ( .a ({signal_3387, signal_3386, signal_3385, signal_3384, signal_1182}), .b ({signal_3951, signal_3950, signal_3949, signal_3948, signal_1323}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1309 ( .a ({signal_3391, signal_3390, signal_3389, signal_3388, signal_1183}), .b ({signal_3955, signal_3954, signal_3953, signal_3952, signal_1324}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1310 ( .a ({signal_3395, signal_3394, signal_3393, signal_3392, signal_1184}), .b ({signal_3959, signal_3958, signal_3957, signal_3956, signal_1325}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1311 ( .a ({signal_3399, signal_3398, signal_3397, signal_3396, signal_1185}), .b ({signal_3963, signal_3962, signal_3961, signal_3960, signal_1326}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1312 ( .a ({signal_3403, signal_3402, signal_3401, signal_3400, signal_1186}), .b ({signal_3967, signal_3966, signal_3965, signal_3964, signal_1327}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1313 ( .a ({signal_3407, signal_3406, signal_3405, signal_3404, signal_1187}), .b ({signal_3971, signal_3970, signal_3969, signal_3968, signal_1328}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1315 ( .a ({signal_3415, signal_3414, signal_3413, signal_3412, signal_1189}), .b ({signal_3979, signal_3978, signal_3977, signal_3976, signal_1330}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1316 ( .a ({signal_3423, signal_3422, signal_3421, signal_3420, signal_1191}), .b ({signal_3983, signal_3982, signal_3981, signal_3980, signal_1331}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1317 ( .a ({signal_3427, signal_3426, signal_3425, signal_3424, signal_1192}), .b ({signal_3987, signal_3986, signal_3985, signal_3984, signal_1332}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1318 ( .a ({signal_3431, signal_3430, signal_3429, signal_3428, signal_1193}), .b ({signal_3991, signal_3990, signal_3989, signal_3988, signal_1333}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1319 ( .a ({signal_3435, signal_3434, signal_3433, signal_3432, signal_1194}), .b ({signal_3995, signal_3994, signal_3993, signal_3992, signal_1334}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1320 ( .a ({signal_3439, signal_3438, signal_3437, signal_3436, signal_1195}), .b ({signal_3999, signal_3998, signal_3997, signal_3996, signal_1335}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1321 ( .a ({signal_3443, signal_3442, signal_3441, signal_3440, signal_1196}), .b ({signal_4003, signal_4002, signal_4001, signal_4000, signal_1336}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1322 ( .a ({signal_3447, signal_3446, signal_3445, signal_3444, signal_1197}), .b ({signal_4007, signal_4006, signal_4005, signal_4004, signal_1337}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1324 ( .a ({signal_3459, signal_3458, signal_3457, signal_3456, signal_1200}), .b ({signal_4015, signal_4014, signal_4013, signal_4012, signal_1339}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1325 ( .a ({signal_3463, signal_3462, signal_3461, signal_3460, signal_1201}), .b ({signal_4019, signal_4018, signal_4017, signal_4016, signal_1340}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1326 ( .a ({signal_3467, signal_3466, signal_3465, signal_3464, signal_1202}), .b ({signal_4023, signal_4022, signal_4021, signal_4020, signal_1341}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1327 ( .a ({signal_3471, signal_3470, signal_3469, signal_3468, signal_1203}), .b ({signal_4027, signal_4026, signal_4025, signal_4024, signal_1342}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1330 ( .a ({signal_3487, signal_3486, signal_3485, signal_3484, signal_1207}), .b ({signal_4039, signal_4038, signal_4037, signal_4036, signal_1345}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1331 ( .a ({signal_3495, signal_3494, signal_3493, signal_3492, signal_1209}), .b ({signal_4043, signal_4042, signal_4041, signal_4040, signal_1346}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1332 ( .a ({signal_3499, signal_3498, signal_3497, signal_3496, signal_1210}), .b ({signal_4047, signal_4046, signal_4045, signal_4044, signal_1347}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1333 ( .a ({signal_3503, signal_3502, signal_3501, signal_3500, signal_1211}), .b ({signal_4051, signal_4050, signal_4049, signal_4048, signal_1348}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1334 ( .a ({signal_3507, signal_3506, signal_3505, signal_3504, signal_1212}), .b ({signal_4055, signal_4054, signal_4053, signal_4052, signal_1349}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1336 ( .a ({signal_3515, signal_3514, signal_3513, signal_3512, signal_1214}), .b ({signal_4063, signal_4062, signal_4061, signal_4060, signal_1351}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1337 ( .a ({signal_3519, signal_3518, signal_3517, signal_3516, signal_1215}), .b ({signal_4067, signal_4066, signal_4065, signal_4064, signal_1352}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1338 ( .a ({signal_3523, signal_3522, signal_3521, signal_3520, signal_1216}), .b ({signal_4071, signal_4070, signal_4069, signal_4068, signal_1353}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1339 ( .a ({signal_3531, signal_3530, signal_3529, signal_3528, signal_1218}), .b ({signal_4075, signal_4074, signal_4073, signal_4072, signal_1354}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1340 ( .a ({signal_3535, signal_3534, signal_3533, signal_3532, signal_1219}), .b ({signal_4079, signal_4078, signal_4077, signal_4076, signal_1355}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1341 ( .a ({signal_3539, signal_3538, signal_3537, signal_3536, signal_1220}), .b ({signal_4083, signal_4082, signal_4081, signal_4080, signal_1356}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1342 ( .a ({signal_3543, signal_3542, signal_3541, signal_3540, signal_1221}), .b ({signal_4087, signal_4086, signal_4085, signal_4084, signal_1357}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1344 ( .a ({signal_3551, signal_3550, signal_3549, signal_3548, signal_1223}), .b ({signal_4095, signal_4094, signal_4093, signal_4092, signal_1359}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1346 ( .a ({signal_3559, signal_3558, signal_3557, signal_3556, signal_1225}), .b ({signal_4103, signal_4102, signal_4101, signal_4100, signal_1361}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1349 ( .a ({signal_3571, signal_3570, signal_3569, signal_3568, signal_1228}), .b ({signal_4115, signal_4114, signal_4113, signal_4112, signal_1364}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1350 ( .a ({signal_3575, signal_3574, signal_3573, signal_3572, signal_1229}), .b ({signal_4119, signal_4118, signal_4117, signal_4116, signal_1365}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1353 ( .a ({signal_17207, signal_17205, signal_17203, signal_17201, signal_17199}), .b ({signal_2843, signal_2842, signal_2841, signal_2840, signal_1046}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150]}), .c ({signal_4131, signal_4130, signal_4129, signal_4128, signal_1368}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1354 ( .a ({signal_17157, signal_17155, signal_17153, signal_17151, signal_17149}), .b ({signal_2827, signal_2826, signal_2825, signal_2824, signal_1042}), .clk ( clk ), .r ({Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_4135, signal_4134, signal_4133, signal_4132, signal_1369}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1355 ( .a ({signal_2783, signal_2782, signal_2781, signal_2780, signal_1031}), .b ({signal_2891, signal_2890, signal_2889, signal_2888, signal_1058}), .clk ( clk ), .r ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170]}), .c ({signal_4139, signal_4138, signal_4137, signal_4136, signal_1370}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1356 ( .a ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}), .b ({signal_2887, signal_2886, signal_2885, signal_2884, signal_1057}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .c ({signal_4143, signal_4142, signal_4141, signal_4140, signal_1371}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1357 ( .a ({signal_2803, signal_2802, signal_2801, signal_2800, signal_1036}), .b ({signal_2807, signal_2806, signal_2805, signal_2804, signal_1037}), .clk ( clk ), .r ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_4147, signal_4146, signal_4145, signal_4144, signal_1372}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1360 ( .a ({signal_2803, signal_2802, signal_2801, signal_2800, signal_1036}), .b ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}), .clk ( clk ), .r ({Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .c ({signal_4159, signal_4158, signal_4157, signal_4156, signal_1375}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1361 ( .a ({signal_2823, signal_2822, signal_2821, signal_2820, signal_1041}), .b ({signal_2867, signal_2866, signal_2865, signal_2864, signal_1052}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210]}), .c ({signal_4163, signal_4162, signal_4161, signal_4160, signal_1376}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1362 ( .a ({signal_2863, signal_2862, signal_2861, signal_2860, signal_1051}), .b ({signal_2871, signal_2870, signal_2869, signal_2868, signal_1053}), .clk ( clk ), .r ({Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_4167, signal_4166, signal_4165, signal_4164, signal_1377}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1365 ( .a ({signal_2783, signal_2782, signal_2781, signal_2780, signal_1031}), .b ({signal_2835, signal_2834, signal_2833, signal_2832, signal_1044}), .clk ( clk ), .r ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230]}), .c ({signal_4179, signal_4178, signal_4177, signal_4176, signal_1380}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1366 ( .a ({signal_2787, signal_2786, signal_2785, signal_2784, signal_1032}), .b ({signal_2867, signal_2866, signal_2865, signal_2864, signal_1052}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .c ({signal_4183, signal_4182, signal_4181, signal_4180, signal_1381}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1367 ( .a ({signal_2827, signal_2826, signal_2825, signal_2824, signal_1042}), .b ({signal_2831, signal_2830, signal_2829, signal_2828, signal_1043}), .clk ( clk ), .r ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_4187, signal_4186, signal_4185, signal_4184, signal_1382}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1368 ( .a ({signal_2807, signal_2806, signal_2805, signal_2804, signal_1037}), .b ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}), .clk ( clk ), .r ({Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .c ({signal_4191, signal_4190, signal_4189, signal_4188, signal_1383}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1369 ( .a ({signal_2555, signal_2554, signal_2553, signal_2552, signal_974}), .b ({signal_2871, signal_2870, signal_2869, signal_2868, signal_1053}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270]}), .c ({signal_4195, signal_4194, signal_4193, signal_4192, signal_1384}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1375 ( .a ({signal_2819, signal_2818, signal_2817, signal_2816, signal_1040}), .b ({signal_2883, signal_2882, signal_2881, signal_2880, signal_1056}), .clk ( clk ), .r ({Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_4219, signal_4218, signal_4217, signal_4216, signal_1390}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1376 ( .a ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}), .b ({signal_2859, signal_2858, signal_2857, signal_2856, signal_1050}), .clk ( clk ), .r ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290]}), .c ({signal_4223, signal_4222, signal_4221, signal_4220, signal_1391}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1383 ( .a ({signal_2791, signal_2790, signal_2789, signal_2788, signal_1033}), .b ({signal_2799, signal_2798, signal_2797, signal_2796, signal_1035}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .c ({signal_4251, signal_4250, signal_4249, signal_4248, signal_1398}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1395 ( .a ({signal_2543, signal_2542, signal_2541, signal_2540, signal_971}), .b ({signal_2855, signal_2854, signal_2853, signal_2852, signal_1049}), .clk ( clk ), .r ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_4299, signal_4298, signal_4297, signal_4296, signal_1410}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1396 ( .a ({signal_2787, signal_2786, signal_2785, signal_2784, signal_1032}), .b ({signal_2847, signal_2846, signal_2845, signal_2844, signal_1047}), .clk ( clk ), .r ({Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .c ({signal_4303, signal_4302, signal_4301, signal_4300, signal_1411}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1401 ( .a ({signal_2527, signal_2526, signal_2525, signal_2524, signal_967}), .b ({signal_2831, signal_2830, signal_2829, signal_2828, signal_1043}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330]}), .c ({signal_4323, signal_4322, signal_4321, signal_4320, signal_1416}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1402 ( .a ({signal_2859, signal_2858, signal_2857, signal_2856, signal_1050}), .b ({signal_2559, signal_2558, signal_2557, signal_2556, signal_975}), .clk ( clk ), .r ({Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_4327, signal_4326, signal_4325, signal_4324, signal_1417}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1403 ( .a ({signal_2547, signal_2546, signal_2545, signal_2544, signal_972}), .b ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1045}), .clk ( clk ), .r ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350]}), .c ({signal_4331, signal_4330, signal_4329, signal_4328, signal_1418}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1407 ( .a ({signal_2811, signal_2810, signal_2809, signal_2808, signal_1038}), .b ({signal_2843, signal_2842, signal_2841, signal_2840, signal_1046}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .c ({signal_4347, signal_4346, signal_4345, signal_4344, signal_1422}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1408 ( .a ({signal_2819, signal_2818, signal_2817, signal_2816, signal_1040}), .b ({signal_2559, signal_2558, signal_2557, signal_2556, signal_975}), .clk ( clk ), .r ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_4351, signal_4350, signal_4349, signal_4348, signal_1423}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1492 ( .a ({signal_4131, signal_4130, signal_4129, signal_4128, signal_1368}), .b ({signal_4687, signal_4686, signal_4685, signal_4684, signal_1507}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1493 ( .a ({signal_4135, signal_4134, signal_4133, signal_4132, signal_1369}), .b ({signal_4691, signal_4690, signal_4689, signal_4688, signal_1508}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1494 ( .a ({signal_4139, signal_4138, signal_4137, signal_4136, signal_1370}), .b ({signal_4695, signal_4694, signal_4693, signal_4692, signal_1509}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1495 ( .a ({signal_4143, signal_4142, signal_4141, signal_4140, signal_1371}), .b ({signal_4699, signal_4698, signal_4697, signal_4696, signal_1510}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1496 ( .a ({signal_4147, signal_4146, signal_4145, signal_4144, signal_1372}), .b ({signal_4703, signal_4702, signal_4701, signal_4700, signal_1511}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1499 ( .a ({signal_4159, signal_4158, signal_4157, signal_4156, signal_1375}), .b ({signal_4715, signal_4714, signal_4713, signal_4712, signal_1514}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1500 ( .a ({signal_4163, signal_4162, signal_4161, signal_4160, signal_1376}), .b ({signal_4719, signal_4718, signal_4717, signal_4716, signal_1515}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1501 ( .a ({signal_4167, signal_4166, signal_4165, signal_4164, signal_1377}), .b ({signal_4723, signal_4722, signal_4721, signal_4720, signal_1516}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1504 ( .a ({signal_4179, signal_4178, signal_4177, signal_4176, signal_1380}), .b ({signal_4735, signal_4734, signal_4733, signal_4732, signal_1519}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1505 ( .a ({signal_4183, signal_4182, signal_4181, signal_4180, signal_1381}), .b ({signal_4739, signal_4738, signal_4737, signal_4736, signal_1520}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1506 ( .a ({signal_4187, signal_4186, signal_4185, signal_4184, signal_1382}), .b ({signal_4743, signal_4742, signal_4741, signal_4740, signal_1521}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1507 ( .a ({signal_4195, signal_4194, signal_4193, signal_4192, signal_1384}), .b ({signal_4747, signal_4746, signal_4745, signal_4744, signal_1522}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1513 ( .a ({signal_4223, signal_4222, signal_4221, signal_4220, signal_1391}), .b ({signal_4771, signal_4770, signal_4769, signal_4768, signal_1528}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1520 ( .a ({signal_4251, signal_4250, signal_4249, signal_4248, signal_1398}), .b ({signal_4799, signal_4798, signal_4797, signal_4796, signal_1535}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1532 ( .a ({signal_4299, signal_4298, signal_4297, signal_4296, signal_1410}), .b ({signal_4847, signal_4846, signal_4845, signal_4844, signal_1547}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1533 ( .a ({signal_4303, signal_4302, signal_4301, signal_4300, signal_1411}), .b ({signal_4851, signal_4850, signal_4849, signal_4848, signal_1548}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1538 ( .a ({signal_4323, signal_4322, signal_4321, signal_4320, signal_1416}), .b ({signal_4871, signal_4870, signal_4869, signal_4868, signal_1553}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1539 ( .a ({signal_4327, signal_4326, signal_4325, signal_4324, signal_1417}), .b ({signal_4875, signal_4874, signal_4873, signal_4872, signal_1554}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1543 ( .a ({signal_4347, signal_4346, signal_4345, signal_4344, signal_1422}), .b ({signal_4891, signal_4890, signal_4889, signal_4888, signal_1558}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1544 ( .a ({signal_4351, signal_4350, signal_4349, signal_4348, signal_1423}), .b ({signal_4895, signal_4894, signal_4893, signal_4892, signal_1559}) ) ;
    buf_clk cell_2518 ( .C ( clk ), .D ( signal_17210 ), .Q ( signal_17211 ) ) ;
    buf_clk cell_2522 ( .C ( clk ), .D ( signal_17214 ), .Q ( signal_17215 ) ) ;
    buf_clk cell_2526 ( .C ( clk ), .D ( signal_17218 ), .Q ( signal_17219 ) ) ;
    buf_clk cell_2530 ( .C ( clk ), .D ( signal_17222 ), .Q ( signal_17223 ) ) ;
    buf_clk cell_2534 ( .C ( clk ), .D ( signal_17226 ), .Q ( signal_17227 ) ) ;
    buf_clk cell_2536 ( .C ( clk ), .D ( signal_17228 ), .Q ( signal_17229 ) ) ;
    buf_clk cell_2538 ( .C ( clk ), .D ( signal_17230 ), .Q ( signal_17231 ) ) ;
    buf_clk cell_2540 ( .C ( clk ), .D ( signal_17232 ), .Q ( signal_17233 ) ) ;
    buf_clk cell_2542 ( .C ( clk ), .D ( signal_17234 ), .Q ( signal_17235 ) ) ;
    buf_clk cell_2544 ( .C ( clk ), .D ( signal_17236 ), .Q ( signal_17237 ) ) ;
    buf_clk cell_2546 ( .C ( clk ), .D ( signal_17238 ), .Q ( signal_17239 ) ) ;
    buf_clk cell_2548 ( .C ( clk ), .D ( signal_17240 ), .Q ( signal_17241 ) ) ;
    buf_clk cell_2550 ( .C ( clk ), .D ( signal_17242 ), .Q ( signal_17243 ) ) ;
    buf_clk cell_2552 ( .C ( clk ), .D ( signal_17244 ), .Q ( signal_17245 ) ) ;
    buf_clk cell_2554 ( .C ( clk ), .D ( signal_17246 ), .Q ( signal_17247 ) ) ;
    buf_clk cell_2556 ( .C ( clk ), .D ( signal_17248 ), .Q ( signal_17249 ) ) ;
    buf_clk cell_2558 ( .C ( clk ), .D ( signal_17250 ), .Q ( signal_17251 ) ) ;
    buf_clk cell_2560 ( .C ( clk ), .D ( signal_17252 ), .Q ( signal_17253 ) ) ;
    buf_clk cell_2562 ( .C ( clk ), .D ( signal_17254 ), .Q ( signal_17255 ) ) ;
    buf_clk cell_2564 ( .C ( clk ), .D ( signal_17256 ), .Q ( signal_17257 ) ) ;
    buf_clk cell_2566 ( .C ( clk ), .D ( signal_17258 ), .Q ( signal_17259 ) ) ;
    buf_clk cell_2568 ( .C ( clk ), .D ( signal_17260 ), .Q ( signal_17261 ) ) ;
    buf_clk cell_2570 ( .C ( clk ), .D ( signal_17262 ), .Q ( signal_17263 ) ) ;
    buf_clk cell_2572 ( .C ( clk ), .D ( signal_17264 ), .Q ( signal_17265 ) ) ;
    buf_clk cell_2574 ( .C ( clk ), .D ( signal_17266 ), .Q ( signal_17267 ) ) ;
    buf_clk cell_2576 ( .C ( clk ), .D ( signal_17268 ), .Q ( signal_17269 ) ) ;
    buf_clk cell_2578 ( .C ( clk ), .D ( signal_17270 ), .Q ( signal_17271 ) ) ;
    buf_clk cell_2580 ( .C ( clk ), .D ( signal_17272 ), .Q ( signal_17273 ) ) ;
    buf_clk cell_2582 ( .C ( clk ), .D ( signal_17274 ), .Q ( signal_17275 ) ) ;
    buf_clk cell_2584 ( .C ( clk ), .D ( signal_17276 ), .Q ( signal_17277 ) ) ;
    buf_clk cell_2586 ( .C ( clk ), .D ( signal_17278 ), .Q ( signal_17279 ) ) ;
    buf_clk cell_2588 ( .C ( clk ), .D ( signal_17280 ), .Q ( signal_17281 ) ) ;
    buf_clk cell_2590 ( .C ( clk ), .D ( signal_17282 ), .Q ( signal_17283 ) ) ;
    buf_clk cell_2592 ( .C ( clk ), .D ( signal_17284 ), .Q ( signal_17285 ) ) ;
    buf_clk cell_2594 ( .C ( clk ), .D ( signal_17286 ), .Q ( signal_17287 ) ) ;
    buf_clk cell_2596 ( .C ( clk ), .D ( signal_17288 ), .Q ( signal_17289 ) ) ;
    buf_clk cell_2598 ( .C ( clk ), .D ( signal_17290 ), .Q ( signal_17291 ) ) ;
    buf_clk cell_2600 ( .C ( clk ), .D ( signal_17292 ), .Q ( signal_17293 ) ) ;
    buf_clk cell_2602 ( .C ( clk ), .D ( signal_17294 ), .Q ( signal_17295 ) ) ;
    buf_clk cell_2604 ( .C ( clk ), .D ( signal_17296 ), .Q ( signal_17297 ) ) ;
    buf_clk cell_2606 ( .C ( clk ), .D ( signal_17298 ), .Q ( signal_17299 ) ) ;
    buf_clk cell_2608 ( .C ( clk ), .D ( signal_17300 ), .Q ( signal_17301 ) ) ;
    buf_clk cell_2610 ( .C ( clk ), .D ( signal_17302 ), .Q ( signal_17303 ) ) ;
    buf_clk cell_2612 ( .C ( clk ), .D ( signal_17304 ), .Q ( signal_17305 ) ) ;
    buf_clk cell_2614 ( .C ( clk ), .D ( signal_17306 ), .Q ( signal_17307 ) ) ;
    buf_clk cell_2616 ( .C ( clk ), .D ( signal_17308 ), .Q ( signal_17309 ) ) ;
    buf_clk cell_2618 ( .C ( clk ), .D ( signal_17310 ), .Q ( signal_17311 ) ) ;
    buf_clk cell_2620 ( .C ( clk ), .D ( signal_17312 ), .Q ( signal_17313 ) ) ;
    buf_clk cell_2622 ( .C ( clk ), .D ( signal_17314 ), .Q ( signal_17315 ) ) ;
    buf_clk cell_2624 ( .C ( clk ), .D ( signal_17316 ), .Q ( signal_17317 ) ) ;
    buf_clk cell_2626 ( .C ( clk ), .D ( signal_17318 ), .Q ( signal_17319 ) ) ;
    buf_clk cell_2628 ( .C ( clk ), .D ( signal_17320 ), .Q ( signal_17321 ) ) ;
    buf_clk cell_2630 ( .C ( clk ), .D ( signal_17322 ), .Q ( signal_17323 ) ) ;
    buf_clk cell_2632 ( .C ( clk ), .D ( signal_17324 ), .Q ( signal_17325 ) ) ;
    buf_clk cell_2634 ( .C ( clk ), .D ( signal_17326 ), .Q ( signal_17327 ) ) ;
    buf_clk cell_2636 ( .C ( clk ), .D ( signal_17328 ), .Q ( signal_17329 ) ) ;
    buf_clk cell_2638 ( .C ( clk ), .D ( signal_17330 ), .Q ( signal_17331 ) ) ;
    buf_clk cell_2640 ( .C ( clk ), .D ( signal_17332 ), .Q ( signal_17333 ) ) ;
    buf_clk cell_2642 ( .C ( clk ), .D ( signal_17334 ), .Q ( signal_17335 ) ) ;
    buf_clk cell_2644 ( .C ( clk ), .D ( signal_17336 ), .Q ( signal_17337 ) ) ;
    buf_clk cell_2646 ( .C ( clk ), .D ( signal_17338 ), .Q ( signal_17339 ) ) ;
    buf_clk cell_2648 ( .C ( clk ), .D ( signal_17340 ), .Q ( signal_17341 ) ) ;
    buf_clk cell_2650 ( .C ( clk ), .D ( signal_17342 ), .Q ( signal_17343 ) ) ;
    buf_clk cell_2652 ( .C ( clk ), .D ( signal_17344 ), .Q ( signal_17345 ) ) ;
    buf_clk cell_2654 ( .C ( clk ), .D ( signal_17346 ), .Q ( signal_17347 ) ) ;
    buf_clk cell_2656 ( .C ( clk ), .D ( signal_17348 ), .Q ( signal_17349 ) ) ;
    buf_clk cell_2658 ( .C ( clk ), .D ( signal_17350 ), .Q ( signal_17351 ) ) ;
    buf_clk cell_2660 ( .C ( clk ), .D ( signal_17352 ), .Q ( signal_17353 ) ) ;
    buf_clk cell_2662 ( .C ( clk ), .D ( signal_17354 ), .Q ( signal_17355 ) ) ;
    buf_clk cell_2664 ( .C ( clk ), .D ( signal_17356 ), .Q ( signal_17357 ) ) ;
    buf_clk cell_2666 ( .C ( clk ), .D ( signal_17358 ), .Q ( signal_17359 ) ) ;
    buf_clk cell_2668 ( .C ( clk ), .D ( signal_17360 ), .Q ( signal_17361 ) ) ;
    buf_clk cell_2670 ( .C ( clk ), .D ( signal_17362 ), .Q ( signal_17363 ) ) ;
    buf_clk cell_2672 ( .C ( clk ), .D ( signal_17364 ), .Q ( signal_17365 ) ) ;
    buf_clk cell_2674 ( .C ( clk ), .D ( signal_17366 ), .Q ( signal_17367 ) ) ;
    buf_clk cell_2676 ( .C ( clk ), .D ( signal_17368 ), .Q ( signal_17369 ) ) ;
    buf_clk cell_2678 ( .C ( clk ), .D ( signal_17370 ), .Q ( signal_17371 ) ) ;
    buf_clk cell_2680 ( .C ( clk ), .D ( signal_17372 ), .Q ( signal_17373 ) ) ;
    buf_clk cell_2682 ( .C ( clk ), .D ( signal_17374 ), .Q ( signal_17375 ) ) ;
    buf_clk cell_2684 ( .C ( clk ), .D ( signal_17376 ), .Q ( signal_17377 ) ) ;
    buf_clk cell_2686 ( .C ( clk ), .D ( signal_17378 ), .Q ( signal_17379 ) ) ;
    buf_clk cell_2688 ( .C ( clk ), .D ( signal_17380 ), .Q ( signal_17381 ) ) ;
    buf_clk cell_2690 ( .C ( clk ), .D ( signal_17382 ), .Q ( signal_17383 ) ) ;
    buf_clk cell_2692 ( .C ( clk ), .D ( signal_17384 ), .Q ( signal_17385 ) ) ;
    buf_clk cell_2694 ( .C ( clk ), .D ( signal_17386 ), .Q ( signal_17387 ) ) ;
    buf_clk cell_2696 ( .C ( clk ), .D ( signal_17388 ), .Q ( signal_17389 ) ) ;
    buf_clk cell_2698 ( .C ( clk ), .D ( signal_17390 ), .Q ( signal_17391 ) ) ;
    buf_clk cell_2700 ( .C ( clk ), .D ( signal_17392 ), .Q ( signal_17393 ) ) ;
    buf_clk cell_2702 ( .C ( clk ), .D ( signal_17394 ), .Q ( signal_17395 ) ) ;
    buf_clk cell_2704 ( .C ( clk ), .D ( signal_17396 ), .Q ( signal_17397 ) ) ;
    buf_clk cell_2706 ( .C ( clk ), .D ( signal_17398 ), .Q ( signal_17399 ) ) ;
    buf_clk cell_2708 ( .C ( clk ), .D ( signal_17400 ), .Q ( signal_17401 ) ) ;
    buf_clk cell_2710 ( .C ( clk ), .D ( signal_17402 ), .Q ( signal_17403 ) ) ;
    buf_clk cell_2712 ( .C ( clk ), .D ( signal_17404 ), .Q ( signal_17405 ) ) ;
    buf_clk cell_2714 ( .C ( clk ), .D ( signal_17406 ), .Q ( signal_17407 ) ) ;
    buf_clk cell_2716 ( .C ( clk ), .D ( signal_17408 ), .Q ( signal_17409 ) ) ;
    buf_clk cell_2718 ( .C ( clk ), .D ( signal_17410 ), .Q ( signal_17411 ) ) ;
    buf_clk cell_2720 ( .C ( clk ), .D ( signal_17412 ), .Q ( signal_17413 ) ) ;
    buf_clk cell_2722 ( .C ( clk ), .D ( signal_17414 ), .Q ( signal_17415 ) ) ;
    buf_clk cell_2724 ( .C ( clk ), .D ( signal_17416 ), .Q ( signal_17417 ) ) ;
    buf_clk cell_2726 ( .C ( clk ), .D ( signal_17418 ), .Q ( signal_17419 ) ) ;
    buf_clk cell_2728 ( .C ( clk ), .D ( signal_17420 ), .Q ( signal_17421 ) ) ;
    buf_clk cell_2730 ( .C ( clk ), .D ( signal_17422 ), .Q ( signal_17423 ) ) ;
    buf_clk cell_2732 ( .C ( clk ), .D ( signal_17424 ), .Q ( signal_17425 ) ) ;
    buf_clk cell_2734 ( .C ( clk ), .D ( signal_17426 ), .Q ( signal_17427 ) ) ;
    buf_clk cell_2736 ( .C ( clk ), .D ( signal_17428 ), .Q ( signal_17429 ) ) ;
    buf_clk cell_2738 ( .C ( clk ), .D ( signal_17430 ), .Q ( signal_17431 ) ) ;
    buf_clk cell_2740 ( .C ( clk ), .D ( signal_17432 ), .Q ( signal_17433 ) ) ;
    buf_clk cell_2742 ( .C ( clk ), .D ( signal_17434 ), .Q ( signal_17435 ) ) ;
    buf_clk cell_2744 ( .C ( clk ), .D ( signal_17436 ), .Q ( signal_17437 ) ) ;
    buf_clk cell_2746 ( .C ( clk ), .D ( signal_17438 ), .Q ( signal_17439 ) ) ;
    buf_clk cell_2748 ( .C ( clk ), .D ( signal_17440 ), .Q ( signal_17441 ) ) ;
    buf_clk cell_2750 ( .C ( clk ), .D ( signal_17442 ), .Q ( signal_17443 ) ) ;
    buf_clk cell_2752 ( .C ( clk ), .D ( signal_17444 ), .Q ( signal_17445 ) ) ;
    buf_clk cell_2754 ( .C ( clk ), .D ( signal_17446 ), .Q ( signal_17447 ) ) ;
    buf_clk cell_2756 ( .C ( clk ), .D ( signal_17448 ), .Q ( signal_17449 ) ) ;
    buf_clk cell_2758 ( .C ( clk ), .D ( signal_17450 ), .Q ( signal_17451 ) ) ;
    buf_clk cell_2760 ( .C ( clk ), .D ( signal_17452 ), .Q ( signal_17453 ) ) ;
    buf_clk cell_2762 ( .C ( clk ), .D ( signal_17454 ), .Q ( signal_17455 ) ) ;
    buf_clk cell_2764 ( .C ( clk ), .D ( signal_17456 ), .Q ( signal_17457 ) ) ;
    buf_clk cell_2766 ( .C ( clk ), .D ( signal_17458 ), .Q ( signal_17459 ) ) ;
    buf_clk cell_2768 ( .C ( clk ), .D ( signal_17460 ), .Q ( signal_17461 ) ) ;
    buf_clk cell_2770 ( .C ( clk ), .D ( signal_17462 ), .Q ( signal_17463 ) ) ;
    buf_clk cell_2772 ( .C ( clk ), .D ( signal_17464 ), .Q ( signal_17465 ) ) ;
    buf_clk cell_2774 ( .C ( clk ), .D ( signal_17466 ), .Q ( signal_17467 ) ) ;
    buf_clk cell_2776 ( .C ( clk ), .D ( signal_17468 ), .Q ( signal_17469 ) ) ;
    buf_clk cell_2778 ( .C ( clk ), .D ( signal_17470 ), .Q ( signal_17471 ) ) ;
    buf_clk cell_2780 ( .C ( clk ), .D ( signal_17472 ), .Q ( signal_17473 ) ) ;
    buf_clk cell_2782 ( .C ( clk ), .D ( signal_17474 ), .Q ( signal_17475 ) ) ;
    buf_clk cell_2784 ( .C ( clk ), .D ( signal_17476 ), .Q ( signal_17477 ) ) ;
    buf_clk cell_2786 ( .C ( clk ), .D ( signal_17478 ), .Q ( signal_17479 ) ) ;
    buf_clk cell_2788 ( .C ( clk ), .D ( signal_17480 ), .Q ( signal_17481 ) ) ;
    buf_clk cell_2790 ( .C ( clk ), .D ( signal_17482 ), .Q ( signal_17483 ) ) ;
    buf_clk cell_2792 ( .C ( clk ), .D ( signal_17484 ), .Q ( signal_17485 ) ) ;
    buf_clk cell_2794 ( .C ( clk ), .D ( signal_17486 ), .Q ( signal_17487 ) ) ;
    buf_clk cell_2796 ( .C ( clk ), .D ( signal_17488 ), .Q ( signal_17489 ) ) ;
    buf_clk cell_2798 ( .C ( clk ), .D ( signal_17490 ), .Q ( signal_17491 ) ) ;
    buf_clk cell_2800 ( .C ( clk ), .D ( signal_17492 ), .Q ( signal_17493 ) ) ;
    buf_clk cell_2802 ( .C ( clk ), .D ( signal_17494 ), .Q ( signal_17495 ) ) ;
    buf_clk cell_2804 ( .C ( clk ), .D ( signal_17496 ), .Q ( signal_17497 ) ) ;
    buf_clk cell_2806 ( .C ( clk ), .D ( signal_17498 ), .Q ( signal_17499 ) ) ;
    buf_clk cell_2808 ( .C ( clk ), .D ( signal_17500 ), .Q ( signal_17501 ) ) ;
    buf_clk cell_2810 ( .C ( clk ), .D ( signal_17502 ), .Q ( signal_17503 ) ) ;
    buf_clk cell_2812 ( .C ( clk ), .D ( signal_17504 ), .Q ( signal_17505 ) ) ;
    buf_clk cell_2814 ( .C ( clk ), .D ( signal_17506 ), .Q ( signal_17507 ) ) ;
    buf_clk cell_2816 ( .C ( clk ), .D ( signal_17508 ), .Q ( signal_17509 ) ) ;
    buf_clk cell_2818 ( .C ( clk ), .D ( signal_17510 ), .Q ( signal_17511 ) ) ;
    buf_clk cell_2820 ( .C ( clk ), .D ( signal_17512 ), .Q ( signal_17513 ) ) ;
    buf_clk cell_2822 ( .C ( clk ), .D ( signal_17514 ), .Q ( signal_17515 ) ) ;
    buf_clk cell_2824 ( .C ( clk ), .D ( signal_17516 ), .Q ( signal_17517 ) ) ;
    buf_clk cell_2826 ( .C ( clk ), .D ( signal_17518 ), .Q ( signal_17519 ) ) ;
    buf_clk cell_2828 ( .C ( clk ), .D ( signal_17520 ), .Q ( signal_17521 ) ) ;
    buf_clk cell_2830 ( .C ( clk ), .D ( signal_17522 ), .Q ( signal_17523 ) ) ;
    buf_clk cell_2832 ( .C ( clk ), .D ( signal_17524 ), .Q ( signal_17525 ) ) ;
    buf_clk cell_2834 ( .C ( clk ), .D ( signal_17526 ), .Q ( signal_17527 ) ) ;
    buf_clk cell_2836 ( .C ( clk ), .D ( signal_17528 ), .Q ( signal_17529 ) ) ;
    buf_clk cell_2838 ( .C ( clk ), .D ( signal_17530 ), .Q ( signal_17531 ) ) ;
    buf_clk cell_2840 ( .C ( clk ), .D ( signal_17532 ), .Q ( signal_17533 ) ) ;
    buf_clk cell_2842 ( .C ( clk ), .D ( signal_17534 ), .Q ( signal_17535 ) ) ;
    buf_clk cell_2844 ( .C ( clk ), .D ( signal_17536 ), .Q ( signal_17537 ) ) ;
    buf_clk cell_2846 ( .C ( clk ), .D ( signal_17538 ), .Q ( signal_17539 ) ) ;
    buf_clk cell_2848 ( .C ( clk ), .D ( signal_17540 ), .Q ( signal_17541 ) ) ;
    buf_clk cell_2850 ( .C ( clk ), .D ( signal_17542 ), .Q ( signal_17543 ) ) ;
    buf_clk cell_2852 ( .C ( clk ), .D ( signal_17544 ), .Q ( signal_17545 ) ) ;
    buf_clk cell_2854 ( .C ( clk ), .D ( signal_17546 ), .Q ( signal_17547 ) ) ;
    buf_clk cell_2856 ( .C ( clk ), .D ( signal_17548 ), .Q ( signal_17549 ) ) ;
    buf_clk cell_2858 ( .C ( clk ), .D ( signal_17550 ), .Q ( signal_17551 ) ) ;
    buf_clk cell_2860 ( .C ( clk ), .D ( signal_17552 ), .Q ( signal_17553 ) ) ;
    buf_clk cell_2862 ( .C ( clk ), .D ( signal_17554 ), .Q ( signal_17555 ) ) ;
    buf_clk cell_2864 ( .C ( clk ), .D ( signal_17556 ), .Q ( signal_17557 ) ) ;
    buf_clk cell_2866 ( .C ( clk ), .D ( signal_17558 ), .Q ( signal_17559 ) ) ;
    buf_clk cell_2868 ( .C ( clk ), .D ( signal_17560 ), .Q ( signal_17561 ) ) ;
    buf_clk cell_2870 ( .C ( clk ), .D ( signal_17562 ), .Q ( signal_17563 ) ) ;
    buf_clk cell_2872 ( .C ( clk ), .D ( signal_17564 ), .Q ( signal_17565 ) ) ;
    buf_clk cell_2874 ( .C ( clk ), .D ( signal_17566 ), .Q ( signal_17567 ) ) ;
    buf_clk cell_2878 ( .C ( clk ), .D ( signal_17570 ), .Q ( signal_17571 ) ) ;
    buf_clk cell_2882 ( .C ( clk ), .D ( signal_17574 ), .Q ( signal_17575 ) ) ;
    buf_clk cell_2886 ( .C ( clk ), .D ( signal_17578 ), .Q ( signal_17579 ) ) ;
    buf_clk cell_2890 ( .C ( clk ), .D ( signal_17582 ), .Q ( signal_17583 ) ) ;
    buf_clk cell_2894 ( .C ( clk ), .D ( signal_17586 ), .Q ( signal_17587 ) ) ;
    buf_clk cell_2896 ( .C ( clk ), .D ( signal_17588 ), .Q ( signal_17589 ) ) ;
    buf_clk cell_2898 ( .C ( clk ), .D ( signal_17590 ), .Q ( signal_17591 ) ) ;
    buf_clk cell_2900 ( .C ( clk ), .D ( signal_17592 ), .Q ( signal_17593 ) ) ;
    buf_clk cell_2902 ( .C ( clk ), .D ( signal_17594 ), .Q ( signal_17595 ) ) ;
    buf_clk cell_2904 ( .C ( clk ), .D ( signal_17596 ), .Q ( signal_17597 ) ) ;
    buf_clk cell_2906 ( .C ( clk ), .D ( signal_17598 ), .Q ( signal_17599 ) ) ;
    buf_clk cell_2908 ( .C ( clk ), .D ( signal_17600 ), .Q ( signal_17601 ) ) ;
    buf_clk cell_2910 ( .C ( clk ), .D ( signal_17602 ), .Q ( signal_17603 ) ) ;
    buf_clk cell_2912 ( .C ( clk ), .D ( signal_17604 ), .Q ( signal_17605 ) ) ;
    buf_clk cell_2914 ( .C ( clk ), .D ( signal_17606 ), .Q ( signal_17607 ) ) ;
    buf_clk cell_2916 ( .C ( clk ), .D ( signal_17608 ), .Q ( signal_17609 ) ) ;
    buf_clk cell_2918 ( .C ( clk ), .D ( signal_17610 ), .Q ( signal_17611 ) ) ;
    buf_clk cell_2920 ( .C ( clk ), .D ( signal_17612 ), .Q ( signal_17613 ) ) ;
    buf_clk cell_2922 ( .C ( clk ), .D ( signal_17614 ), .Q ( signal_17615 ) ) ;
    buf_clk cell_2924 ( .C ( clk ), .D ( signal_17616 ), .Q ( signal_17617 ) ) ;
    buf_clk cell_2926 ( .C ( clk ), .D ( signal_17618 ), .Q ( signal_17619 ) ) ;
    buf_clk cell_2928 ( .C ( clk ), .D ( signal_17620 ), .Q ( signal_17621 ) ) ;
    buf_clk cell_2930 ( .C ( clk ), .D ( signal_17622 ), .Q ( signal_17623 ) ) ;
    buf_clk cell_2932 ( .C ( clk ), .D ( signal_17624 ), .Q ( signal_17625 ) ) ;
    buf_clk cell_2934 ( .C ( clk ), .D ( signal_17626 ), .Q ( signal_17627 ) ) ;
    buf_clk cell_2936 ( .C ( clk ), .D ( signal_17628 ), .Q ( signal_17629 ) ) ;
    buf_clk cell_2938 ( .C ( clk ), .D ( signal_17630 ), .Q ( signal_17631 ) ) ;
    buf_clk cell_2940 ( .C ( clk ), .D ( signal_17632 ), .Q ( signal_17633 ) ) ;
    buf_clk cell_2942 ( .C ( clk ), .D ( signal_17634 ), .Q ( signal_17635 ) ) ;
    buf_clk cell_2944 ( .C ( clk ), .D ( signal_17636 ), .Q ( signal_17637 ) ) ;
    buf_clk cell_2946 ( .C ( clk ), .D ( signal_17638 ), .Q ( signal_17639 ) ) ;
    buf_clk cell_2948 ( .C ( clk ), .D ( signal_17640 ), .Q ( signal_17641 ) ) ;
    buf_clk cell_2950 ( .C ( clk ), .D ( signal_17642 ), .Q ( signal_17643 ) ) ;
    buf_clk cell_2952 ( .C ( clk ), .D ( signal_17644 ), .Q ( signal_17645 ) ) ;
    buf_clk cell_2954 ( .C ( clk ), .D ( signal_17646 ), .Q ( signal_17647 ) ) ;
    buf_clk cell_2956 ( .C ( clk ), .D ( signal_17648 ), .Q ( signal_17649 ) ) ;
    buf_clk cell_2958 ( .C ( clk ), .D ( signal_17650 ), .Q ( signal_17651 ) ) ;
    buf_clk cell_2960 ( .C ( clk ), .D ( signal_17652 ), .Q ( signal_17653 ) ) ;
    buf_clk cell_2962 ( .C ( clk ), .D ( signal_17654 ), .Q ( signal_17655 ) ) ;
    buf_clk cell_2964 ( .C ( clk ), .D ( signal_17656 ), .Q ( signal_17657 ) ) ;
    buf_clk cell_2966 ( .C ( clk ), .D ( signal_17658 ), .Q ( signal_17659 ) ) ;
    buf_clk cell_2968 ( .C ( clk ), .D ( signal_17660 ), .Q ( signal_17661 ) ) ;
    buf_clk cell_2970 ( .C ( clk ), .D ( signal_17662 ), .Q ( signal_17663 ) ) ;
    buf_clk cell_2972 ( .C ( clk ), .D ( signal_17664 ), .Q ( signal_17665 ) ) ;
    buf_clk cell_2974 ( .C ( clk ), .D ( signal_17666 ), .Q ( signal_17667 ) ) ;
    buf_clk cell_2976 ( .C ( clk ), .D ( signal_17668 ), .Q ( signal_17669 ) ) ;
    buf_clk cell_2978 ( .C ( clk ), .D ( signal_17670 ), .Q ( signal_17671 ) ) ;
    buf_clk cell_2980 ( .C ( clk ), .D ( signal_17672 ), .Q ( signal_17673 ) ) ;
    buf_clk cell_2982 ( .C ( clk ), .D ( signal_17674 ), .Q ( signal_17675 ) ) ;
    buf_clk cell_2984 ( .C ( clk ), .D ( signal_17676 ), .Q ( signal_17677 ) ) ;
    buf_clk cell_2986 ( .C ( clk ), .D ( signal_17678 ), .Q ( signal_17679 ) ) ;
    buf_clk cell_2988 ( .C ( clk ), .D ( signal_17680 ), .Q ( signal_17681 ) ) ;
    buf_clk cell_2990 ( .C ( clk ), .D ( signal_17682 ), .Q ( signal_17683 ) ) ;
    buf_clk cell_2992 ( .C ( clk ), .D ( signal_17684 ), .Q ( signal_17685 ) ) ;
    buf_clk cell_2994 ( .C ( clk ), .D ( signal_17686 ), .Q ( signal_17687 ) ) ;
    buf_clk cell_2996 ( .C ( clk ), .D ( signal_17688 ), .Q ( signal_17689 ) ) ;
    buf_clk cell_2998 ( .C ( clk ), .D ( signal_17690 ), .Q ( signal_17691 ) ) ;
    buf_clk cell_3000 ( .C ( clk ), .D ( signal_17692 ), .Q ( signal_17693 ) ) ;
    buf_clk cell_3002 ( .C ( clk ), .D ( signal_17694 ), .Q ( signal_17695 ) ) ;
    buf_clk cell_3004 ( .C ( clk ), .D ( signal_17696 ), .Q ( signal_17697 ) ) ;
    buf_clk cell_3006 ( .C ( clk ), .D ( signal_17698 ), .Q ( signal_17699 ) ) ;
    buf_clk cell_3008 ( .C ( clk ), .D ( signal_17700 ), .Q ( signal_17701 ) ) ;
    buf_clk cell_3010 ( .C ( clk ), .D ( signal_17702 ), .Q ( signal_17703 ) ) ;
    buf_clk cell_3012 ( .C ( clk ), .D ( signal_17704 ), .Q ( signal_17705 ) ) ;
    buf_clk cell_3014 ( .C ( clk ), .D ( signal_17706 ), .Q ( signal_17707 ) ) ;
    buf_clk cell_3016 ( .C ( clk ), .D ( signal_17708 ), .Q ( signal_17709 ) ) ;
    buf_clk cell_3018 ( .C ( clk ), .D ( signal_17710 ), .Q ( signal_17711 ) ) ;
    buf_clk cell_3020 ( .C ( clk ), .D ( signal_17712 ), .Q ( signal_17713 ) ) ;
    buf_clk cell_3022 ( .C ( clk ), .D ( signal_17714 ), .Q ( signal_17715 ) ) ;
    buf_clk cell_3024 ( .C ( clk ), .D ( signal_17716 ), .Q ( signal_17717 ) ) ;
    buf_clk cell_3026 ( .C ( clk ), .D ( signal_17718 ), .Q ( signal_17719 ) ) ;
    buf_clk cell_3028 ( .C ( clk ), .D ( signal_17720 ), .Q ( signal_17721 ) ) ;
    buf_clk cell_3030 ( .C ( clk ), .D ( signal_17722 ), .Q ( signal_17723 ) ) ;
    buf_clk cell_3032 ( .C ( clk ), .D ( signal_17724 ), .Q ( signal_17725 ) ) ;
    buf_clk cell_3034 ( .C ( clk ), .D ( signal_17726 ), .Q ( signal_17727 ) ) ;
    buf_clk cell_3036 ( .C ( clk ), .D ( signal_17728 ), .Q ( signal_17729 ) ) ;
    buf_clk cell_3038 ( .C ( clk ), .D ( signal_17730 ), .Q ( signal_17731 ) ) ;
    buf_clk cell_3040 ( .C ( clk ), .D ( signal_17732 ), .Q ( signal_17733 ) ) ;
    buf_clk cell_3042 ( .C ( clk ), .D ( signal_17734 ), .Q ( signal_17735 ) ) ;
    buf_clk cell_3044 ( .C ( clk ), .D ( signal_17736 ), .Q ( signal_17737 ) ) ;
    buf_clk cell_3046 ( .C ( clk ), .D ( signal_17738 ), .Q ( signal_17739 ) ) ;
    buf_clk cell_3048 ( .C ( clk ), .D ( signal_17740 ), .Q ( signal_17741 ) ) ;
    buf_clk cell_3050 ( .C ( clk ), .D ( signal_17742 ), .Q ( signal_17743 ) ) ;
    buf_clk cell_3052 ( .C ( clk ), .D ( signal_17744 ), .Q ( signal_17745 ) ) ;
    buf_clk cell_3054 ( .C ( clk ), .D ( signal_17746 ), .Q ( signal_17747 ) ) ;
    buf_clk cell_3056 ( .C ( clk ), .D ( signal_17748 ), .Q ( signal_17749 ) ) ;
    buf_clk cell_3058 ( .C ( clk ), .D ( signal_17750 ), .Q ( signal_17751 ) ) ;
    buf_clk cell_3060 ( .C ( clk ), .D ( signal_17752 ), .Q ( signal_17753 ) ) ;
    buf_clk cell_3062 ( .C ( clk ), .D ( signal_17754 ), .Q ( signal_17755 ) ) ;
    buf_clk cell_3064 ( .C ( clk ), .D ( signal_17756 ), .Q ( signal_17757 ) ) ;
    buf_clk cell_3066 ( .C ( clk ), .D ( signal_17758 ), .Q ( signal_17759 ) ) ;
    buf_clk cell_3068 ( .C ( clk ), .D ( signal_17760 ), .Q ( signal_17761 ) ) ;
    buf_clk cell_3070 ( .C ( clk ), .D ( signal_17762 ), .Q ( signal_17763 ) ) ;
    buf_clk cell_3072 ( .C ( clk ), .D ( signal_17764 ), .Q ( signal_17765 ) ) ;
    buf_clk cell_3074 ( .C ( clk ), .D ( signal_17766 ), .Q ( signal_17767 ) ) ;
    buf_clk cell_3076 ( .C ( clk ), .D ( signal_17768 ), .Q ( signal_17769 ) ) ;
    buf_clk cell_3078 ( .C ( clk ), .D ( signal_17770 ), .Q ( signal_17771 ) ) ;
    buf_clk cell_3080 ( .C ( clk ), .D ( signal_17772 ), .Q ( signal_17773 ) ) ;
    buf_clk cell_3082 ( .C ( clk ), .D ( signal_17774 ), .Q ( signal_17775 ) ) ;
    buf_clk cell_3084 ( .C ( clk ), .D ( signal_17776 ), .Q ( signal_17777 ) ) ;
    buf_clk cell_3086 ( .C ( clk ), .D ( signal_17778 ), .Q ( signal_17779 ) ) ;
    buf_clk cell_3088 ( .C ( clk ), .D ( signal_17780 ), .Q ( signal_17781 ) ) ;
    buf_clk cell_3090 ( .C ( clk ), .D ( signal_17782 ), .Q ( signal_17783 ) ) ;
    buf_clk cell_3092 ( .C ( clk ), .D ( signal_17784 ), .Q ( signal_17785 ) ) ;
    buf_clk cell_3094 ( .C ( clk ), .D ( signal_17786 ), .Q ( signal_17787 ) ) ;
    buf_clk cell_3096 ( .C ( clk ), .D ( signal_17788 ), .Q ( signal_17789 ) ) ;
    buf_clk cell_3098 ( .C ( clk ), .D ( signal_17790 ), .Q ( signal_17791 ) ) ;
    buf_clk cell_3100 ( .C ( clk ), .D ( signal_17792 ), .Q ( signal_17793 ) ) ;
    buf_clk cell_3102 ( .C ( clk ), .D ( signal_17794 ), .Q ( signal_17795 ) ) ;
    buf_clk cell_3104 ( .C ( clk ), .D ( signal_17796 ), .Q ( signal_17797 ) ) ;
    buf_clk cell_3106 ( .C ( clk ), .D ( signal_17798 ), .Q ( signal_17799 ) ) ;
    buf_clk cell_3108 ( .C ( clk ), .D ( signal_17800 ), .Q ( signal_17801 ) ) ;
    buf_clk cell_3110 ( .C ( clk ), .D ( signal_17802 ), .Q ( signal_17803 ) ) ;
    buf_clk cell_3112 ( .C ( clk ), .D ( signal_17804 ), .Q ( signal_17805 ) ) ;
    buf_clk cell_3114 ( .C ( clk ), .D ( signal_17806 ), .Q ( signal_17807 ) ) ;
    buf_clk cell_3228 ( .C ( clk ), .D ( signal_17920 ), .Q ( signal_17921 ) ) ;
    buf_clk cell_3234 ( .C ( clk ), .D ( signal_17926 ), .Q ( signal_17927 ) ) ;
    buf_clk cell_3240 ( .C ( clk ), .D ( signal_17932 ), .Q ( signal_17933 ) ) ;
    buf_clk cell_3246 ( .C ( clk ), .D ( signal_17938 ), .Q ( signal_17939 ) ) ;
    buf_clk cell_3252 ( .C ( clk ), .D ( signal_17944 ), .Q ( signal_17945 ) ) ;
    buf_clk cell_3456 ( .C ( clk ), .D ( signal_18148 ), .Q ( signal_18149 ) ) ;
    buf_clk cell_3460 ( .C ( clk ), .D ( signal_18152 ), .Q ( signal_18153 ) ) ;
    buf_clk cell_3464 ( .C ( clk ), .D ( signal_18156 ), .Q ( signal_18157 ) ) ;
    buf_clk cell_3468 ( .C ( clk ), .D ( signal_18160 ), .Q ( signal_18161 ) ) ;
    buf_clk cell_3472 ( .C ( clk ), .D ( signal_18164 ), .Q ( signal_18165 ) ) ;
    buf_clk cell_3496 ( .C ( clk ), .D ( signal_18188 ), .Q ( signal_18189 ) ) ;
    buf_clk cell_3500 ( .C ( clk ), .D ( signal_18192 ), .Q ( signal_18193 ) ) ;
    buf_clk cell_3504 ( .C ( clk ), .D ( signal_18196 ), .Q ( signal_18197 ) ) ;
    buf_clk cell_3508 ( .C ( clk ), .D ( signal_18200 ), .Q ( signal_18201 ) ) ;
    buf_clk cell_3512 ( .C ( clk ), .D ( signal_18204 ), .Q ( signal_18205 ) ) ;
    buf_clk cell_3626 ( .C ( clk ), .D ( signal_18318 ), .Q ( signal_18319 ) ) ;
    buf_clk cell_3630 ( .C ( clk ), .D ( signal_18322 ), .Q ( signal_18323 ) ) ;
    buf_clk cell_3634 ( .C ( clk ), .D ( signal_18326 ), .Q ( signal_18327 ) ) ;
    buf_clk cell_3638 ( .C ( clk ), .D ( signal_18330 ), .Q ( signal_18331 ) ) ;
    buf_clk cell_3642 ( .C ( clk ), .D ( signal_18334 ), .Q ( signal_18335 ) ) ;
    buf_clk cell_3656 ( .C ( clk ), .D ( signal_18348 ), .Q ( signal_18349 ) ) ;
    buf_clk cell_3660 ( .C ( clk ), .D ( signal_18352 ), .Q ( signal_18353 ) ) ;
    buf_clk cell_3664 ( .C ( clk ), .D ( signal_18356 ), .Q ( signal_18357 ) ) ;
    buf_clk cell_3668 ( .C ( clk ), .D ( signal_18360 ), .Q ( signal_18361 ) ) ;
    buf_clk cell_3672 ( .C ( clk ), .D ( signal_18364 ), .Q ( signal_18365 ) ) ;
    buf_clk cell_3708 ( .C ( clk ), .D ( signal_18400 ), .Q ( signal_18401 ) ) ;
    buf_clk cell_3714 ( .C ( clk ), .D ( signal_18406 ), .Q ( signal_18407 ) ) ;
    buf_clk cell_3720 ( .C ( clk ), .D ( signal_18412 ), .Q ( signal_18413 ) ) ;
    buf_clk cell_3726 ( .C ( clk ), .D ( signal_18418 ), .Q ( signal_18419 ) ) ;
    buf_clk cell_3732 ( .C ( clk ), .D ( signal_18424 ), .Q ( signal_18425 ) ) ;
    buf_clk cell_3776 ( .C ( clk ), .D ( signal_18468 ), .Q ( signal_18469 ) ) ;
    buf_clk cell_3780 ( .C ( clk ), .D ( signal_18472 ), .Q ( signal_18473 ) ) ;
    buf_clk cell_3784 ( .C ( clk ), .D ( signal_18476 ), .Q ( signal_18477 ) ) ;
    buf_clk cell_3788 ( .C ( clk ), .D ( signal_18480 ), .Q ( signal_18481 ) ) ;
    buf_clk cell_3792 ( .C ( clk ), .D ( signal_18484 ), .Q ( signal_18485 ) ) ;
    buf_clk cell_3886 ( .C ( clk ), .D ( signal_18578 ), .Q ( signal_18579 ) ) ;
    buf_clk cell_3890 ( .C ( clk ), .D ( signal_18582 ), .Q ( signal_18583 ) ) ;
    buf_clk cell_3894 ( .C ( clk ), .D ( signal_18586 ), .Q ( signal_18587 ) ) ;
    buf_clk cell_3898 ( .C ( clk ), .D ( signal_18590 ), .Q ( signal_18591 ) ) ;
    buf_clk cell_3902 ( .C ( clk ), .D ( signal_18594 ), .Q ( signal_18595 ) ) ;
    buf_clk cell_4078 ( .C ( clk ), .D ( signal_18770 ), .Q ( signal_18771 ) ) ;
    buf_clk cell_4086 ( .C ( clk ), .D ( signal_18778 ), .Q ( signal_18779 ) ) ;
    buf_clk cell_4094 ( .C ( clk ), .D ( signal_18786 ), .Q ( signal_18787 ) ) ;
    buf_clk cell_4102 ( .C ( clk ), .D ( signal_18794 ), .Q ( signal_18795 ) ) ;
    buf_clk cell_4110 ( .C ( clk ), .D ( signal_18802 ), .Q ( signal_18803 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_3115 ( .C ( clk ), .D ( signal_1293 ), .Q ( signal_17808 ) ) ;
    buf_clk cell_3117 ( .C ( clk ), .D ( signal_3828 ), .Q ( signal_17810 ) ) ;
    buf_clk cell_3119 ( .C ( clk ), .D ( signal_3829 ), .Q ( signal_17812 ) ) ;
    buf_clk cell_3121 ( .C ( clk ), .D ( signal_3830 ), .Q ( signal_17814 ) ) ;
    buf_clk cell_3123 ( .C ( clk ), .D ( signal_3831 ), .Q ( signal_17816 ) ) ;
    buf_clk cell_3125 ( .C ( clk ), .D ( signal_17549 ), .Q ( signal_17818 ) ) ;
    buf_clk cell_3127 ( .C ( clk ), .D ( signal_17551 ), .Q ( signal_17820 ) ) ;
    buf_clk cell_3129 ( .C ( clk ), .D ( signal_17553 ), .Q ( signal_17822 ) ) ;
    buf_clk cell_3131 ( .C ( clk ), .D ( signal_17555 ), .Q ( signal_17824 ) ) ;
    buf_clk cell_3133 ( .C ( clk ), .D ( signal_17557 ), .Q ( signal_17826 ) ) ;
    buf_clk cell_3135 ( .C ( clk ), .D ( signal_1328 ), .Q ( signal_17828 ) ) ;
    buf_clk cell_3137 ( .C ( clk ), .D ( signal_3968 ), .Q ( signal_17830 ) ) ;
    buf_clk cell_3139 ( .C ( clk ), .D ( signal_3969 ), .Q ( signal_17832 ) ) ;
    buf_clk cell_3141 ( .C ( clk ), .D ( signal_3970 ), .Q ( signal_17834 ) ) ;
    buf_clk cell_3143 ( .C ( clk ), .D ( signal_3971 ), .Q ( signal_17836 ) ) ;
    buf_clk cell_3145 ( .C ( clk ), .D ( signal_1342 ), .Q ( signal_17838 ) ) ;
    buf_clk cell_3147 ( .C ( clk ), .D ( signal_4024 ), .Q ( signal_17840 ) ) ;
    buf_clk cell_3149 ( .C ( clk ), .D ( signal_4025 ), .Q ( signal_17842 ) ) ;
    buf_clk cell_3151 ( .C ( clk ), .D ( signal_4026 ), .Q ( signal_17844 ) ) ;
    buf_clk cell_3153 ( .C ( clk ), .D ( signal_4027 ), .Q ( signal_17846 ) ) ;
    buf_clk cell_3155 ( .C ( clk ), .D ( signal_1282 ), .Q ( signal_17848 ) ) ;
    buf_clk cell_3157 ( .C ( clk ), .D ( signal_3784 ), .Q ( signal_17850 ) ) ;
    buf_clk cell_3159 ( .C ( clk ), .D ( signal_3785 ), .Q ( signal_17852 ) ) ;
    buf_clk cell_3161 ( .C ( clk ), .D ( signal_3786 ), .Q ( signal_17854 ) ) ;
    buf_clk cell_3163 ( .C ( clk ), .D ( signal_3787 ), .Q ( signal_17856 ) ) ;
    buf_clk cell_3165 ( .C ( clk ), .D ( signal_1291 ), .Q ( signal_17858 ) ) ;
    buf_clk cell_3167 ( .C ( clk ), .D ( signal_3820 ), .Q ( signal_17860 ) ) ;
    buf_clk cell_3169 ( .C ( clk ), .D ( signal_3821 ), .Q ( signal_17862 ) ) ;
    buf_clk cell_3171 ( .C ( clk ), .D ( signal_3822 ), .Q ( signal_17864 ) ) ;
    buf_clk cell_3173 ( .C ( clk ), .D ( signal_3823 ), .Q ( signal_17866 ) ) ;
    buf_clk cell_3175 ( .C ( clk ), .D ( signal_17299 ), .Q ( signal_17868 ) ) ;
    buf_clk cell_3177 ( .C ( clk ), .D ( signal_17301 ), .Q ( signal_17870 ) ) ;
    buf_clk cell_3179 ( .C ( clk ), .D ( signal_17303 ), .Q ( signal_17872 ) ) ;
    buf_clk cell_3181 ( .C ( clk ), .D ( signal_17305 ), .Q ( signal_17874 ) ) ;
    buf_clk cell_3183 ( .C ( clk ), .D ( signal_17307 ), .Q ( signal_17876 ) ) ;
    buf_clk cell_3185 ( .C ( clk ), .D ( signal_17379 ), .Q ( signal_17878 ) ) ;
    buf_clk cell_3187 ( .C ( clk ), .D ( signal_17381 ), .Q ( signal_17880 ) ) ;
    buf_clk cell_3189 ( .C ( clk ), .D ( signal_17383 ), .Q ( signal_17882 ) ) ;
    buf_clk cell_3191 ( .C ( clk ), .D ( signal_17385 ), .Q ( signal_17884 ) ) ;
    buf_clk cell_3193 ( .C ( clk ), .D ( signal_17387 ), .Q ( signal_17886 ) ) ;
    buf_clk cell_3195 ( .C ( clk ), .D ( signal_17389 ), .Q ( signal_17888 ) ) ;
    buf_clk cell_3197 ( .C ( clk ), .D ( signal_17391 ), .Q ( signal_17890 ) ) ;
    buf_clk cell_3199 ( .C ( clk ), .D ( signal_17393 ), .Q ( signal_17892 ) ) ;
    buf_clk cell_3201 ( .C ( clk ), .D ( signal_17395 ), .Q ( signal_17894 ) ) ;
    buf_clk cell_3203 ( .C ( clk ), .D ( signal_17397 ), .Q ( signal_17896 ) ) ;
    buf_clk cell_3205 ( .C ( clk ), .D ( signal_17709 ), .Q ( signal_17898 ) ) ;
    buf_clk cell_3207 ( .C ( clk ), .D ( signal_17711 ), .Q ( signal_17900 ) ) ;
    buf_clk cell_3209 ( .C ( clk ), .D ( signal_17713 ), .Q ( signal_17902 ) ) ;
    buf_clk cell_3211 ( .C ( clk ), .D ( signal_17715 ), .Q ( signal_17904 ) ) ;
    buf_clk cell_3213 ( .C ( clk ), .D ( signal_17717 ), .Q ( signal_17906 ) ) ;
    buf_clk cell_3215 ( .C ( clk ), .D ( signal_17479 ), .Q ( signal_17908 ) ) ;
    buf_clk cell_3217 ( .C ( clk ), .D ( signal_17481 ), .Q ( signal_17910 ) ) ;
    buf_clk cell_3219 ( .C ( clk ), .D ( signal_17483 ), .Q ( signal_17912 ) ) ;
    buf_clk cell_3221 ( .C ( clk ), .D ( signal_17485 ), .Q ( signal_17914 ) ) ;
    buf_clk cell_3223 ( .C ( clk ), .D ( signal_17487 ), .Q ( signal_17916 ) ) ;
    buf_clk cell_3229 ( .C ( clk ), .D ( signal_17921 ), .Q ( signal_17922 ) ) ;
    buf_clk cell_3235 ( .C ( clk ), .D ( signal_17927 ), .Q ( signal_17928 ) ) ;
    buf_clk cell_3241 ( .C ( clk ), .D ( signal_17933 ), .Q ( signal_17934 ) ) ;
    buf_clk cell_3247 ( .C ( clk ), .D ( signal_17939 ), .Q ( signal_17940 ) ) ;
    buf_clk cell_3253 ( .C ( clk ), .D ( signal_17945 ), .Q ( signal_17946 ) ) ;
    buf_clk cell_3255 ( .C ( clk ), .D ( signal_17539 ), .Q ( signal_17948 ) ) ;
    buf_clk cell_3257 ( .C ( clk ), .D ( signal_17541 ), .Q ( signal_17950 ) ) ;
    buf_clk cell_3259 ( .C ( clk ), .D ( signal_17543 ), .Q ( signal_17952 ) ) ;
    buf_clk cell_3261 ( .C ( clk ), .D ( signal_17545 ), .Q ( signal_17954 ) ) ;
    buf_clk cell_3263 ( .C ( clk ), .D ( signal_17547 ), .Q ( signal_17956 ) ) ;
    buf_clk cell_3265 ( .C ( clk ), .D ( signal_17739 ), .Q ( signal_17958 ) ) ;
    buf_clk cell_3267 ( .C ( clk ), .D ( signal_17741 ), .Q ( signal_17960 ) ) ;
    buf_clk cell_3269 ( .C ( clk ), .D ( signal_17743 ), .Q ( signal_17962 ) ) ;
    buf_clk cell_3271 ( .C ( clk ), .D ( signal_17745 ), .Q ( signal_17964 ) ) ;
    buf_clk cell_3273 ( .C ( clk ), .D ( signal_17747 ), .Q ( signal_17966 ) ) ;
    buf_clk cell_3275 ( .C ( clk ), .D ( signal_17259 ), .Q ( signal_17968 ) ) ;
    buf_clk cell_3277 ( .C ( clk ), .D ( signal_17261 ), .Q ( signal_17970 ) ) ;
    buf_clk cell_3279 ( .C ( clk ), .D ( signal_17263 ), .Q ( signal_17972 ) ) ;
    buf_clk cell_3281 ( .C ( clk ), .D ( signal_17265 ), .Q ( signal_17974 ) ) ;
    buf_clk cell_3283 ( .C ( clk ), .D ( signal_17267 ), .Q ( signal_17976 ) ) ;
    buf_clk cell_3285 ( .C ( clk ), .D ( signal_17369 ), .Q ( signal_17978 ) ) ;
    buf_clk cell_3287 ( .C ( clk ), .D ( signal_17371 ), .Q ( signal_17980 ) ) ;
    buf_clk cell_3289 ( .C ( clk ), .D ( signal_17373 ), .Q ( signal_17982 ) ) ;
    buf_clk cell_3291 ( .C ( clk ), .D ( signal_17375 ), .Q ( signal_17984 ) ) ;
    buf_clk cell_3293 ( .C ( clk ), .D ( signal_17377 ), .Q ( signal_17986 ) ) ;
    buf_clk cell_3295 ( .C ( clk ), .D ( signal_1048 ), .Q ( signal_17988 ) ) ;
    buf_clk cell_3297 ( .C ( clk ), .D ( signal_2848 ), .Q ( signal_17990 ) ) ;
    buf_clk cell_3299 ( .C ( clk ), .D ( signal_2849 ), .Q ( signal_17992 ) ) ;
    buf_clk cell_3301 ( .C ( clk ), .D ( signal_2850 ), .Q ( signal_17994 ) ) ;
    buf_clk cell_3303 ( .C ( clk ), .D ( signal_2851 ), .Q ( signal_17996 ) ) ;
    buf_clk cell_3305 ( .C ( clk ), .D ( signal_17339 ), .Q ( signal_17998 ) ) ;
    buf_clk cell_3307 ( .C ( clk ), .D ( signal_17341 ), .Q ( signal_18000 ) ) ;
    buf_clk cell_3309 ( .C ( clk ), .D ( signal_17343 ), .Q ( signal_18002 ) ) ;
    buf_clk cell_3311 ( .C ( clk ), .D ( signal_17345 ), .Q ( signal_18004 ) ) ;
    buf_clk cell_3313 ( .C ( clk ), .D ( signal_17347 ), .Q ( signal_18006 ) ) ;
    buf_clk cell_3315 ( .C ( clk ), .D ( signal_1262 ), .Q ( signal_18008 ) ) ;
    buf_clk cell_3317 ( .C ( clk ), .D ( signal_3704 ), .Q ( signal_18010 ) ) ;
    buf_clk cell_3319 ( .C ( clk ), .D ( signal_3705 ), .Q ( signal_18012 ) ) ;
    buf_clk cell_3321 ( .C ( clk ), .D ( signal_3706 ), .Q ( signal_18014 ) ) ;
    buf_clk cell_3323 ( .C ( clk ), .D ( signal_3707 ), .Q ( signal_18016 ) ) ;
    buf_clk cell_3325 ( .C ( clk ), .D ( signal_1244 ), .Q ( signal_18018 ) ) ;
    buf_clk cell_3327 ( .C ( clk ), .D ( signal_3632 ), .Q ( signal_18020 ) ) ;
    buf_clk cell_3329 ( .C ( clk ), .D ( signal_3633 ), .Q ( signal_18022 ) ) ;
    buf_clk cell_3331 ( .C ( clk ), .D ( signal_3634 ), .Q ( signal_18024 ) ) ;
    buf_clk cell_3333 ( .C ( clk ), .D ( signal_3635 ), .Q ( signal_18026 ) ) ;
    buf_clk cell_3335 ( .C ( clk ), .D ( signal_1275 ), .Q ( signal_18028 ) ) ;
    buf_clk cell_3337 ( .C ( clk ), .D ( signal_3756 ), .Q ( signal_18030 ) ) ;
    buf_clk cell_3339 ( .C ( clk ), .D ( signal_3757 ), .Q ( signal_18032 ) ) ;
    buf_clk cell_3341 ( .C ( clk ), .D ( signal_3758 ), .Q ( signal_18034 ) ) ;
    buf_clk cell_3343 ( .C ( clk ), .D ( signal_3759 ), .Q ( signal_18036 ) ) ;
    buf_clk cell_3345 ( .C ( clk ), .D ( signal_1255 ), .Q ( signal_18038 ) ) ;
    buf_clk cell_3347 ( .C ( clk ), .D ( signal_3676 ), .Q ( signal_18040 ) ) ;
    buf_clk cell_3349 ( .C ( clk ), .D ( signal_3677 ), .Q ( signal_18042 ) ) ;
    buf_clk cell_3351 ( .C ( clk ), .D ( signal_3678 ), .Q ( signal_18044 ) ) ;
    buf_clk cell_3353 ( .C ( clk ), .D ( signal_3679 ), .Q ( signal_18046 ) ) ;
    buf_clk cell_3355 ( .C ( clk ), .D ( signal_1353 ), .Q ( signal_18048 ) ) ;
    buf_clk cell_3357 ( .C ( clk ), .D ( signal_4068 ), .Q ( signal_18050 ) ) ;
    buf_clk cell_3359 ( .C ( clk ), .D ( signal_4069 ), .Q ( signal_18052 ) ) ;
    buf_clk cell_3361 ( .C ( clk ), .D ( signal_4070 ), .Q ( signal_18054 ) ) ;
    buf_clk cell_3363 ( .C ( clk ), .D ( signal_4071 ), .Q ( signal_18056 ) ) ;
    buf_clk cell_3365 ( .C ( clk ), .D ( signal_1349 ), .Q ( signal_18058 ) ) ;
    buf_clk cell_3367 ( .C ( clk ), .D ( signal_4052 ), .Q ( signal_18060 ) ) ;
    buf_clk cell_3369 ( .C ( clk ), .D ( signal_4053 ), .Q ( signal_18062 ) ) ;
    buf_clk cell_3371 ( .C ( clk ), .D ( signal_4054 ), .Q ( signal_18064 ) ) ;
    buf_clk cell_3373 ( .C ( clk ), .D ( signal_4055 ), .Q ( signal_18066 ) ) ;
    buf_clk cell_3375 ( .C ( clk ), .D ( signal_1232 ), .Q ( signal_18068 ) ) ;
    buf_clk cell_3377 ( .C ( clk ), .D ( signal_3584 ), .Q ( signal_18070 ) ) ;
    buf_clk cell_3379 ( .C ( clk ), .D ( signal_3585 ), .Q ( signal_18072 ) ) ;
    buf_clk cell_3381 ( .C ( clk ), .D ( signal_3586 ), .Q ( signal_18074 ) ) ;
    buf_clk cell_3383 ( .C ( clk ), .D ( signal_3587 ), .Q ( signal_18076 ) ) ;
    buf_clk cell_3385 ( .C ( clk ), .D ( signal_1285 ), .Q ( signal_18078 ) ) ;
    buf_clk cell_3387 ( .C ( clk ), .D ( signal_3796 ), .Q ( signal_18080 ) ) ;
    buf_clk cell_3389 ( .C ( clk ), .D ( signal_3797 ), .Q ( signal_18082 ) ) ;
    buf_clk cell_3391 ( .C ( clk ), .D ( signal_3798 ), .Q ( signal_18084 ) ) ;
    buf_clk cell_3393 ( .C ( clk ), .D ( signal_3799 ), .Q ( signal_18086 ) ) ;
    buf_clk cell_3395 ( .C ( clk ), .D ( signal_1245 ), .Q ( signal_18088 ) ) ;
    buf_clk cell_3397 ( .C ( clk ), .D ( signal_3636 ), .Q ( signal_18090 ) ) ;
    buf_clk cell_3399 ( .C ( clk ), .D ( signal_3637 ), .Q ( signal_18092 ) ) ;
    buf_clk cell_3401 ( .C ( clk ), .D ( signal_3638 ), .Q ( signal_18094 ) ) ;
    buf_clk cell_3403 ( .C ( clk ), .D ( signal_3639 ), .Q ( signal_18096 ) ) ;
    buf_clk cell_3405 ( .C ( clk ), .D ( signal_1246 ), .Q ( signal_18098 ) ) ;
    buf_clk cell_3407 ( .C ( clk ), .D ( signal_3640 ), .Q ( signal_18100 ) ) ;
    buf_clk cell_3409 ( .C ( clk ), .D ( signal_3641 ), .Q ( signal_18102 ) ) ;
    buf_clk cell_3411 ( .C ( clk ), .D ( signal_3642 ), .Q ( signal_18104 ) ) ;
    buf_clk cell_3413 ( .C ( clk ), .D ( signal_3643 ), .Q ( signal_18106 ) ) ;
    buf_clk cell_3415 ( .C ( clk ), .D ( signal_1063 ), .Q ( signal_18108 ) ) ;
    buf_clk cell_3417 ( .C ( clk ), .D ( signal_2908 ), .Q ( signal_18110 ) ) ;
    buf_clk cell_3419 ( .C ( clk ), .D ( signal_2909 ), .Q ( signal_18112 ) ) ;
    buf_clk cell_3421 ( .C ( clk ), .D ( signal_2910 ), .Q ( signal_18114 ) ) ;
    buf_clk cell_3423 ( .C ( clk ), .D ( signal_2911 ), .Q ( signal_18116 ) ) ;
    buf_clk cell_3425 ( .C ( clk ), .D ( signal_1301 ), .Q ( signal_18118 ) ) ;
    buf_clk cell_3427 ( .C ( clk ), .D ( signal_3860 ), .Q ( signal_18120 ) ) ;
    buf_clk cell_3429 ( .C ( clk ), .D ( signal_3861 ), .Q ( signal_18122 ) ) ;
    buf_clk cell_3431 ( .C ( clk ), .D ( signal_3862 ), .Q ( signal_18124 ) ) ;
    buf_clk cell_3433 ( .C ( clk ), .D ( signal_3863 ), .Q ( signal_18126 ) ) ;
    buf_clk cell_3435 ( .C ( clk ), .D ( signal_1249 ), .Q ( signal_18128 ) ) ;
    buf_clk cell_3437 ( .C ( clk ), .D ( signal_3652 ), .Q ( signal_18130 ) ) ;
    buf_clk cell_3439 ( .C ( clk ), .D ( signal_3653 ), .Q ( signal_18132 ) ) ;
    buf_clk cell_3441 ( .C ( clk ), .D ( signal_3654 ), .Q ( signal_18134 ) ) ;
    buf_clk cell_3443 ( .C ( clk ), .D ( signal_3655 ), .Q ( signal_18136 ) ) ;
    buf_clk cell_3445 ( .C ( clk ), .D ( signal_1303 ), .Q ( signal_18138 ) ) ;
    buf_clk cell_3447 ( .C ( clk ), .D ( signal_3868 ), .Q ( signal_18140 ) ) ;
    buf_clk cell_3449 ( .C ( clk ), .D ( signal_3869 ), .Q ( signal_18142 ) ) ;
    buf_clk cell_3451 ( .C ( clk ), .D ( signal_3870 ), .Q ( signal_18144 ) ) ;
    buf_clk cell_3453 ( .C ( clk ), .D ( signal_3871 ), .Q ( signal_18146 ) ) ;
    buf_clk cell_3457 ( .C ( clk ), .D ( signal_18149 ), .Q ( signal_18150 ) ) ;
    buf_clk cell_3461 ( .C ( clk ), .D ( signal_18153 ), .Q ( signal_18154 ) ) ;
    buf_clk cell_3465 ( .C ( clk ), .D ( signal_18157 ), .Q ( signal_18158 ) ) ;
    buf_clk cell_3469 ( .C ( clk ), .D ( signal_18161 ), .Q ( signal_18162 ) ) ;
    buf_clk cell_3473 ( .C ( clk ), .D ( signal_18165 ), .Q ( signal_18166 ) ) ;
    buf_clk cell_3475 ( .C ( clk ), .D ( signal_1253 ), .Q ( signal_18168 ) ) ;
    buf_clk cell_3477 ( .C ( clk ), .D ( signal_3668 ), .Q ( signal_18170 ) ) ;
    buf_clk cell_3479 ( .C ( clk ), .D ( signal_3669 ), .Q ( signal_18172 ) ) ;
    buf_clk cell_3481 ( .C ( clk ), .D ( signal_3670 ), .Q ( signal_18174 ) ) ;
    buf_clk cell_3483 ( .C ( clk ), .D ( signal_3671 ), .Q ( signal_18176 ) ) ;
    buf_clk cell_3485 ( .C ( clk ), .D ( signal_1259 ), .Q ( signal_18178 ) ) ;
    buf_clk cell_3487 ( .C ( clk ), .D ( signal_3692 ), .Q ( signal_18180 ) ) ;
    buf_clk cell_3489 ( .C ( clk ), .D ( signal_3693 ), .Q ( signal_18182 ) ) ;
    buf_clk cell_3491 ( .C ( clk ), .D ( signal_3694 ), .Q ( signal_18184 ) ) ;
    buf_clk cell_3493 ( .C ( clk ), .D ( signal_3695 ), .Q ( signal_18186 ) ) ;
    buf_clk cell_3497 ( .C ( clk ), .D ( signal_18189 ), .Q ( signal_18190 ) ) ;
    buf_clk cell_3501 ( .C ( clk ), .D ( signal_18193 ), .Q ( signal_18194 ) ) ;
    buf_clk cell_3505 ( .C ( clk ), .D ( signal_18197 ), .Q ( signal_18198 ) ) ;
    buf_clk cell_3509 ( .C ( clk ), .D ( signal_18201 ), .Q ( signal_18202 ) ) ;
    buf_clk cell_3513 ( .C ( clk ), .D ( signal_18205 ), .Q ( signal_18206 ) ) ;
    buf_clk cell_3515 ( .C ( clk ), .D ( signal_1339 ), .Q ( signal_18208 ) ) ;
    buf_clk cell_3517 ( .C ( clk ), .D ( signal_4012 ), .Q ( signal_18210 ) ) ;
    buf_clk cell_3519 ( .C ( clk ), .D ( signal_4013 ), .Q ( signal_18212 ) ) ;
    buf_clk cell_3521 ( .C ( clk ), .D ( signal_4014 ), .Q ( signal_18214 ) ) ;
    buf_clk cell_3523 ( .C ( clk ), .D ( signal_4015 ), .Q ( signal_18216 ) ) ;
    buf_clk cell_3525 ( .C ( clk ), .D ( signal_17419 ), .Q ( signal_18218 ) ) ;
    buf_clk cell_3527 ( .C ( clk ), .D ( signal_17421 ), .Q ( signal_18220 ) ) ;
    buf_clk cell_3529 ( .C ( clk ), .D ( signal_17423 ), .Q ( signal_18222 ) ) ;
    buf_clk cell_3531 ( .C ( clk ), .D ( signal_17425 ), .Q ( signal_18224 ) ) ;
    buf_clk cell_3533 ( .C ( clk ), .D ( signal_17427 ), .Q ( signal_18226 ) ) ;
    buf_clk cell_3535 ( .C ( clk ), .D ( signal_1272 ), .Q ( signal_18228 ) ) ;
    buf_clk cell_3537 ( .C ( clk ), .D ( signal_3744 ), .Q ( signal_18230 ) ) ;
    buf_clk cell_3539 ( .C ( clk ), .D ( signal_3745 ), .Q ( signal_18232 ) ) ;
    buf_clk cell_3541 ( .C ( clk ), .D ( signal_3746 ), .Q ( signal_18234 ) ) ;
    buf_clk cell_3543 ( .C ( clk ), .D ( signal_3747 ), .Q ( signal_18236 ) ) ;
    buf_clk cell_3545 ( .C ( clk ), .D ( signal_1062 ), .Q ( signal_18238 ) ) ;
    buf_clk cell_3547 ( .C ( clk ), .D ( signal_2904 ), .Q ( signal_18240 ) ) ;
    buf_clk cell_3549 ( .C ( clk ), .D ( signal_2905 ), .Q ( signal_18242 ) ) ;
    buf_clk cell_3551 ( .C ( clk ), .D ( signal_2906 ), .Q ( signal_18244 ) ) ;
    buf_clk cell_3553 ( .C ( clk ), .D ( signal_2907 ), .Q ( signal_18246 ) ) ;
    buf_clk cell_3555 ( .C ( clk ), .D ( signal_1345 ), .Q ( signal_18248 ) ) ;
    buf_clk cell_3557 ( .C ( clk ), .D ( signal_4036 ), .Q ( signal_18250 ) ) ;
    buf_clk cell_3559 ( .C ( clk ), .D ( signal_4037 ), .Q ( signal_18252 ) ) ;
    buf_clk cell_3561 ( .C ( clk ), .D ( signal_4038 ), .Q ( signal_18254 ) ) ;
    buf_clk cell_3563 ( .C ( clk ), .D ( signal_4039 ), .Q ( signal_18256 ) ) ;
    buf_clk cell_3565 ( .C ( clk ), .D ( signal_1278 ), .Q ( signal_18258 ) ) ;
    buf_clk cell_3567 ( .C ( clk ), .D ( signal_3768 ), .Q ( signal_18260 ) ) ;
    buf_clk cell_3569 ( .C ( clk ), .D ( signal_3769 ), .Q ( signal_18262 ) ) ;
    buf_clk cell_3571 ( .C ( clk ), .D ( signal_3770 ), .Q ( signal_18264 ) ) ;
    buf_clk cell_3573 ( .C ( clk ), .D ( signal_3771 ), .Q ( signal_18266 ) ) ;
    buf_clk cell_3575 ( .C ( clk ), .D ( signal_1238 ), .Q ( signal_18268 ) ) ;
    buf_clk cell_3577 ( .C ( clk ), .D ( signal_3608 ), .Q ( signal_18270 ) ) ;
    buf_clk cell_3579 ( .C ( clk ), .D ( signal_3609 ), .Q ( signal_18272 ) ) ;
    buf_clk cell_3581 ( .C ( clk ), .D ( signal_3610 ), .Q ( signal_18274 ) ) ;
    buf_clk cell_3583 ( .C ( clk ), .D ( signal_3611 ), .Q ( signal_18276 ) ) ;
    buf_clk cell_3585 ( .C ( clk ), .D ( signal_1279 ), .Q ( signal_18278 ) ) ;
    buf_clk cell_3587 ( .C ( clk ), .D ( signal_3772 ), .Q ( signal_18280 ) ) ;
    buf_clk cell_3589 ( .C ( clk ), .D ( signal_3773 ), .Q ( signal_18282 ) ) ;
    buf_clk cell_3591 ( .C ( clk ), .D ( signal_3774 ), .Q ( signal_18284 ) ) ;
    buf_clk cell_3593 ( .C ( clk ), .D ( signal_3775 ), .Q ( signal_18286 ) ) ;
    buf_clk cell_3595 ( .C ( clk ), .D ( signal_1233 ), .Q ( signal_18288 ) ) ;
    buf_clk cell_3597 ( .C ( clk ), .D ( signal_3588 ), .Q ( signal_18290 ) ) ;
    buf_clk cell_3599 ( .C ( clk ), .D ( signal_3589 ), .Q ( signal_18292 ) ) ;
    buf_clk cell_3601 ( .C ( clk ), .D ( signal_3590 ), .Q ( signal_18294 ) ) ;
    buf_clk cell_3603 ( .C ( clk ), .D ( signal_3591 ), .Q ( signal_18296 ) ) ;
    buf_clk cell_3605 ( .C ( clk ), .D ( signal_1286 ), .Q ( signal_18298 ) ) ;
    buf_clk cell_3607 ( .C ( clk ), .D ( signal_3800 ), .Q ( signal_18300 ) ) ;
    buf_clk cell_3609 ( .C ( clk ), .D ( signal_3801 ), .Q ( signal_18302 ) ) ;
    buf_clk cell_3611 ( .C ( clk ), .D ( signal_3802 ), .Q ( signal_18304 ) ) ;
    buf_clk cell_3613 ( .C ( clk ), .D ( signal_3803 ), .Q ( signal_18306 ) ) ;
    buf_clk cell_3615 ( .C ( clk ), .D ( signal_1265 ), .Q ( signal_18308 ) ) ;
    buf_clk cell_3617 ( .C ( clk ), .D ( signal_3716 ), .Q ( signal_18310 ) ) ;
    buf_clk cell_3619 ( .C ( clk ), .D ( signal_3717 ), .Q ( signal_18312 ) ) ;
    buf_clk cell_3621 ( .C ( clk ), .D ( signal_3718 ), .Q ( signal_18314 ) ) ;
    buf_clk cell_3623 ( .C ( clk ), .D ( signal_3719 ), .Q ( signal_18316 ) ) ;
    buf_clk cell_3627 ( .C ( clk ), .D ( signal_18319 ), .Q ( signal_18320 ) ) ;
    buf_clk cell_3631 ( .C ( clk ), .D ( signal_18323 ), .Q ( signal_18324 ) ) ;
    buf_clk cell_3635 ( .C ( clk ), .D ( signal_18327 ), .Q ( signal_18328 ) ) ;
    buf_clk cell_3639 ( .C ( clk ), .D ( signal_18331 ), .Q ( signal_18332 ) ) ;
    buf_clk cell_3643 ( .C ( clk ), .D ( signal_18335 ), .Q ( signal_18336 ) ) ;
    buf_clk cell_3645 ( .C ( clk ), .D ( signal_17529 ), .Q ( signal_18338 ) ) ;
    buf_clk cell_3647 ( .C ( clk ), .D ( signal_17531 ), .Q ( signal_18340 ) ) ;
    buf_clk cell_3649 ( .C ( clk ), .D ( signal_17533 ), .Q ( signal_18342 ) ) ;
    buf_clk cell_3651 ( .C ( clk ), .D ( signal_17535 ), .Q ( signal_18344 ) ) ;
    buf_clk cell_3653 ( .C ( clk ), .D ( signal_17537 ), .Q ( signal_18346 ) ) ;
    buf_clk cell_3657 ( .C ( clk ), .D ( signal_18349 ), .Q ( signal_18350 ) ) ;
    buf_clk cell_3661 ( .C ( clk ), .D ( signal_18353 ), .Q ( signal_18354 ) ) ;
    buf_clk cell_3665 ( .C ( clk ), .D ( signal_18357 ), .Q ( signal_18358 ) ) ;
    buf_clk cell_3669 ( .C ( clk ), .D ( signal_18361 ), .Q ( signal_18362 ) ) ;
    buf_clk cell_3673 ( .C ( clk ), .D ( signal_18365 ), .Q ( signal_18366 ) ) ;
    buf_clk cell_3675 ( .C ( clk ), .D ( signal_1333 ), .Q ( signal_18368 ) ) ;
    buf_clk cell_3677 ( .C ( clk ), .D ( signal_3988 ), .Q ( signal_18370 ) ) ;
    buf_clk cell_3679 ( .C ( clk ), .D ( signal_3989 ), .Q ( signal_18372 ) ) ;
    buf_clk cell_3681 ( .C ( clk ), .D ( signal_3990 ), .Q ( signal_18374 ) ) ;
    buf_clk cell_3683 ( .C ( clk ), .D ( signal_3991 ), .Q ( signal_18376 ) ) ;
    buf_clk cell_3685 ( .C ( clk ), .D ( signal_17609 ), .Q ( signal_18378 ) ) ;
    buf_clk cell_3687 ( .C ( clk ), .D ( signal_17611 ), .Q ( signal_18380 ) ) ;
    buf_clk cell_3689 ( .C ( clk ), .D ( signal_17613 ), .Q ( signal_18382 ) ) ;
    buf_clk cell_3691 ( .C ( clk ), .D ( signal_17615 ), .Q ( signal_18384 ) ) ;
    buf_clk cell_3693 ( .C ( clk ), .D ( signal_17617 ), .Q ( signal_18386 ) ) ;
    buf_clk cell_3695 ( .C ( clk ), .D ( signal_17571 ), .Q ( signal_18388 ) ) ;
    buf_clk cell_3697 ( .C ( clk ), .D ( signal_17575 ), .Q ( signal_18390 ) ) ;
    buf_clk cell_3699 ( .C ( clk ), .D ( signal_17579 ), .Q ( signal_18392 ) ) ;
    buf_clk cell_3701 ( .C ( clk ), .D ( signal_17583 ), .Q ( signal_18394 ) ) ;
    buf_clk cell_3703 ( .C ( clk ), .D ( signal_17587 ), .Q ( signal_18396 ) ) ;
    buf_clk cell_3709 ( .C ( clk ), .D ( signal_18401 ), .Q ( signal_18402 ) ) ;
    buf_clk cell_3715 ( .C ( clk ), .D ( signal_18407 ), .Q ( signal_18408 ) ) ;
    buf_clk cell_3721 ( .C ( clk ), .D ( signal_18413 ), .Q ( signal_18414 ) ) ;
    buf_clk cell_3727 ( .C ( clk ), .D ( signal_18419 ), .Q ( signal_18420 ) ) ;
    buf_clk cell_3733 ( .C ( clk ), .D ( signal_18425 ), .Q ( signal_18426 ) ) ;
    buf_clk cell_3735 ( .C ( clk ), .D ( signal_17489 ), .Q ( signal_18428 ) ) ;
    buf_clk cell_3737 ( .C ( clk ), .D ( signal_17491 ), .Q ( signal_18430 ) ) ;
    buf_clk cell_3739 ( .C ( clk ), .D ( signal_17493 ), .Q ( signal_18432 ) ) ;
    buf_clk cell_3741 ( .C ( clk ), .D ( signal_17495 ), .Q ( signal_18434 ) ) ;
    buf_clk cell_3743 ( .C ( clk ), .D ( signal_17497 ), .Q ( signal_18436 ) ) ;
    buf_clk cell_3745 ( .C ( clk ), .D ( signal_17279 ), .Q ( signal_18438 ) ) ;
    buf_clk cell_3747 ( .C ( clk ), .D ( signal_17281 ), .Q ( signal_18440 ) ) ;
    buf_clk cell_3749 ( .C ( clk ), .D ( signal_17283 ), .Q ( signal_18442 ) ) ;
    buf_clk cell_3751 ( .C ( clk ), .D ( signal_17285 ), .Q ( signal_18444 ) ) ;
    buf_clk cell_3753 ( .C ( clk ), .D ( signal_17287 ), .Q ( signal_18446 ) ) ;
    buf_clk cell_3755 ( .C ( clk ), .D ( signal_17619 ), .Q ( signal_18448 ) ) ;
    buf_clk cell_3757 ( .C ( clk ), .D ( signal_17621 ), .Q ( signal_18450 ) ) ;
    buf_clk cell_3759 ( .C ( clk ), .D ( signal_17623 ), .Q ( signal_18452 ) ) ;
    buf_clk cell_3761 ( .C ( clk ), .D ( signal_17625 ), .Q ( signal_18454 ) ) ;
    buf_clk cell_3763 ( .C ( clk ), .D ( signal_17627 ), .Q ( signal_18456 ) ) ;
    buf_clk cell_3765 ( .C ( clk ), .D ( signal_1145 ), .Q ( signal_18458 ) ) ;
    buf_clk cell_3767 ( .C ( clk ), .D ( signal_3236 ), .Q ( signal_18460 ) ) ;
    buf_clk cell_3769 ( .C ( clk ), .D ( signal_3237 ), .Q ( signal_18462 ) ) ;
    buf_clk cell_3771 ( .C ( clk ), .D ( signal_3238 ), .Q ( signal_18464 ) ) ;
    buf_clk cell_3773 ( .C ( clk ), .D ( signal_3239 ), .Q ( signal_18466 ) ) ;
    buf_clk cell_3777 ( .C ( clk ), .D ( signal_18469 ), .Q ( signal_18470 ) ) ;
    buf_clk cell_3781 ( .C ( clk ), .D ( signal_18473 ), .Q ( signal_18474 ) ) ;
    buf_clk cell_3785 ( .C ( clk ), .D ( signal_18477 ), .Q ( signal_18478 ) ) ;
    buf_clk cell_3789 ( .C ( clk ), .D ( signal_18481 ), .Q ( signal_18482 ) ) ;
    buf_clk cell_3793 ( .C ( clk ), .D ( signal_18485 ), .Q ( signal_18486 ) ) ;
    buf_clk cell_3795 ( .C ( clk ), .D ( signal_1095 ), .Q ( signal_18488 ) ) ;
    buf_clk cell_3797 ( .C ( clk ), .D ( signal_3036 ), .Q ( signal_18490 ) ) ;
    buf_clk cell_3799 ( .C ( clk ), .D ( signal_3037 ), .Q ( signal_18492 ) ) ;
    buf_clk cell_3801 ( .C ( clk ), .D ( signal_3038 ), .Q ( signal_18494 ) ) ;
    buf_clk cell_3803 ( .C ( clk ), .D ( signal_3039 ), .Q ( signal_18496 ) ) ;
    buf_clk cell_3805 ( .C ( clk ), .D ( signal_1078 ), .Q ( signal_18498 ) ) ;
    buf_clk cell_3807 ( .C ( clk ), .D ( signal_2968 ), .Q ( signal_18500 ) ) ;
    buf_clk cell_3809 ( .C ( clk ), .D ( signal_2969 ), .Q ( signal_18502 ) ) ;
    buf_clk cell_3811 ( .C ( clk ), .D ( signal_2970 ), .Q ( signal_18504 ) ) ;
    buf_clk cell_3813 ( .C ( clk ), .D ( signal_2971 ), .Q ( signal_18506 ) ) ;
    buf_clk cell_3815 ( .C ( clk ), .D ( signal_1073 ), .Q ( signal_18508 ) ) ;
    buf_clk cell_3817 ( .C ( clk ), .D ( signal_2948 ), .Q ( signal_18510 ) ) ;
    buf_clk cell_3819 ( .C ( clk ), .D ( signal_2949 ), .Q ( signal_18512 ) ) ;
    buf_clk cell_3821 ( .C ( clk ), .D ( signal_2950 ), .Q ( signal_18514 ) ) ;
    buf_clk cell_3823 ( .C ( clk ), .D ( signal_2951 ), .Q ( signal_18516 ) ) ;
    buf_clk cell_3825 ( .C ( clk ), .D ( signal_1158 ), .Q ( signal_18518 ) ) ;
    buf_clk cell_3827 ( .C ( clk ), .D ( signal_3288 ), .Q ( signal_18520 ) ) ;
    buf_clk cell_3829 ( .C ( clk ), .D ( signal_3289 ), .Q ( signal_18522 ) ) ;
    buf_clk cell_3831 ( .C ( clk ), .D ( signal_3290 ), .Q ( signal_18524 ) ) ;
    buf_clk cell_3833 ( .C ( clk ), .D ( signal_3291 ), .Q ( signal_18526 ) ) ;
    buf_clk cell_3835 ( .C ( clk ), .D ( signal_1020 ), .Q ( signal_18528 ) ) ;
    buf_clk cell_3837 ( .C ( clk ), .D ( signal_2736 ), .Q ( signal_18530 ) ) ;
    buf_clk cell_3839 ( .C ( clk ), .D ( signal_2737 ), .Q ( signal_18532 ) ) ;
    buf_clk cell_3841 ( .C ( clk ), .D ( signal_2738 ), .Q ( signal_18534 ) ) ;
    buf_clk cell_3843 ( .C ( clk ), .D ( signal_2739 ), .Q ( signal_18536 ) ) ;
    buf_clk cell_3845 ( .C ( clk ), .D ( signal_17749 ), .Q ( signal_18538 ) ) ;
    buf_clk cell_3847 ( .C ( clk ), .D ( signal_17751 ), .Q ( signal_18540 ) ) ;
    buf_clk cell_3849 ( .C ( clk ), .D ( signal_17753 ), .Q ( signal_18542 ) ) ;
    buf_clk cell_3851 ( .C ( clk ), .D ( signal_17755 ), .Q ( signal_18544 ) ) ;
    buf_clk cell_3853 ( .C ( clk ), .D ( signal_17757 ), .Q ( signal_18546 ) ) ;
    buf_clk cell_3855 ( .C ( clk ), .D ( signal_17559 ), .Q ( signal_18548 ) ) ;
    buf_clk cell_3857 ( .C ( clk ), .D ( signal_17561 ), .Q ( signal_18550 ) ) ;
    buf_clk cell_3859 ( .C ( clk ), .D ( signal_17563 ), .Q ( signal_18552 ) ) ;
    buf_clk cell_3861 ( .C ( clk ), .D ( signal_17565 ), .Q ( signal_18554 ) ) ;
    buf_clk cell_3863 ( .C ( clk ), .D ( signal_17567 ), .Q ( signal_18556 ) ) ;
    buf_clk cell_3865 ( .C ( clk ), .D ( signal_1162 ), .Q ( signal_18558 ) ) ;
    buf_clk cell_3867 ( .C ( clk ), .D ( signal_3304 ), .Q ( signal_18560 ) ) ;
    buf_clk cell_3869 ( .C ( clk ), .D ( signal_3305 ), .Q ( signal_18562 ) ) ;
    buf_clk cell_3871 ( .C ( clk ), .D ( signal_3306 ), .Q ( signal_18564 ) ) ;
    buf_clk cell_3873 ( .C ( clk ), .D ( signal_3307 ), .Q ( signal_18566 ) ) ;
    buf_clk cell_3875 ( .C ( clk ), .D ( signal_1071 ), .Q ( signal_18568 ) ) ;
    buf_clk cell_3877 ( .C ( clk ), .D ( signal_2940 ), .Q ( signal_18570 ) ) ;
    buf_clk cell_3879 ( .C ( clk ), .D ( signal_2941 ), .Q ( signal_18572 ) ) ;
    buf_clk cell_3881 ( .C ( clk ), .D ( signal_2942 ), .Q ( signal_18574 ) ) ;
    buf_clk cell_3883 ( .C ( clk ), .D ( signal_2943 ), .Q ( signal_18576 ) ) ;
    buf_clk cell_3887 ( .C ( clk ), .D ( signal_18579 ), .Q ( signal_18580 ) ) ;
    buf_clk cell_3891 ( .C ( clk ), .D ( signal_18583 ), .Q ( signal_18584 ) ) ;
    buf_clk cell_3895 ( .C ( clk ), .D ( signal_18587 ), .Q ( signal_18588 ) ) ;
    buf_clk cell_3899 ( .C ( clk ), .D ( signal_18591 ), .Q ( signal_18592 ) ) ;
    buf_clk cell_3903 ( .C ( clk ), .D ( signal_18595 ), .Q ( signal_18596 ) ) ;
    buf_clk cell_3905 ( .C ( clk ), .D ( signal_1081 ), .Q ( signal_18598 ) ) ;
    buf_clk cell_3907 ( .C ( clk ), .D ( signal_2980 ), .Q ( signal_18600 ) ) ;
    buf_clk cell_3909 ( .C ( clk ), .D ( signal_2981 ), .Q ( signal_18602 ) ) ;
    buf_clk cell_3911 ( .C ( clk ), .D ( signal_2982 ), .Q ( signal_18604 ) ) ;
    buf_clk cell_3913 ( .C ( clk ), .D ( signal_2983 ), .Q ( signal_18606 ) ) ;
    buf_clk cell_3915 ( .C ( clk ), .D ( signal_17679 ), .Q ( signal_18608 ) ) ;
    buf_clk cell_3917 ( .C ( clk ), .D ( signal_17681 ), .Q ( signal_18610 ) ) ;
    buf_clk cell_3919 ( .C ( clk ), .D ( signal_17683 ), .Q ( signal_18612 ) ) ;
    buf_clk cell_3921 ( .C ( clk ), .D ( signal_17685 ), .Q ( signal_18614 ) ) ;
    buf_clk cell_3923 ( .C ( clk ), .D ( signal_17687 ), .Q ( signal_18616 ) ) ;
    buf_clk cell_3925 ( .C ( clk ), .D ( signal_17629 ), .Q ( signal_18618 ) ) ;
    buf_clk cell_3927 ( .C ( clk ), .D ( signal_17631 ), .Q ( signal_18620 ) ) ;
    buf_clk cell_3929 ( .C ( clk ), .D ( signal_17633 ), .Q ( signal_18622 ) ) ;
    buf_clk cell_3931 ( .C ( clk ), .D ( signal_17635 ), .Q ( signal_18624 ) ) ;
    buf_clk cell_3933 ( .C ( clk ), .D ( signal_17637 ), .Q ( signal_18626 ) ) ;
    buf_clk cell_3935 ( .C ( clk ), .D ( signal_1304 ), .Q ( signal_18628 ) ) ;
    buf_clk cell_3937 ( .C ( clk ), .D ( signal_3872 ), .Q ( signal_18630 ) ) ;
    buf_clk cell_3939 ( .C ( clk ), .D ( signal_3873 ), .Q ( signal_18632 ) ) ;
    buf_clk cell_3941 ( .C ( clk ), .D ( signal_3874 ), .Q ( signal_18634 ) ) ;
    buf_clk cell_3943 ( .C ( clk ), .D ( signal_3875 ), .Q ( signal_18636 ) ) ;
    buf_clk cell_3945 ( .C ( clk ), .D ( signal_1250 ), .Q ( signal_18638 ) ) ;
    buf_clk cell_3947 ( .C ( clk ), .D ( signal_3656 ), .Q ( signal_18640 ) ) ;
    buf_clk cell_3949 ( .C ( clk ), .D ( signal_3657 ), .Q ( signal_18642 ) ) ;
    buf_clk cell_3951 ( .C ( clk ), .D ( signal_3658 ), .Q ( signal_18644 ) ) ;
    buf_clk cell_3953 ( .C ( clk ), .D ( signal_3659 ), .Q ( signal_18646 ) ) ;
    buf_clk cell_3955 ( .C ( clk ), .D ( signal_1327 ), .Q ( signal_18648 ) ) ;
    buf_clk cell_3957 ( .C ( clk ), .D ( signal_3964 ), .Q ( signal_18650 ) ) ;
    buf_clk cell_3959 ( .C ( clk ), .D ( signal_3965 ), .Q ( signal_18652 ) ) ;
    buf_clk cell_3961 ( .C ( clk ), .D ( signal_3966 ), .Q ( signal_18654 ) ) ;
    buf_clk cell_3963 ( .C ( clk ), .D ( signal_3967 ), .Q ( signal_18656 ) ) ;
    buf_clk cell_3985 ( .C ( clk ), .D ( signal_17789 ), .Q ( signal_18678 ) ) ;
    buf_clk cell_3989 ( .C ( clk ), .D ( signal_17791 ), .Q ( signal_18682 ) ) ;
    buf_clk cell_3993 ( .C ( clk ), .D ( signal_17793 ), .Q ( signal_18686 ) ) ;
    buf_clk cell_3997 ( .C ( clk ), .D ( signal_17795 ), .Q ( signal_18690 ) ) ;
    buf_clk cell_4001 ( .C ( clk ), .D ( signal_17797 ), .Q ( signal_18694 ) ) ;
    buf_clk cell_4015 ( .C ( clk ), .D ( signal_1290 ), .Q ( signal_18708 ) ) ;
    buf_clk cell_4019 ( .C ( clk ), .D ( signal_3816 ), .Q ( signal_18712 ) ) ;
    buf_clk cell_4023 ( .C ( clk ), .D ( signal_3817 ), .Q ( signal_18716 ) ) ;
    buf_clk cell_4027 ( .C ( clk ), .D ( signal_3818 ), .Q ( signal_18720 ) ) ;
    buf_clk cell_4031 ( .C ( clk ), .D ( signal_3819 ), .Q ( signal_18724 ) ) ;
    buf_clk cell_4035 ( .C ( clk ), .D ( signal_1354 ), .Q ( signal_18728 ) ) ;
    buf_clk cell_4039 ( .C ( clk ), .D ( signal_4072 ), .Q ( signal_18732 ) ) ;
    buf_clk cell_4043 ( .C ( clk ), .D ( signal_4073 ), .Q ( signal_18736 ) ) ;
    buf_clk cell_4047 ( .C ( clk ), .D ( signal_4074 ), .Q ( signal_18740 ) ) ;
    buf_clk cell_4051 ( .C ( clk ), .D ( signal_4075 ), .Q ( signal_18744 ) ) ;
    buf_clk cell_4055 ( .C ( clk ), .D ( signal_1234 ), .Q ( signal_18748 ) ) ;
    buf_clk cell_4059 ( .C ( clk ), .D ( signal_3592 ), .Q ( signal_18752 ) ) ;
    buf_clk cell_4063 ( .C ( clk ), .D ( signal_3593 ), .Q ( signal_18756 ) ) ;
    buf_clk cell_4067 ( .C ( clk ), .D ( signal_3594 ), .Q ( signal_18760 ) ) ;
    buf_clk cell_4071 ( .C ( clk ), .D ( signal_3595 ), .Q ( signal_18764 ) ) ;
    buf_clk cell_4079 ( .C ( clk ), .D ( signal_18771 ), .Q ( signal_18772 ) ) ;
    buf_clk cell_4087 ( .C ( clk ), .D ( signal_18779 ), .Q ( signal_18780 ) ) ;
    buf_clk cell_4095 ( .C ( clk ), .D ( signal_18787 ), .Q ( signal_18788 ) ) ;
    buf_clk cell_4103 ( .C ( clk ), .D ( signal_18795 ), .Q ( signal_18796 ) ) ;
    buf_clk cell_4111 ( .C ( clk ), .D ( signal_18803 ), .Q ( signal_18804 ) ) ;
    buf_clk cell_4135 ( .C ( clk ), .D ( signal_1313 ), .Q ( signal_18828 ) ) ;
    buf_clk cell_4139 ( .C ( clk ), .D ( signal_3908 ), .Q ( signal_18832 ) ) ;
    buf_clk cell_4143 ( .C ( clk ), .D ( signal_3909 ), .Q ( signal_18836 ) ) ;
    buf_clk cell_4147 ( .C ( clk ), .D ( signal_3910 ), .Q ( signal_18840 ) ) ;
    buf_clk cell_4151 ( .C ( clk ), .D ( signal_3911 ), .Q ( signal_18844 ) ) ;
    buf_clk cell_4175 ( .C ( clk ), .D ( signal_1335 ), .Q ( signal_18868 ) ) ;
    buf_clk cell_4179 ( .C ( clk ), .D ( signal_3996 ), .Q ( signal_18872 ) ) ;
    buf_clk cell_4183 ( .C ( clk ), .D ( signal_3997 ), .Q ( signal_18876 ) ) ;
    buf_clk cell_4187 ( .C ( clk ), .D ( signal_3998 ), .Q ( signal_18880 ) ) ;
    buf_clk cell_4191 ( .C ( clk ), .D ( signal_3999 ), .Q ( signal_18884 ) ) ;
    buf_clk cell_4245 ( .C ( clk ), .D ( signal_1061 ), .Q ( signal_18938 ) ) ;
    buf_clk cell_4249 ( .C ( clk ), .D ( signal_2900 ), .Q ( signal_18942 ) ) ;
    buf_clk cell_4253 ( .C ( clk ), .D ( signal_2901 ), .Q ( signal_18946 ) ) ;
    buf_clk cell_4257 ( .C ( clk ), .D ( signal_2902 ), .Q ( signal_18950 ) ) ;
    buf_clk cell_4261 ( .C ( clk ), .D ( signal_2903 ), .Q ( signal_18954 ) ) ;
    buf_clk cell_4305 ( .C ( clk ), .D ( signal_1361 ), .Q ( signal_18998 ) ) ;
    buf_clk cell_4309 ( .C ( clk ), .D ( signal_4100 ), .Q ( signal_19002 ) ) ;
    buf_clk cell_4313 ( .C ( clk ), .D ( signal_4101 ), .Q ( signal_19006 ) ) ;
    buf_clk cell_4317 ( .C ( clk ), .D ( signal_4102 ), .Q ( signal_19010 ) ) ;
    buf_clk cell_4321 ( .C ( clk ), .D ( signal_4103 ), .Q ( signal_19014 ) ) ;
    buf_clk cell_4345 ( .C ( clk ), .D ( signal_17359 ), .Q ( signal_19038 ) ) ;
    buf_clk cell_4349 ( .C ( clk ), .D ( signal_17361 ), .Q ( signal_19042 ) ) ;
    buf_clk cell_4353 ( .C ( clk ), .D ( signal_17363 ), .Q ( signal_19046 ) ) ;
    buf_clk cell_4357 ( .C ( clk ), .D ( signal_17365 ), .Q ( signal_19050 ) ) ;
    buf_clk cell_4361 ( .C ( clk ), .D ( signal_17367 ), .Q ( signal_19054 ) ) ;
    buf_clk cell_4365 ( .C ( clk ), .D ( signal_17409 ), .Q ( signal_19058 ) ) ;
    buf_clk cell_4369 ( .C ( clk ), .D ( signal_17411 ), .Q ( signal_19062 ) ) ;
    buf_clk cell_4373 ( .C ( clk ), .D ( signal_17413 ), .Q ( signal_19066 ) ) ;
    buf_clk cell_4377 ( .C ( clk ), .D ( signal_17415 ), .Q ( signal_19070 ) ) ;
    buf_clk cell_4381 ( .C ( clk ), .D ( signal_17417 ), .Q ( signal_19074 ) ) ;
    buf_clk cell_4385 ( .C ( clk ), .D ( signal_17589 ), .Q ( signal_19078 ) ) ;
    buf_clk cell_4389 ( .C ( clk ), .D ( signal_17591 ), .Q ( signal_19082 ) ) ;
    buf_clk cell_4393 ( .C ( clk ), .D ( signal_17593 ), .Q ( signal_19086 ) ) ;
    buf_clk cell_4397 ( .C ( clk ), .D ( signal_17595 ), .Q ( signal_19090 ) ) ;
    buf_clk cell_4401 ( .C ( clk ), .D ( signal_17597 ), .Q ( signal_19094 ) ) ;
    buf_clk cell_4405 ( .C ( clk ), .D ( signal_17289 ), .Q ( signal_19098 ) ) ;
    buf_clk cell_4409 ( .C ( clk ), .D ( signal_17291 ), .Q ( signal_19102 ) ) ;
    buf_clk cell_4413 ( .C ( clk ), .D ( signal_17293 ), .Q ( signal_19106 ) ) ;
    buf_clk cell_4417 ( .C ( clk ), .D ( signal_17295 ), .Q ( signal_19110 ) ) ;
    buf_clk cell_4421 ( .C ( clk ), .D ( signal_17297 ), .Q ( signal_19114 ) ) ;
    buf_clk cell_4475 ( .C ( clk ), .D ( signal_17319 ), .Q ( signal_19168 ) ) ;
    buf_clk cell_4479 ( .C ( clk ), .D ( signal_17321 ), .Q ( signal_19172 ) ) ;
    buf_clk cell_4483 ( .C ( clk ), .D ( signal_17323 ), .Q ( signal_19176 ) ) ;
    buf_clk cell_4487 ( .C ( clk ), .D ( signal_17325 ), .Q ( signal_19180 ) ) ;
    buf_clk cell_4491 ( .C ( clk ), .D ( signal_17327 ), .Q ( signal_19184 ) ) ;
    buf_clk cell_4495 ( .C ( clk ), .D ( signal_17309 ), .Q ( signal_19188 ) ) ;
    buf_clk cell_4499 ( .C ( clk ), .D ( signal_17311 ), .Q ( signal_19192 ) ) ;
    buf_clk cell_4503 ( .C ( clk ), .D ( signal_17313 ), .Q ( signal_19196 ) ) ;
    buf_clk cell_4507 ( .C ( clk ), .D ( signal_17315 ), .Q ( signal_19200 ) ) ;
    buf_clk cell_4511 ( .C ( clk ), .D ( signal_17317 ), .Q ( signal_19204 ) ) ;
    buf_clk cell_4515 ( .C ( clk ), .D ( signal_17499 ), .Q ( signal_19208 ) ) ;
    buf_clk cell_4519 ( .C ( clk ), .D ( signal_17501 ), .Q ( signal_19212 ) ) ;
    buf_clk cell_4523 ( .C ( clk ), .D ( signal_17503 ), .Q ( signal_19216 ) ) ;
    buf_clk cell_4527 ( .C ( clk ), .D ( signal_17505 ), .Q ( signal_19220 ) ) ;
    buf_clk cell_4531 ( .C ( clk ), .D ( signal_17507 ), .Q ( signal_19224 ) ) ;
    buf_clk cell_4545 ( .C ( clk ), .D ( signal_17399 ), .Q ( signal_19238 ) ) ;
    buf_clk cell_4549 ( .C ( clk ), .D ( signal_17401 ), .Q ( signal_19242 ) ) ;
    buf_clk cell_4553 ( .C ( clk ), .D ( signal_17403 ), .Q ( signal_19246 ) ) ;
    buf_clk cell_4557 ( .C ( clk ), .D ( signal_17405 ), .Q ( signal_19250 ) ) ;
    buf_clk cell_4561 ( .C ( clk ), .D ( signal_17407 ), .Q ( signal_19254 ) ) ;
    buf_clk cell_4615 ( .C ( clk ), .D ( signal_1080 ), .Q ( signal_19308 ) ) ;
    buf_clk cell_4619 ( .C ( clk ), .D ( signal_2976 ), .Q ( signal_19312 ) ) ;
    buf_clk cell_4623 ( .C ( clk ), .D ( signal_2977 ), .Q ( signal_19316 ) ) ;
    buf_clk cell_4627 ( .C ( clk ), .D ( signal_2978 ), .Q ( signal_19320 ) ) ;
    buf_clk cell_4631 ( .C ( clk ), .D ( signal_2979 ), .Q ( signal_19324 ) ) ;
    buf_clk cell_4635 ( .C ( clk ), .D ( signal_1365 ), .Q ( signal_19328 ) ) ;
    buf_clk cell_4639 ( .C ( clk ), .D ( signal_4116 ), .Q ( signal_19332 ) ) ;
    buf_clk cell_4643 ( .C ( clk ), .D ( signal_4117 ), .Q ( signal_19336 ) ) ;
    buf_clk cell_4647 ( .C ( clk ), .D ( signal_4118 ), .Q ( signal_19340 ) ) ;
    buf_clk cell_4651 ( .C ( clk ), .D ( signal_4119 ), .Q ( signal_19344 ) ) ;
    buf_clk cell_4665 ( .C ( clk ), .D ( signal_1242 ), .Q ( signal_19358 ) ) ;
    buf_clk cell_4669 ( .C ( clk ), .D ( signal_3624 ), .Q ( signal_19362 ) ) ;
    buf_clk cell_4673 ( .C ( clk ), .D ( signal_3625 ), .Q ( signal_19366 ) ) ;
    buf_clk cell_4677 ( .C ( clk ), .D ( signal_3626 ), .Q ( signal_19370 ) ) ;
    buf_clk cell_4681 ( .C ( clk ), .D ( signal_3627 ), .Q ( signal_19374 ) ) ;
    buf_clk cell_4705 ( .C ( clk ), .D ( signal_1296 ), .Q ( signal_19398 ) ) ;
    buf_clk cell_4709 ( .C ( clk ), .D ( signal_3840 ), .Q ( signal_19402 ) ) ;
    buf_clk cell_4713 ( .C ( clk ), .D ( signal_3841 ), .Q ( signal_19406 ) ) ;
    buf_clk cell_4717 ( .C ( clk ), .D ( signal_3842 ), .Q ( signal_19410 ) ) ;
    buf_clk cell_4721 ( .C ( clk ), .D ( signal_3843 ), .Q ( signal_19414 ) ) ;
    buf_clk cell_4725 ( .C ( clk ), .D ( signal_1308 ), .Q ( signal_19418 ) ) ;
    buf_clk cell_4729 ( .C ( clk ), .D ( signal_3888 ), .Q ( signal_19422 ) ) ;
    buf_clk cell_4733 ( .C ( clk ), .D ( signal_3889 ), .Q ( signal_19426 ) ) ;
    buf_clk cell_4737 ( .C ( clk ), .D ( signal_3890 ), .Q ( signal_19430 ) ) ;
    buf_clk cell_4741 ( .C ( clk ), .D ( signal_3891 ), .Q ( signal_19434 ) ) ;
    buf_clk cell_4745 ( .C ( clk ), .D ( signal_1251 ), .Q ( signal_19438 ) ) ;
    buf_clk cell_4749 ( .C ( clk ), .D ( signal_3660 ), .Q ( signal_19442 ) ) ;
    buf_clk cell_4753 ( .C ( clk ), .D ( signal_3661 ), .Q ( signal_19446 ) ) ;
    buf_clk cell_4757 ( .C ( clk ), .D ( signal_3662 ), .Q ( signal_19450 ) ) ;
    buf_clk cell_4761 ( .C ( clk ), .D ( signal_3663 ), .Q ( signal_19454 ) ) ;
    buf_clk cell_4775 ( .C ( clk ), .D ( signal_1326 ), .Q ( signal_19468 ) ) ;
    buf_clk cell_4779 ( .C ( clk ), .D ( signal_3960 ), .Q ( signal_19472 ) ) ;
    buf_clk cell_4783 ( .C ( clk ), .D ( signal_3961 ), .Q ( signal_19476 ) ) ;
    buf_clk cell_4787 ( .C ( clk ), .D ( signal_3962 ), .Q ( signal_19480 ) ) ;
    buf_clk cell_4791 ( .C ( clk ), .D ( signal_3963 ), .Q ( signal_19484 ) ) ;
    buf_clk cell_4795 ( .C ( clk ), .D ( signal_1261 ), .Q ( signal_19488 ) ) ;
    buf_clk cell_4799 ( .C ( clk ), .D ( signal_3700 ), .Q ( signal_19492 ) ) ;
    buf_clk cell_4803 ( .C ( clk ), .D ( signal_3701 ), .Q ( signal_19496 ) ) ;
    buf_clk cell_4807 ( .C ( clk ), .D ( signal_3702 ), .Q ( signal_19500 ) ) ;
    buf_clk cell_4811 ( .C ( clk ), .D ( signal_3703 ), .Q ( signal_19504 ) ) ;
    buf_clk cell_4825 ( .C ( clk ), .D ( signal_1271 ), .Q ( signal_19518 ) ) ;
    buf_clk cell_4829 ( .C ( clk ), .D ( signal_3740 ), .Q ( signal_19522 ) ) ;
    buf_clk cell_4833 ( .C ( clk ), .D ( signal_3741 ), .Q ( signal_19526 ) ) ;
    buf_clk cell_4837 ( .C ( clk ), .D ( signal_3742 ), .Q ( signal_19530 ) ) ;
    buf_clk cell_4841 ( .C ( clk ), .D ( signal_3743 ), .Q ( signal_19534 ) ) ;
    buf_clk cell_4875 ( .C ( clk ), .D ( signal_17269 ), .Q ( signal_19568 ) ) ;
    buf_clk cell_4879 ( .C ( clk ), .D ( signal_17271 ), .Q ( signal_19572 ) ) ;
    buf_clk cell_4883 ( .C ( clk ), .D ( signal_17273 ), .Q ( signal_19576 ) ) ;
    buf_clk cell_4887 ( .C ( clk ), .D ( signal_17275 ), .Q ( signal_19580 ) ) ;
    buf_clk cell_4891 ( .C ( clk ), .D ( signal_17277 ), .Q ( signal_19584 ) ) ;
    buf_clk cell_4905 ( .C ( clk ), .D ( signal_17799 ), .Q ( signal_19598 ) ) ;
    buf_clk cell_4911 ( .C ( clk ), .D ( signal_17801 ), .Q ( signal_19604 ) ) ;
    buf_clk cell_4917 ( .C ( clk ), .D ( signal_17803 ), .Q ( signal_19610 ) ) ;
    buf_clk cell_4923 ( .C ( clk ), .D ( signal_17805 ), .Q ( signal_19616 ) ) ;
    buf_clk cell_4929 ( .C ( clk ), .D ( signal_17807 ), .Q ( signal_19622 ) ) ;
    buf_clk cell_4935 ( .C ( clk ), .D ( signal_1248 ), .Q ( signal_19628 ) ) ;
    buf_clk cell_4941 ( .C ( clk ), .D ( signal_3648 ), .Q ( signal_19634 ) ) ;
    buf_clk cell_4947 ( .C ( clk ), .D ( signal_3649 ), .Q ( signal_19640 ) ) ;
    buf_clk cell_4953 ( .C ( clk ), .D ( signal_3650 ), .Q ( signal_19646 ) ) ;
    buf_clk cell_4959 ( .C ( clk ), .D ( signal_3651 ), .Q ( signal_19652 ) ) ;
    buf_clk cell_4965 ( .C ( clk ), .D ( signal_1314 ), .Q ( signal_19658 ) ) ;
    buf_clk cell_4971 ( .C ( clk ), .D ( signal_3912 ), .Q ( signal_19664 ) ) ;
    buf_clk cell_4977 ( .C ( clk ), .D ( signal_3913 ), .Q ( signal_19670 ) ) ;
    buf_clk cell_4983 ( .C ( clk ), .D ( signal_3914 ), .Q ( signal_19676 ) ) ;
    buf_clk cell_4989 ( .C ( clk ), .D ( signal_3915 ), .Q ( signal_19682 ) ) ;
    buf_clk cell_5015 ( .C ( clk ), .D ( signal_1336 ), .Q ( signal_19708 ) ) ;
    buf_clk cell_5021 ( .C ( clk ), .D ( signal_4000 ), .Q ( signal_19714 ) ) ;
    buf_clk cell_5027 ( .C ( clk ), .D ( signal_4001 ), .Q ( signal_19720 ) ) ;
    buf_clk cell_5033 ( .C ( clk ), .D ( signal_4002 ), .Q ( signal_19726 ) ) ;
    buf_clk cell_5039 ( .C ( clk ), .D ( signal_4003 ), .Q ( signal_19732 ) ) ;
    buf_clk cell_5145 ( .C ( clk ), .D ( signal_17509 ), .Q ( signal_19838 ) ) ;
    buf_clk cell_5151 ( .C ( clk ), .D ( signal_17511 ), .Q ( signal_19844 ) ) ;
    buf_clk cell_5157 ( .C ( clk ), .D ( signal_17513 ), .Q ( signal_19850 ) ) ;
    buf_clk cell_5163 ( .C ( clk ), .D ( signal_17515 ), .Q ( signal_19856 ) ) ;
    buf_clk cell_5169 ( .C ( clk ), .D ( signal_17517 ), .Q ( signal_19862 ) ) ;
    buf_clk cell_5295 ( .C ( clk ), .D ( signal_17239 ), .Q ( signal_19988 ) ) ;
    buf_clk cell_5301 ( .C ( clk ), .D ( signal_17241 ), .Q ( signal_19994 ) ) ;
    buf_clk cell_5307 ( .C ( clk ), .D ( signal_17243 ), .Q ( signal_20000 ) ) ;
    buf_clk cell_5313 ( .C ( clk ), .D ( signal_17245 ), .Q ( signal_20006 ) ) ;
    buf_clk cell_5319 ( .C ( clk ), .D ( signal_17247 ), .Q ( signal_20012 ) ) ;
    buf_clk cell_5375 ( .C ( clk ), .D ( signal_1298 ), .Q ( signal_20068 ) ) ;
    buf_clk cell_5381 ( .C ( clk ), .D ( signal_3848 ), .Q ( signal_20074 ) ) ;
    buf_clk cell_5387 ( .C ( clk ), .D ( signal_3849 ), .Q ( signal_20080 ) ) ;
    buf_clk cell_5393 ( .C ( clk ), .D ( signal_3850 ), .Q ( signal_20086 ) ) ;
    buf_clk cell_5399 ( .C ( clk ), .D ( signal_3851 ), .Q ( signal_20092 ) ) ;
    buf_clk cell_5515 ( .C ( clk ), .D ( signal_1064 ), .Q ( signal_20208 ) ) ;
    buf_clk cell_5521 ( .C ( clk ), .D ( signal_2912 ), .Q ( signal_20214 ) ) ;
    buf_clk cell_5527 ( .C ( clk ), .D ( signal_2913 ), .Q ( signal_20220 ) ) ;
    buf_clk cell_5533 ( .C ( clk ), .D ( signal_2914 ), .Q ( signal_20226 ) ) ;
    buf_clk cell_5539 ( .C ( clk ), .D ( signal_2915 ), .Q ( signal_20232 ) ) ;
    buf_clk cell_5565 ( .C ( clk ), .D ( signal_1316 ), .Q ( signal_20258 ) ) ;
    buf_clk cell_5571 ( .C ( clk ), .D ( signal_3920 ), .Q ( signal_20264 ) ) ;
    buf_clk cell_5577 ( .C ( clk ), .D ( signal_3921 ), .Q ( signal_20270 ) ) ;
    buf_clk cell_5583 ( .C ( clk ), .D ( signal_3922 ), .Q ( signal_20276 ) ) ;
    buf_clk cell_5589 ( .C ( clk ), .D ( signal_3923 ), .Q ( signal_20282 ) ) ;
    buf_clk cell_5705 ( .C ( clk ), .D ( signal_1289 ), .Q ( signal_20398 ) ) ;
    buf_clk cell_5711 ( .C ( clk ), .D ( signal_3812 ), .Q ( signal_20404 ) ) ;
    buf_clk cell_5717 ( .C ( clk ), .D ( signal_3813 ), .Q ( signal_20410 ) ) ;
    buf_clk cell_5723 ( .C ( clk ), .D ( signal_3814 ), .Q ( signal_20416 ) ) ;
    buf_clk cell_5729 ( .C ( clk ), .D ( signal_3815 ), .Q ( signal_20422 ) ) ;
    buf_clk cell_5775 ( .C ( clk ), .D ( signal_1359 ), .Q ( signal_20468 ) ) ;
    buf_clk cell_5781 ( .C ( clk ), .D ( signal_4092 ), .Q ( signal_20474 ) ) ;
    buf_clk cell_5787 ( .C ( clk ), .D ( signal_4093 ), .Q ( signal_20480 ) ) ;
    buf_clk cell_5793 ( .C ( clk ), .D ( signal_4094 ), .Q ( signal_20486 ) ) ;
    buf_clk cell_5799 ( .C ( clk ), .D ( signal_4095 ), .Q ( signal_20492 ) ) ;
    buf_clk cell_5805 ( .C ( clk ), .D ( signal_1307 ), .Q ( signal_20498 ) ) ;
    buf_clk cell_5811 ( .C ( clk ), .D ( signal_3884 ), .Q ( signal_20504 ) ) ;
    buf_clk cell_5817 ( .C ( clk ), .D ( signal_3885 ), .Q ( signal_20510 ) ) ;
    buf_clk cell_5823 ( .C ( clk ), .D ( signal_3886 ), .Q ( signal_20516 ) ) ;
    buf_clk cell_5829 ( .C ( clk ), .D ( signal_3887 ), .Q ( signal_20522 ) ) ;
    buf_clk cell_5835 ( .C ( clk ), .D ( signal_17599 ), .Q ( signal_20528 ) ) ;
    buf_clk cell_5841 ( .C ( clk ), .D ( signal_17601 ), .Q ( signal_20534 ) ) ;
    buf_clk cell_5847 ( .C ( clk ), .D ( signal_17603 ), .Q ( signal_20540 ) ) ;
    buf_clk cell_5853 ( .C ( clk ), .D ( signal_17605 ), .Q ( signal_20546 ) ) ;
    buf_clk cell_5859 ( .C ( clk ), .D ( signal_17607 ), .Q ( signal_20552 ) ) ;
    buf_clk cell_5905 ( .C ( clk ), .D ( signal_1315 ), .Q ( signal_20598 ) ) ;
    buf_clk cell_5913 ( .C ( clk ), .D ( signal_3916 ), .Q ( signal_20606 ) ) ;
    buf_clk cell_5921 ( .C ( clk ), .D ( signal_3917 ), .Q ( signal_20614 ) ) ;
    buf_clk cell_5929 ( .C ( clk ), .D ( signal_3918 ), .Q ( signal_20622 ) ) ;
    buf_clk cell_5937 ( .C ( clk ), .D ( signal_3919 ), .Q ( signal_20630 ) ) ;
    buf_clk cell_6335 ( .C ( clk ), .D ( signal_1239 ), .Q ( signal_21028 ) ) ;
    buf_clk cell_6343 ( .C ( clk ), .D ( signal_3612 ), .Q ( signal_21036 ) ) ;
    buf_clk cell_6351 ( .C ( clk ), .D ( signal_3613 ), .Q ( signal_21044 ) ) ;
    buf_clk cell_6359 ( .C ( clk ), .D ( signal_3614 ), .Q ( signal_21052 ) ) ;
    buf_clk cell_6367 ( .C ( clk ), .D ( signal_3615 ), .Q ( signal_21060 ) ) ;
    buf_clk cell_6495 ( .C ( clk ), .D ( signal_1060 ), .Q ( signal_21188 ) ) ;
    buf_clk cell_6503 ( .C ( clk ), .D ( signal_2896 ), .Q ( signal_21196 ) ) ;
    buf_clk cell_6511 ( .C ( clk ), .D ( signal_2897 ), .Q ( signal_21204 ) ) ;
    buf_clk cell_6519 ( .C ( clk ), .D ( signal_2898 ), .Q ( signal_21212 ) ) ;
    buf_clk cell_6527 ( .C ( clk ), .D ( signal_2899 ), .Q ( signal_21220 ) ) ;
    buf_clk cell_6745 ( .C ( clk ), .D ( signal_1254 ), .Q ( signal_21438 ) ) ;
    buf_clk cell_6755 ( .C ( clk ), .D ( signal_3672 ), .Q ( signal_21448 ) ) ;
    buf_clk cell_6765 ( .C ( clk ), .D ( signal_3673 ), .Q ( signal_21458 ) ) ;
    buf_clk cell_6775 ( .C ( clk ), .D ( signal_3674 ), .Q ( signal_21468 ) ) ;
    buf_clk cell_6785 ( .C ( clk ), .D ( signal_3675 ), .Q ( signal_21478 ) ) ;
    buf_clk cell_6985 ( .C ( clk ), .D ( signal_1247 ), .Q ( signal_21678 ) ) ;
    buf_clk cell_6995 ( .C ( clk ), .D ( signal_3644 ), .Q ( signal_21688 ) ) ;
    buf_clk cell_7005 ( .C ( clk ), .D ( signal_3645 ), .Q ( signal_21698 ) ) ;
    buf_clk cell_7015 ( .C ( clk ), .D ( signal_3646 ), .Q ( signal_21708 ) ) ;
    buf_clk cell_7025 ( .C ( clk ), .D ( signal_3647 ), .Q ( signal_21718 ) ) ;
    buf_clk cell_7265 ( .C ( clk ), .D ( signal_1066 ), .Q ( signal_21958 ) ) ;
    buf_clk cell_7275 ( .C ( clk ), .D ( signal_2920 ), .Q ( signal_21968 ) ) ;
    buf_clk cell_7285 ( .C ( clk ), .D ( signal_2921 ), .Q ( signal_21978 ) ) ;
    buf_clk cell_7295 ( .C ( clk ), .D ( signal_2922 ), .Q ( signal_21988 ) ) ;
    buf_clk cell_7305 ( .C ( clk ), .D ( signal_2923 ), .Q ( signal_21998 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1085 ( .a ({signal_17227, signal_17223, signal_17219, signal_17215, signal_17211}), .b ({signal_2715, signal_2714, signal_2713, signal_2712, signal_1014}), .clk ( clk ), .r ({Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .c ({signal_3059, signal_3058, signal_3057, signal_3056, signal_1100}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1124 ( .a ({signal_17237, signal_17235, signal_17233, signal_17231, signal_17229}), .b ({signal_2735, signal_2734, signal_2733, signal_2732, signal_1019}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390]}), .c ({signal_3215, signal_3214, signal_3213, signal_3212, signal_1139}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1132 ( .a ({signal_17247, signal_17245, signal_17243, signal_17241, signal_17239}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_3247, signal_3246, signal_3245, signal_3244, signal_1147}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1140 ( .a ({signal_17257, signal_17255, signal_17253, signal_17251, signal_17249}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410]}), .c ({signal_3279, signal_3278, signal_3277, signal_3276, signal_1155}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1155 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1020}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .c ({signal_3339, signal_3338, signal_3337, signal_3336, signal_1170}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1173 ( .a ({signal_17277, signal_17275, signal_17273, signal_17271, signal_17269}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_3411, signal_3410, signal_3409, signal_3408, signal_1188}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1184 ( .a ({signal_17287, signal_17285, signal_17283, signal_17281, signal_17279}), .b ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1024}), .clk ( clk ), .r ({Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .c ({signal_3455, signal_3454, signal_3453, signal_3452, signal_1199}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1189 ( .a ({signal_17297, signal_17295, signal_17293, signal_17291, signal_17289}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450]}), .c ({signal_3475, signal_3474, signal_3473, signal_3472, signal_1204}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1190 ( .a ({signal_17307, signal_17305, signal_17303, signal_17301, signal_17299}), .b ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1024}), .clk ( clk ), .r ({Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_3479, signal_3478, signal_3477, signal_3476, signal_1205}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1198 ( .a ({signal_17317, signal_17315, signal_17313, signal_17311, signal_17309}), .b ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1024}), .clk ( clk ), .r ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470]}), .c ({signal_3511, signal_3510, signal_3509, signal_3508, signal_1213}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1207 ( .a ({signal_17327, signal_17325, signal_17323, signal_17321, signal_17319}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .c ({signal_3547, signal_3546, signal_3545, signal_3544, signal_1222}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1209 ( .a ({signal_17337, signal_17335, signal_17333, signal_17331, signal_17329}), .b ({signal_2763, signal_2762, signal_2761, signal_2760, signal_1026}), .clk ( clk ), .r ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_3555, signal_3554, signal_3553, signal_3552, signal_1224}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1211 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1020}), .clk ( clk ), .r ({Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .c ({signal_3563, signal_3562, signal_3561, signal_3560, signal_1226}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1212 ( .a ({signal_17357, signal_17355, signal_17353, signal_17351, signal_17349}), .b ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1020}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510]}), .c ({signal_3567, signal_3566, signal_3565, signal_3564, signal_1227}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1243 ( .a ({signal_3059, signal_3058, signal_3057, signal_3056, signal_1100}), .b ({signal_3691, signal_3690, signal_3689, signal_3688, signal_1258}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1272 ( .a ({signal_3215, signal_3214, signal_3213, signal_3212, signal_1139}), .b ({signal_3807, signal_3806, signal_3805, signal_3804, signal_1287}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1277 ( .a ({signal_3247, signal_3246, signal_3245, signal_3244, signal_1147}), .b ({signal_3827, signal_3826, signal_3825, signal_3824, signal_1292}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1284 ( .a ({signal_3279, signal_3278, signal_3277, signal_3276, signal_1155}), .b ({signal_3855, signal_3854, signal_3853, signal_3852, signal_1299}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1297 ( .a ({signal_3339, signal_3338, signal_3337, signal_3336, signal_1170}), .b ({signal_3907, signal_3906, signal_3905, signal_3904, signal_1312}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1314 ( .a ({signal_3411, signal_3410, signal_3409, signal_3408, signal_1188}), .b ({signal_3975, signal_3974, signal_3973, signal_3972, signal_1329}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1323 ( .a ({signal_3455, signal_3454, signal_3453, signal_3452, signal_1199}), .b ({signal_4011, signal_4010, signal_4009, signal_4008, signal_1338}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1328 ( .a ({signal_3475, signal_3474, signal_3473, signal_3472, signal_1204}), .b ({signal_4031, signal_4030, signal_4029, signal_4028, signal_1343}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1329 ( .a ({signal_3479, signal_3478, signal_3477, signal_3476, signal_1205}), .b ({signal_4035, signal_4034, signal_4033, signal_4032, signal_1344}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1335 ( .a ({signal_3511, signal_3510, signal_3509, signal_3508, signal_1213}), .b ({signal_4059, signal_4058, signal_4057, signal_4056, signal_1350}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1343 ( .a ({signal_3547, signal_3546, signal_3545, signal_3544, signal_1222}), .b ({signal_4091, signal_4090, signal_4089, signal_4088, signal_1358}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1345 ( .a ({signal_3555, signal_3554, signal_3553, signal_3552, signal_1224}), .b ({signal_4099, signal_4098, signal_4097, signal_4096, signal_1360}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1347 ( .a ({signal_3563, signal_3562, signal_3561, signal_3560, signal_1226}), .b ({signal_4107, signal_4106, signal_4105, signal_4104, signal_1362}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1348 ( .a ({signal_3567, signal_3566, signal_3565, signal_3564, signal_1227}), .b ({signal_4111, signal_4110, signal_4109, signal_4108, signal_1363}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1351 ( .a ({signal_17367, signal_17365, signal_17363, signal_17361, signal_17359}), .b ({signal_2927, signal_2926, signal_2925, signal_2924, signal_1067}), .clk ( clk ), .r ({Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_4123, signal_4122, signal_4121, signal_4120, signal_1366}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1352 ( .a ({signal_17377, signal_17375, signal_17373, signal_17371, signal_17369}), .b ({signal_2931, signal_2930, signal_2929, signal_2928, signal_1068}), .clk ( clk ), .r ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530]}), .c ({signal_4127, signal_4126, signal_4125, signal_4124, signal_1367}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1358 ( .a ({signal_17277, signal_17275, signal_17273, signal_17271, signal_17269}), .b ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1080}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .c ({signal_4151, signal_4150, signal_4149, signal_4148, signal_1373}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1359 ( .a ({signal_17327, signal_17325, signal_17323, signal_17321, signal_17319}), .b ({signal_2999, signal_2998, signal_2997, signal_2996, signal_1085}), .clk ( clk ), .r ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_4155, signal_4154, signal_4153, signal_4152, signal_1374}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1363 ( .a ({signal_17307, signal_17305, signal_17303, signal_17301, signal_17299}), .b ({signal_3015, signal_3014, signal_3013, signal_3012, signal_1089}), .clk ( clk ), .r ({Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .c ({signal_4171, signal_4170, signal_4169, signal_4168, signal_1378}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1364 ( .a ({signal_17387, signal_17385, signal_17383, signal_17381, signal_17379}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570]}), .c ({signal_4175, signal_4174, signal_4173, signal_4172, signal_1379}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1370 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .clk ( clk ), .r ({Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_4199, signal_4198, signal_4197, signal_4196, signal_1385}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1371 ( .a ({signal_17407, signal_17405, signal_17403, signal_17401, signal_17399}), .b ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .clk ( clk ), .r ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590]}), .c ({signal_4203, signal_4202, signal_4201, signal_4200, signal_1386}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1372 ( .a ({signal_17417, signal_17415, signal_17413, signal_17411, signal_17409}), .b ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .c ({signal_4207, signal_4206, signal_4205, signal_4204, signal_1387}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1373 ( .a ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_4211, signal_4210, signal_4209, signal_4208, signal_1388}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1374 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3047, signal_3046, signal_3045, signal_3044, signal_1097}), .clk ( clk ), .r ({Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .c ({signal_4215, signal_4214, signal_4213, signal_4212, signal_1389}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1377 ( .a ({signal_17437, signal_17435, signal_17433, signal_17431, signal_17429}), .b ({signal_3075, signal_3074, signal_3073, signal_3072, signal_1104}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630]}), .c ({signal_4227, signal_4226, signal_4225, signal_4224, signal_1392}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1378 ( .a ({signal_17447, signal_17445, signal_17443, signal_17441, signal_17439}), .b ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1078}), .clk ( clk ), .r ({Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_4231, signal_4230, signal_4229, signal_4228, signal_1393}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1379 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650]}), .c ({signal_4235, signal_4234, signal_4233, signal_4232, signal_1394}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1380 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3015, signal_3014, signal_3013, signal_3012, signal_1089}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .c ({signal_4239, signal_4238, signal_4237, signal_4236, signal_1395}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1381 ( .a ({signal_17307, signal_17305, signal_17303, signal_17301, signal_17299}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_4243, signal_4242, signal_4241, signal_4240, signal_1396}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1382 ( .a ({signal_17457, signal_17455, signal_17453, signal_17451, signal_17449}), .b ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .clk ( clk ), .r ({Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .c ({signal_4247, signal_4246, signal_4245, signal_4244, signal_1397}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1384 ( .a ({signal_17467, signal_17465, signal_17463, signal_17461, signal_17459}), .b ({signal_3087, signal_3086, signal_3085, signal_3084, signal_1107}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690]}), .c ({signal_4255, signal_4254, signal_4253, signal_4252, signal_1399}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1385 ( .a ({signal_17287, signal_17285, signal_17283, signal_17281, signal_17279}), .b ({signal_3027, signal_3026, signal_3025, signal_3024, signal_1092}), .clk ( clk ), .r ({Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_4259, signal_4258, signal_4257, signal_4256, signal_1400}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1386 ( .a ({signal_17477, signal_17475, signal_17473, signal_17471, signal_17469}), .b ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1080}), .clk ( clk ), .r ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710]}), .c ({signal_4263, signal_4262, signal_4261, signal_4260, signal_1401}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1387 ( .a ({signal_17487, signal_17485, signal_17483, signal_17481, signal_17479}), .b ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .c ({signal_4267, signal_4266, signal_4265, signal_4264, signal_1402}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1388 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_3115, signal_3114, signal_3113, signal_3112, signal_1114}), .clk ( clk ), .r ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_4271, signal_4270, signal_4269, signal_4268, signal_1403}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1389 ( .a ({signal_17507, signal_17505, signal_17503, signal_17501, signal_17499}), .b ({signal_3091, signal_3090, signal_3089, signal_3088, signal_1108}), .clk ( clk ), .r ({Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .c ({signal_4275, signal_4274, signal_4273, signal_4272, signal_1404}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1390 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750]}), .c ({signal_4279, signal_4278, signal_4277, signal_4276, signal_1405}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1391 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_3047, signal_3046, signal_3045, signal_3044, signal_1097}), .clk ( clk ), .r ({Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_4283, signal_4282, signal_4281, signal_4280, signal_1406}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1392 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770]}), .c ({signal_4287, signal_4286, signal_4285, signal_4284, signal_1407}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1393 ( .a ({signal_17517, signal_17515, signal_17513, signal_17511, signal_17509}), .b ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .c ({signal_4291, signal_4290, signal_4289, signal_4288, signal_1408}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1394 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_3115, signal_3114, signal_3113, signal_3112, signal_1114}), .clk ( clk ), .r ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_4295, signal_4294, signal_4293, signal_4292, signal_1409}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1397 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_3067, signal_3066, signal_3065, signal_3064, signal_1102}), .clk ( clk ), .r ({Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .c ({signal_4307, signal_4306, signal_4305, signal_4304, signal_1412}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1398 ( .a ({signal_17357, signal_17355, signal_17353, signal_17351, signal_17349}), .b ({signal_3151, signal_3150, signal_3149, signal_3148, signal_1123}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810]}), .c ({signal_4311, signal_4310, signal_4309, signal_4308, signal_1413}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1399 ( .a ({signal_17527, signal_17525, signal_17523, signal_17521, signal_17519}), .b ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .clk ( clk ), .r ({Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_4315, signal_4314, signal_4313, signal_4312, signal_1414}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1400 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .clk ( clk ), .r ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830]}), .c ({signal_4319, signal_4318, signal_4317, signal_4316, signal_1415}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1404 ( .a ({signal_17417, signal_17415, signal_17413, signal_17411, signal_17409}), .b ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1078}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .c ({signal_4335, signal_4334, signal_4333, signal_4332, signal_1419}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1405 ( .a ({signal_17307, signal_17305, signal_17303, signal_17301, signal_17299}), .b ({signal_3067, signal_3066, signal_3065, signal_3064, signal_1102}), .clk ( clk ), .r ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_4339, signal_4338, signal_4337, signal_4336, signal_1420}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1406 ( .a ({signal_17537, signal_17535, signal_17533, signal_17531, signal_17529}), .b ({signal_3119, signal_3118, signal_3117, signal_3116, signal_1115}), .clk ( clk ), .r ({Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .c ({signal_4343, signal_4342, signal_4341, signal_4340, signal_1421}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1409 ( .a ({signal_17547, signal_17545, signal_17543, signal_17541, signal_17539}), .b ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870]}), .c ({signal_4355, signal_4354, signal_4353, signal_4352, signal_1424}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1410 ( .a ({signal_17237, signal_17235, signal_17233, signal_17231, signal_17229}), .b ({signal_3087, signal_3086, signal_3085, signal_3084, signal_1107}), .clk ( clk ), .r ({Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_4359, signal_4358, signal_4357, signal_4356, signal_1425}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1411 ( .a ({signal_17417, signal_17415, signal_17413, signal_17411, signal_17409}), .b ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}), .clk ( clk ), .r ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890]}), .c ({signal_4363, signal_4362, signal_4361, signal_4360, signal_1426}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1412 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_3171, signal_3170, signal_3169, signal_3168, signal_1128}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .c ({signal_4367, signal_4366, signal_4365, signal_4364, signal_1427}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1413 ( .a ({signal_17557, signal_17555, signal_17553, signal_17551, signal_17549}), .b ({signal_2947, signal_2946, signal_2945, signal_2944, signal_1072}), .clk ( clk ), .r ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_4371, signal_4370, signal_4369, signal_4368, signal_1428}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1414 ( .a ({signal_17567, signal_17565, signal_17563, signal_17561, signal_17559}), .b ({signal_3191, signal_3190, signal_3189, signal_3188, signal_1133}), .clk ( clk ), .r ({Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .c ({signal_4375, signal_4374, signal_4373, signal_4372, signal_1429}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1415 ( .a ({signal_17407, signal_17405, signal_17403, signal_17401, signal_17399}), .b ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930]}), .c ({signal_4379, signal_4378, signal_4377, signal_4376, signal_1430}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1416 ( .a ({signal_17587, signal_17583, signal_17579, signal_17575, signal_17571}), .b ({signal_3211, signal_3210, signal_3209, signal_3208, signal_1138}), .clk ( clk ), .r ({Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_4383, signal_4382, signal_4381, signal_4380, signal_1431}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1417 ( .a ({signal_17357, signal_17355, signal_17353, signal_17351, signal_17349}), .b ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .clk ( clk ), .r ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950]}), .c ({signal_4387, signal_4386, signal_4385, signal_4384, signal_1432}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1418 ( .a ({signal_17597, signal_17595, signal_17593, signal_17591, signal_17589}), .b ({signal_3219, signal_3218, signal_3217, signal_3216, signal_1140}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .c ({signal_4391, signal_4390, signal_4389, signal_4388, signal_1433}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1419 ( .a ({signal_17607, signal_17605, signal_17603, signal_17601, signal_17599}), .b ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .clk ( clk ), .r ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_4395, signal_4394, signal_4393, signal_4392, signal_1434}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1420 ( .a ({signal_17377, signal_17375, signal_17373, signal_17371, signal_17369}), .b ({signal_3227, signal_3226, signal_3225, signal_3224, signal_1142}), .clk ( clk ), .r ({Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .c ({signal_4399, signal_4398, signal_4397, signal_4396, signal_1435}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1421 ( .a ({signal_17527, signal_17525, signal_17523, signal_17521, signal_17519}), .b ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990]}), .c ({signal_4403, signal_4402, signal_4401, signal_4400, signal_1436}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1422 ( .a ({signal_17377, signal_17375, signal_17373, signal_17371, signal_17369}), .b ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .clk ( clk ), .r ({Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_4407, signal_4406, signal_4405, signal_4404, signal_1437}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1423 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3263, signal_3262, signal_3261, signal_3260, signal_1151}), .clk ( clk ), .r ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010]}), .c ({signal_4411, signal_4410, signal_4409, signal_4408, signal_1438}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1424 ( .a ({signal_17617, signal_17615, signal_17613, signal_17611, signal_17609}), .b ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .c ({signal_4415, signal_4414, signal_4413, signal_4412, signal_1439}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1425 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_3283, signal_3282, signal_3281, signal_3280, signal_1156}), .clk ( clk ), .r ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_4419, signal_4418, signal_4417, signal_4416, signal_1440}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1426 ( .a ({signal_17437, signal_17435, signal_17433, signal_17431, signal_17429}), .b ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}), .clk ( clk ), .r ({Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .c ({signal_4423, signal_4422, signal_4421, signal_4420, signal_1441}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1427 ( .a ({signal_17377, signal_17375, signal_17373, signal_17371, signal_17369}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050]}), .c ({signal_4427, signal_4426, signal_4425, signal_4424, signal_1442}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1428 ( .a ({signal_17537, signal_17535, signal_17533, signal_17531, signal_17529}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_4431, signal_4430, signal_4429, signal_4428, signal_1443}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1429 ( .a ({signal_17367, signal_17365, signal_17363, signal_17361, signal_17359}), .b ({signal_3323, signal_3322, signal_3321, signal_3320, signal_1166}), .clk ( clk ), .r ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070]}), .c ({signal_4435, signal_4434, signal_4433, signal_4432, signal_1444}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1430 ( .a ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}), .b ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .c ({signal_4439, signal_4438, signal_4437, signal_4436, signal_1445}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1431 ( .a ({signal_17627, signal_17625, signal_17623, signal_17621, signal_17619}), .b ({signal_3331, signal_3330, signal_3329, signal_3328, signal_1168}), .clk ( clk ), .r ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_4443, signal_4442, signal_4441, signal_4440, signal_1446}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1432 ( .a ({signal_2747, signal_2746, signal_2745, signal_2744, signal_1022}), .b ({signal_3227, signal_3226, signal_3225, signal_3224, signal_1142}), .clk ( clk ), .r ({Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .c ({signal_4447, signal_4446, signal_4445, signal_4444, signal_1447}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1433 ( .a ({signal_17287, signal_17285, signal_17283, signal_17281, signal_17279}), .b ({signal_3203, signal_3202, signal_3201, signal_3200, signal_1136}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110]}), .c ({signal_4451, signal_4450, signal_4449, signal_4448, signal_1448}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1434 ( .a ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .b ({signal_3239, signal_3238, signal_3237, signal_3236, signal_1145}), .clk ( clk ), .r ({Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_4455, signal_4454, signal_4453, signal_4452, signal_1449}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1435 ( .a ({signal_17467, signal_17465, signal_17463, signal_17461, signal_17459}), .b ({signal_3323, signal_3322, signal_3321, signal_3320, signal_1166}), .clk ( clk ), .r ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130]}), .c ({signal_4459, signal_4458, signal_4457, signal_4456, signal_1450}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1436 ( .a ({signal_17637, signal_17635, signal_17633, signal_17631, signal_17629}), .b ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .c ({signal_4463, signal_4462, signal_4461, signal_4460, signal_1451}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1437 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_3363, signal_3362, signal_3361, signal_3360, signal_1176}), .clk ( clk ), .r ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_4467, signal_4466, signal_4465, signal_4464, signal_1452}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1438 ( .a ({signal_3203, signal_3202, signal_3201, signal_3200, signal_1136}), .b ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .clk ( clk ), .r ({Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .c ({signal_4471, signal_4470, signal_4469, signal_4468, signal_1453}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1439 ( .a ({signal_3023, signal_3022, signal_3021, signal_3020, signal_1091}), .b ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170]}), .c ({signal_4475, signal_4474, signal_4473, signal_4472, signal_1454}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1440 ( .a ({signal_17337, signal_17335, signal_17333, signal_17331, signal_17329}), .b ({signal_3287, signal_3286, signal_3285, signal_3284, signal_1157}), .clk ( clk ), .r ({Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_4479, signal_4478, signal_4477, signal_4476, signal_1455}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1441 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_3371, signal_3370, signal_3369, signal_3368, signal_1178}), .clk ( clk ), .r ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190]}), .c ({signal_4483, signal_4482, signal_4481, signal_4480, signal_1456}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1442 ( .a ({signal_17547, signal_17545, signal_17543, signal_17541, signal_17539}), .b ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .c ({signal_4487, signal_4486, signal_4485, signal_4484, signal_1457}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1443 ( .a ({signal_17567, signal_17565, signal_17563, signal_17561, signal_17559}), .b ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}), .clk ( clk ), .r ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_4491, signal_4490, signal_4489, signal_4488, signal_1458}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1444 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .clk ( clk ), .r ({Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .c ({signal_4495, signal_4494, signal_4493, signal_4492, signal_1459}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1445 ( .a ({signal_17407, signal_17405, signal_17403, signal_17401, signal_17399}), .b ({signal_3415, signal_3414, signal_3413, signal_3412, signal_1189}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230]}), .c ({signal_4499, signal_4498, signal_4497, signal_4496, signal_1460}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1446 ( .a ({signal_17647, signal_17645, signal_17643, signal_17641, signal_17639}), .b ({signal_3419, signal_3418, signal_3417, signal_3416, signal_1190}), .clk ( clk ), .r ({Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_4503, signal_4502, signal_4501, signal_4500, signal_1461}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1447 ( .a ({signal_17407, signal_17405, signal_17403, signal_17401, signal_17399}), .b ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .clk ( clk ), .r ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250]}), .c ({signal_4507, signal_4506, signal_4505, signal_4504, signal_1462}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1448 ( .a ({signal_17657, signal_17655, signal_17653, signal_17651, signal_17649}), .b ({signal_3287, signal_3286, signal_3285, signal_3284, signal_1157}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .c ({signal_4511, signal_4510, signal_4509, signal_4508, signal_1463}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1449 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .clk ( clk ), .r ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_4515, signal_4514, signal_4513, signal_4512, signal_1464}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1450 ( .a ({signal_17617, signal_17615, signal_17613, signal_17611, signal_17609}), .b ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}), .clk ( clk ), .r ({Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .c ({signal_4519, signal_4518, signal_4517, signal_4516, signal_1465}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1451 ( .a ({signal_17667, signal_17665, signal_17663, signal_17661, signal_17659}), .b ({signal_3451, signal_3450, signal_3449, signal_3448, signal_1198}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290]}), .c ({signal_4523, signal_4522, signal_4521, signal_4520, signal_1466}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1452 ( .a ({signal_17677, signal_17675, signal_17673, signal_17671, signal_17669}), .b ({signal_3239, signal_3238, signal_3237, signal_3236, signal_1145}), .clk ( clk ), .r ({Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_4527, signal_4526, signal_4525, signal_4524, signal_1467}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1453 ( .a ({signal_17687, signal_17685, signal_17683, signal_17681, signal_17679}), .b ({signal_3427, signal_3426, signal_3425, signal_3424, signal_1192}), .clk ( clk ), .r ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310]}), .c ({signal_4531, signal_4530, signal_4529, signal_4528, signal_1468}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1454 ( .a ({signal_3067, signal_3066, signal_3065, signal_3064, signal_1102}), .b ({signal_3291, signal_3290, signal_3289, signal_3288, signal_1158}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .c ({signal_4535, signal_4534, signal_4533, signal_4532, signal_1469}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1455 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_3367, signal_3366, signal_3365, signal_3364, signal_1177}), .clk ( clk ), .r ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_4539, signal_4538, signal_4537, signal_4536, signal_1470}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1456 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}), .clk ( clk ), .r ({Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .c ({signal_4543, signal_4542, signal_4541, signal_4540, signal_1471}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1457 ( .a ({signal_17537, signal_17535, signal_17533, signal_17531, signal_17529}), .b ({signal_3423, signal_3422, signal_3421, signal_3420, signal_1191}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350]}), .c ({signal_4547, signal_4546, signal_4545, signal_4544, signal_1472}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1458 ( .a ({signal_17457, signal_17455, signal_17453, signal_17451, signal_17449}), .b ({signal_3235, signal_3234, signal_3233, signal_3232, signal_1144}), .clk ( clk ), .r ({Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_4551, signal_4550, signal_4549, signal_4548, signal_1473}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1459 ( .a ({signal_17407, signal_17405, signal_17403, signal_17401, signal_17399}), .b ({signal_3367, signal_3366, signal_3365, signal_3364, signal_1177}), .clk ( clk ), .r ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370]}), .c ({signal_4555, signal_4554, signal_4553, signal_4552, signal_1474}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1460 ( .a ({signal_17507, signal_17505, signal_17503, signal_17501, signal_17499}), .b ({signal_3403, signal_3402, signal_3401, signal_3400, signal_1186}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .c ({signal_4559, signal_4558, signal_4557, signal_4556, signal_1475}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1461 ( .a ({signal_17417, signal_17415, signal_17413, signal_17411, signal_17409}), .b ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}), .clk ( clk ), .r ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_4563, signal_4562, signal_4561, signal_4560, signal_1476}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1462 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}), .clk ( clk ), .r ({Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .c ({signal_4567, signal_4566, signal_4565, signal_4564, signal_1477}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1463 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3483, signal_3482, signal_3481, signal_3480, signal_1206}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410]}), .c ({signal_4571, signal_4570, signal_4569, signal_4568, signal_1478}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1464 ( .a ({signal_17567, signal_17565, signal_17563, signal_17561, signal_17559}), .b ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .clk ( clk ), .r ({Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_4575, signal_4574, signal_4573, signal_4572, signal_1479}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1465 ( .a ({signal_17277, signal_17275, signal_17273, signal_17271, signal_17269}), .b ({signal_3403, signal_3402, signal_3401, signal_3400, signal_1186}), .clk ( clk ), .r ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430]}), .c ({signal_4579, signal_4578, signal_4577, signal_4576, signal_1480}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1466 ( .a ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1075}), .b ({signal_2983, signal_2982, signal_2981, signal_2980, signal_1081}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .c ({signal_4583, signal_4582, signal_4581, signal_4580, signal_1481}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1467 ( .a ({signal_17317, signal_17315, signal_17313, signal_17311, signal_17309}), .b ({signal_3331, signal_3330, signal_3329, signal_3328, signal_1168}), .clk ( clk ), .r ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_4587, signal_4586, signal_4585, signal_4584, signal_1482}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1468 ( .a ({signal_17537, signal_17535, signal_17533, signal_17531, signal_17529}), .b ({signal_3303, signal_3302, signal_3301, signal_3300, signal_1161}), .clk ( clk ), .r ({Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .c ({signal_4591, signal_4590, signal_4589, signal_4588, signal_1483}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1469 ( .a ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1021}), .b ({signal_3187, signal_3186, signal_3185, signal_3184, signal_1132}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470]}), .c ({signal_4595, signal_4594, signal_4593, signal_4592, signal_1484}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1470 ( .a ({signal_17487, signal_17485, signal_17483, signal_17481, signal_17479}), .b ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}), .clk ( clk ), .r ({Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_4599, signal_4598, signal_4597, signal_4596, signal_1485}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1471 ( .a ({signal_17697, signal_17695, signal_17693, signal_17691, signal_17689}), .b ({signal_3491, signal_3490, signal_3489, signal_3488, signal_1208}), .clk ( clk ), .r ({Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490]}), .c ({signal_4603, signal_4602, signal_4601, signal_4600, signal_1486}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1472 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_2995, signal_2994, signal_2993, signal_2992, signal_1084}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500]}), .c ({signal_4607, signal_4606, signal_4605, signal_4604, signal_1487}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1473 ( .a ({signal_17457, signal_17455, signal_17453, signal_17451, signal_17449}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_4611, signal_4610, signal_4609, signal_4608, signal_1488}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1474 ( .a ({signal_17707, signal_17705, signal_17703, signal_17701, signal_17699}), .b ({signal_3463, signal_3462, signal_3461, signal_3460, signal_1201}), .clk ( clk ), .r ({Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520]}), .c ({signal_4615, signal_4614, signal_4613, signal_4612, signal_1489}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1475 ( .a ({signal_17307, signal_17305, signal_17303, signal_17301, signal_17299}), .b ({signal_3303, signal_3302, signal_3301, signal_3300, signal_1161}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530]}), .c ({signal_4619, signal_4618, signal_4617, signal_4616, signal_1490}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1476 ( .a ({signal_17227, signal_17223, signal_17219, signal_17215, signal_17211}), .b ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .clk ( clk ), .r ({Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_4623, signal_4622, signal_4621, signal_4620, signal_1491}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1477 ( .a ({signal_17567, signal_17565, signal_17563, signal_17561, signal_17559}), .b ({signal_3527, signal_3526, signal_3525, signal_3524, signal_1217}), .clk ( clk ), .r ({Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550]}), .c ({signal_4627, signal_4626, signal_4625, signal_4624, signal_1492}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1478 ( .a ({signal_17557, signal_17555, signal_17553, signal_17551, signal_17549}), .b ({signal_3039, signal_3038, signal_3037, signal_3036, signal_1095}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560]}), .c ({signal_4631, signal_4630, signal_4629, signal_4628, signal_1493}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1479 ( .a ({signal_17227, signal_17223, signal_17219, signal_17215, signal_17211}), .b ({signal_3415, signal_3414, signal_3413, signal_3412, signal_1189}), .clk ( clk ), .r ({Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_4635, signal_4634, signal_4633, signal_4632, signal_1494}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1480 ( .a ({signal_17717, signal_17715, signal_17713, signal_17711, signal_17709}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580]}), .c ({signal_4639, signal_4638, signal_4637, signal_4636, signal_1495}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1481 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1073}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590]}), .c ({signal_4643, signal_4642, signal_4641, signal_4640, signal_1496}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1482 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3235, signal_3234, signal_3233, signal_3232, signal_1144}), .clk ( clk ), .r ({Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_4647, signal_4646, signal_4645, signal_4644, signal_1497}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1483 ( .a ({signal_17417, signal_17415, signal_17413, signal_17411, signal_17409}), .b ({signal_3235, signal_3234, signal_3233, signal_3232, signal_1144}), .clk ( clk ), .r ({Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610]}), .c ({signal_4651, signal_4650, signal_4649, signal_4648, signal_1498}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1484 ( .a ({signal_17357, signal_17355, signal_17353, signal_17351, signal_17349}), .b ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620]}), .c ({signal_4655, signal_4654, signal_4653, signal_4652, signal_1499}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1485 ( .a ({signal_17227, signal_17223, signal_17219, signal_17215, signal_17211}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_4659, signal_4658, signal_4657, signal_4656, signal_1500}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1486 ( .a ({signal_17547, signal_17545, signal_17543, signal_17541, signal_17539}), .b ({signal_3307, signal_3306, signal_3305, signal_3304, signal_1162}), .clk ( clk ), .r ({Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640]}), .c ({signal_4663, signal_4662, signal_4661, signal_4660, signal_1501}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1487 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650]}), .c ({signal_4667, signal_4666, signal_4665, signal_4664, signal_1502}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1488 ( .a ({signal_17427, signal_17425, signal_17423, signal_17421, signal_17419}), .b ({signal_3231, signal_3230, signal_3229, signal_3228, signal_1143}), .clk ( clk ), .r ({Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_4671, signal_4670, signal_4669, signal_4668, signal_1503}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1489 ( .a ({signal_17367, signal_17365, signal_17363, signal_17361, signal_17359}), .b ({signal_3135, signal_3134, signal_3133, signal_3132, signal_1119}), .clk ( clk ), .r ({Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670]}), .c ({signal_4675, signal_4674, signal_4673, signal_4672, signal_1504}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1490 ( .a ({signal_4123, signal_4122, signal_4121, signal_4120, signal_1366}), .b ({signal_4679, signal_4678, signal_4677, signal_4676, signal_1505}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1491 ( .a ({signal_4127, signal_4126, signal_4125, signal_4124, signal_1367}), .b ({signal_4683, signal_4682, signal_4681, signal_4680, signal_1506}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1497 ( .a ({signal_4151, signal_4150, signal_4149, signal_4148, signal_1373}), .b ({signal_4707, signal_4706, signal_4705, signal_4704, signal_1512}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1498 ( .a ({signal_4155, signal_4154, signal_4153, signal_4152, signal_1374}), .b ({signal_4711, signal_4710, signal_4709, signal_4708, signal_1513}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1502 ( .a ({signal_4171, signal_4170, signal_4169, signal_4168, signal_1378}), .b ({signal_4727, signal_4726, signal_4725, signal_4724, signal_1517}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1503 ( .a ({signal_4175, signal_4174, signal_4173, signal_4172, signal_1379}), .b ({signal_4731, signal_4730, signal_4729, signal_4728, signal_1518}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1508 ( .a ({signal_4199, signal_4198, signal_4197, signal_4196, signal_1385}), .b ({signal_4751, signal_4750, signal_4749, signal_4748, signal_1523}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1509 ( .a ({signal_4203, signal_4202, signal_4201, signal_4200, signal_1386}), .b ({signal_4755, signal_4754, signal_4753, signal_4752, signal_1524}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1510 ( .a ({signal_4207, signal_4206, signal_4205, signal_4204, signal_1387}), .b ({signal_4759, signal_4758, signal_4757, signal_4756, signal_1525}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1511 ( .a ({signal_4211, signal_4210, signal_4209, signal_4208, signal_1388}), .b ({signal_4763, signal_4762, signal_4761, signal_4760, signal_1526}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1512 ( .a ({signal_4215, signal_4214, signal_4213, signal_4212, signal_1389}), .b ({signal_4767, signal_4766, signal_4765, signal_4764, signal_1527}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1514 ( .a ({signal_4227, signal_4226, signal_4225, signal_4224, signal_1392}), .b ({signal_4775, signal_4774, signal_4773, signal_4772, signal_1529}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1515 ( .a ({signal_4231, signal_4230, signal_4229, signal_4228, signal_1393}), .b ({signal_4779, signal_4778, signal_4777, signal_4776, signal_1530}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1516 ( .a ({signal_4235, signal_4234, signal_4233, signal_4232, signal_1394}), .b ({signal_4783, signal_4782, signal_4781, signal_4780, signal_1531}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1517 ( .a ({signal_4239, signal_4238, signal_4237, signal_4236, signal_1395}), .b ({signal_4787, signal_4786, signal_4785, signal_4784, signal_1532}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1518 ( .a ({signal_4243, signal_4242, signal_4241, signal_4240, signal_1396}), .b ({signal_4791, signal_4790, signal_4789, signal_4788, signal_1533}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1519 ( .a ({signal_4247, signal_4246, signal_4245, signal_4244, signal_1397}), .b ({signal_4795, signal_4794, signal_4793, signal_4792, signal_1534}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1521 ( .a ({signal_4255, signal_4254, signal_4253, signal_4252, signal_1399}), .b ({signal_4803, signal_4802, signal_4801, signal_4800, signal_1536}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1522 ( .a ({signal_4259, signal_4258, signal_4257, signal_4256, signal_1400}), .b ({signal_4807, signal_4806, signal_4805, signal_4804, signal_1537}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1523 ( .a ({signal_4263, signal_4262, signal_4261, signal_4260, signal_1401}), .b ({signal_4811, signal_4810, signal_4809, signal_4808, signal_1538}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1524 ( .a ({signal_4267, signal_4266, signal_4265, signal_4264, signal_1402}), .b ({signal_4815, signal_4814, signal_4813, signal_4812, signal_1539}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1525 ( .a ({signal_4271, signal_4270, signal_4269, signal_4268, signal_1403}), .b ({signal_4819, signal_4818, signal_4817, signal_4816, signal_1540}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1526 ( .a ({signal_4275, signal_4274, signal_4273, signal_4272, signal_1404}), .b ({signal_4823, signal_4822, signal_4821, signal_4820, signal_1541}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1527 ( .a ({signal_4279, signal_4278, signal_4277, signal_4276, signal_1405}), .b ({signal_4827, signal_4826, signal_4825, signal_4824, signal_1542}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1528 ( .a ({signal_4283, signal_4282, signal_4281, signal_4280, signal_1406}), .b ({signal_4831, signal_4830, signal_4829, signal_4828, signal_1543}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1529 ( .a ({signal_4287, signal_4286, signal_4285, signal_4284, signal_1407}), .b ({signal_4835, signal_4834, signal_4833, signal_4832, signal_1544}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1530 ( .a ({signal_4291, signal_4290, signal_4289, signal_4288, signal_1408}), .b ({signal_4839, signal_4838, signal_4837, signal_4836, signal_1545}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1531 ( .a ({signal_4295, signal_4294, signal_4293, signal_4292, signal_1409}), .b ({signal_4843, signal_4842, signal_4841, signal_4840, signal_1546}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1534 ( .a ({signal_4307, signal_4306, signal_4305, signal_4304, signal_1412}), .b ({signal_4855, signal_4854, signal_4853, signal_4852, signal_1549}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1535 ( .a ({signal_4311, signal_4310, signal_4309, signal_4308, signal_1413}), .b ({signal_4859, signal_4858, signal_4857, signal_4856, signal_1550}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1536 ( .a ({signal_4315, signal_4314, signal_4313, signal_4312, signal_1414}), .b ({signal_4863, signal_4862, signal_4861, signal_4860, signal_1551}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1537 ( .a ({signal_4319, signal_4318, signal_4317, signal_4316, signal_1415}), .b ({signal_4867, signal_4866, signal_4865, signal_4864, signal_1552}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1540 ( .a ({signal_4335, signal_4334, signal_4333, signal_4332, signal_1419}), .b ({signal_4879, signal_4878, signal_4877, signal_4876, signal_1555}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1541 ( .a ({signal_4339, signal_4338, signal_4337, signal_4336, signal_1420}), .b ({signal_4883, signal_4882, signal_4881, signal_4880, signal_1556}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1542 ( .a ({signal_4343, signal_4342, signal_4341, signal_4340, signal_1421}), .b ({signal_4887, signal_4886, signal_4885, signal_4884, signal_1557}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1545 ( .a ({signal_4355, signal_4354, signal_4353, signal_4352, signal_1424}), .b ({signal_4899, signal_4898, signal_4897, signal_4896, signal_1560}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1546 ( .a ({signal_4359, signal_4358, signal_4357, signal_4356, signal_1425}), .b ({signal_4903, signal_4902, signal_4901, signal_4900, signal_1561}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1547 ( .a ({signal_4363, signal_4362, signal_4361, signal_4360, signal_1426}), .b ({signal_4907, signal_4906, signal_4905, signal_4904, signal_1562}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1548 ( .a ({signal_4367, signal_4366, signal_4365, signal_4364, signal_1427}), .b ({signal_4911, signal_4910, signal_4909, signal_4908, signal_1563}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1549 ( .a ({signal_4371, signal_4370, signal_4369, signal_4368, signal_1428}), .b ({signal_4915, signal_4914, signal_4913, signal_4912, signal_1564}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1550 ( .a ({signal_4375, signal_4374, signal_4373, signal_4372, signal_1429}), .b ({signal_4919, signal_4918, signal_4917, signal_4916, signal_1565}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1551 ( .a ({signal_4379, signal_4378, signal_4377, signal_4376, signal_1430}), .b ({signal_4923, signal_4922, signal_4921, signal_4920, signal_1566}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1552 ( .a ({signal_4383, signal_4382, signal_4381, signal_4380, signal_1431}), .b ({signal_4927, signal_4926, signal_4925, signal_4924, signal_1567}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1553 ( .a ({signal_4387, signal_4386, signal_4385, signal_4384, signal_1432}), .b ({signal_4931, signal_4930, signal_4929, signal_4928, signal_1568}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1554 ( .a ({signal_4391, signal_4390, signal_4389, signal_4388, signal_1433}), .b ({signal_4935, signal_4934, signal_4933, signal_4932, signal_1569}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1555 ( .a ({signal_4395, signal_4394, signal_4393, signal_4392, signal_1434}), .b ({signal_4939, signal_4938, signal_4937, signal_4936, signal_1570}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1556 ( .a ({signal_4399, signal_4398, signal_4397, signal_4396, signal_1435}), .b ({signal_4943, signal_4942, signal_4941, signal_4940, signal_1571}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1557 ( .a ({signal_4403, signal_4402, signal_4401, signal_4400, signal_1436}), .b ({signal_4947, signal_4946, signal_4945, signal_4944, signal_1572}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1558 ( .a ({signal_4407, signal_4406, signal_4405, signal_4404, signal_1437}), .b ({signal_4951, signal_4950, signal_4949, signal_4948, signal_1573}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1559 ( .a ({signal_4411, signal_4410, signal_4409, signal_4408, signal_1438}), .b ({signal_4955, signal_4954, signal_4953, signal_4952, signal_1574}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1560 ( .a ({signal_4415, signal_4414, signal_4413, signal_4412, signal_1439}), .b ({signal_4959, signal_4958, signal_4957, signal_4956, signal_1575}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1561 ( .a ({signal_4419, signal_4418, signal_4417, signal_4416, signal_1440}), .b ({signal_4963, signal_4962, signal_4961, signal_4960, signal_1576}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1562 ( .a ({signal_4423, signal_4422, signal_4421, signal_4420, signal_1441}), .b ({signal_4967, signal_4966, signal_4965, signal_4964, signal_1577}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1563 ( .a ({signal_4427, signal_4426, signal_4425, signal_4424, signal_1442}), .b ({signal_4971, signal_4970, signal_4969, signal_4968, signal_1578}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1564 ( .a ({signal_4431, signal_4430, signal_4429, signal_4428, signal_1443}), .b ({signal_4975, signal_4974, signal_4973, signal_4972, signal_1579}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1565 ( .a ({signal_4435, signal_4434, signal_4433, signal_4432, signal_1444}), .b ({signal_4979, signal_4978, signal_4977, signal_4976, signal_1580}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1566 ( .a ({signal_4439, signal_4438, signal_4437, signal_4436, signal_1445}), .b ({signal_4983, signal_4982, signal_4981, signal_4980, signal_1581}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1567 ( .a ({signal_4447, signal_4446, signal_4445, signal_4444, signal_1447}), .b ({signal_4987, signal_4986, signal_4985, signal_4984, signal_1582}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1568 ( .a ({signal_4451, signal_4450, signal_4449, signal_4448, signal_1448}), .b ({signal_4991, signal_4990, signal_4989, signal_4988, signal_1583}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1569 ( .a ({signal_4455, signal_4454, signal_4453, signal_4452, signal_1449}), .b ({signal_4995, signal_4994, signal_4993, signal_4992, signal_1584}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1570 ( .a ({signal_4459, signal_4458, signal_4457, signal_4456, signal_1450}), .b ({signal_4999, signal_4998, signal_4997, signal_4996, signal_1585}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1571 ( .a ({signal_4463, signal_4462, signal_4461, signal_4460, signal_1451}), .b ({signal_5003, signal_5002, signal_5001, signal_5000, signal_1586}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1572 ( .a ({signal_4467, signal_4466, signal_4465, signal_4464, signal_1452}), .b ({signal_5007, signal_5006, signal_5005, signal_5004, signal_1587}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1573 ( .a ({signal_4471, signal_4470, signal_4469, signal_4468, signal_1453}), .b ({signal_5011, signal_5010, signal_5009, signal_5008, signal_1588}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1574 ( .a ({signal_4475, signal_4474, signal_4473, signal_4472, signal_1454}), .b ({signal_5015, signal_5014, signal_5013, signal_5012, signal_1589}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1575 ( .a ({signal_4479, signal_4478, signal_4477, signal_4476, signal_1455}), .b ({signal_5019, signal_5018, signal_5017, signal_5016, signal_1590}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1576 ( .a ({signal_4483, signal_4482, signal_4481, signal_4480, signal_1456}), .b ({signal_5023, signal_5022, signal_5021, signal_5020, signal_1591}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1577 ( .a ({signal_4487, signal_4486, signal_4485, signal_4484, signal_1457}), .b ({signal_5027, signal_5026, signal_5025, signal_5024, signal_1592}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1578 ( .a ({signal_4491, signal_4490, signal_4489, signal_4488, signal_1458}), .b ({signal_5031, signal_5030, signal_5029, signal_5028, signal_1593}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1579 ( .a ({signal_4495, signal_4494, signal_4493, signal_4492, signal_1459}), .b ({signal_5035, signal_5034, signal_5033, signal_5032, signal_1594}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1580 ( .a ({signal_4499, signal_4498, signal_4497, signal_4496, signal_1460}), .b ({signal_5039, signal_5038, signal_5037, signal_5036, signal_1595}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1581 ( .a ({signal_4507, signal_4506, signal_4505, signal_4504, signal_1462}), .b ({signal_5043, signal_5042, signal_5041, signal_5040, signal_1596}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1582 ( .a ({signal_4511, signal_4510, signal_4509, signal_4508, signal_1463}), .b ({signal_5047, signal_5046, signal_5045, signal_5044, signal_1597}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1583 ( .a ({signal_4515, signal_4514, signal_4513, signal_4512, signal_1464}), .b ({signal_5051, signal_5050, signal_5049, signal_5048, signal_1598}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1584 ( .a ({signal_4519, signal_4518, signal_4517, signal_4516, signal_1465}), .b ({signal_5055, signal_5054, signal_5053, signal_5052, signal_1599}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1585 ( .a ({signal_4523, signal_4522, signal_4521, signal_4520, signal_1466}), .b ({signal_5059, signal_5058, signal_5057, signal_5056, signal_1600}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1586 ( .a ({signal_4527, signal_4526, signal_4525, signal_4524, signal_1467}), .b ({signal_5063, signal_5062, signal_5061, signal_5060, signal_1601}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1587 ( .a ({signal_4531, signal_4530, signal_4529, signal_4528, signal_1468}), .b ({signal_5067, signal_5066, signal_5065, signal_5064, signal_1602}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1588 ( .a ({signal_4535, signal_4534, signal_4533, signal_4532, signal_1469}), .b ({signal_5071, signal_5070, signal_5069, signal_5068, signal_1603}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1589 ( .a ({signal_4539, signal_4538, signal_4537, signal_4536, signal_1470}), .b ({signal_5075, signal_5074, signal_5073, signal_5072, signal_1604}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1590 ( .a ({signal_4543, signal_4542, signal_4541, signal_4540, signal_1471}), .b ({signal_5079, signal_5078, signal_5077, signal_5076, signal_1605}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1591 ( .a ({signal_4547, signal_4546, signal_4545, signal_4544, signal_1472}), .b ({signal_5083, signal_5082, signal_5081, signal_5080, signal_1606}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1592 ( .a ({signal_4551, signal_4550, signal_4549, signal_4548, signal_1473}), .b ({signal_5087, signal_5086, signal_5085, signal_5084, signal_1607}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1593 ( .a ({signal_4555, signal_4554, signal_4553, signal_4552, signal_1474}), .b ({signal_5091, signal_5090, signal_5089, signal_5088, signal_1608}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1594 ( .a ({signal_4559, signal_4558, signal_4557, signal_4556, signal_1475}), .b ({signal_5095, signal_5094, signal_5093, signal_5092, signal_1609}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1595 ( .a ({signal_4563, signal_4562, signal_4561, signal_4560, signal_1476}), .b ({signal_5099, signal_5098, signal_5097, signal_5096, signal_1610}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1596 ( .a ({signal_4567, signal_4566, signal_4565, signal_4564, signal_1477}), .b ({signal_5103, signal_5102, signal_5101, signal_5100, signal_1611}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1597 ( .a ({signal_4575, signal_4574, signal_4573, signal_4572, signal_1479}), .b ({signal_5107, signal_5106, signal_5105, signal_5104, signal_1612}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1598 ( .a ({signal_4579, signal_4578, signal_4577, signal_4576, signal_1480}), .b ({signal_5111, signal_5110, signal_5109, signal_5108, signal_1613}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1599 ( .a ({signal_4583, signal_4582, signal_4581, signal_4580, signal_1481}), .b ({signal_5115, signal_5114, signal_5113, signal_5112, signal_1614}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1600 ( .a ({signal_4587, signal_4586, signal_4585, signal_4584, signal_1482}), .b ({signal_5119, signal_5118, signal_5117, signal_5116, signal_1615}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1601 ( .a ({signal_4591, signal_4590, signal_4589, signal_4588, signal_1483}), .b ({signal_5123, signal_5122, signal_5121, signal_5120, signal_1616}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1602 ( .a ({signal_4595, signal_4594, signal_4593, signal_4592, signal_1484}), .b ({signal_5127, signal_5126, signal_5125, signal_5124, signal_1617}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1603 ( .a ({signal_4599, signal_4598, signal_4597, signal_4596, signal_1485}), .b ({signal_5131, signal_5130, signal_5129, signal_5128, signal_1618}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1604 ( .a ({signal_4603, signal_4602, signal_4601, signal_4600, signal_1486}), .b ({signal_5135, signal_5134, signal_5133, signal_5132, signal_1619}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1605 ( .a ({signal_4607, signal_4606, signal_4605, signal_4604, signal_1487}), .b ({signal_5139, signal_5138, signal_5137, signal_5136, signal_1620}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1606 ( .a ({signal_4611, signal_4610, signal_4609, signal_4608, signal_1488}), .b ({signal_5143, signal_5142, signal_5141, signal_5140, signal_1621}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1607 ( .a ({signal_4615, signal_4614, signal_4613, signal_4612, signal_1489}), .b ({signal_5147, signal_5146, signal_5145, signal_5144, signal_1622}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1608 ( .a ({signal_4619, signal_4618, signal_4617, signal_4616, signal_1490}), .b ({signal_5151, signal_5150, signal_5149, signal_5148, signal_1623}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1609 ( .a ({signal_4623, signal_4622, signal_4621, signal_4620, signal_1491}), .b ({signal_5155, signal_5154, signal_5153, signal_5152, signal_1624}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1610 ( .a ({signal_4627, signal_4626, signal_4625, signal_4624, signal_1492}), .b ({signal_5159, signal_5158, signal_5157, signal_5156, signal_1625}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1611 ( .a ({signal_4631, signal_4630, signal_4629, signal_4628, signal_1493}), .b ({signal_5163, signal_5162, signal_5161, signal_5160, signal_1626}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1612 ( .a ({signal_4635, signal_4634, signal_4633, signal_4632, signal_1494}), .b ({signal_5167, signal_5166, signal_5165, signal_5164, signal_1627}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1613 ( .a ({signal_4639, signal_4638, signal_4637, signal_4636, signal_1495}), .b ({signal_5171, signal_5170, signal_5169, signal_5168, signal_1628}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1614 ( .a ({signal_4643, signal_4642, signal_4641, signal_4640, signal_1496}), .b ({signal_5175, signal_5174, signal_5173, signal_5172, signal_1629}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1615 ( .a ({signal_4647, signal_4646, signal_4645, signal_4644, signal_1497}), .b ({signal_5179, signal_5178, signal_5177, signal_5176, signal_1630}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1616 ( .a ({signal_4651, signal_4650, signal_4649, signal_4648, signal_1498}), .b ({signal_5183, signal_5182, signal_5181, signal_5180, signal_1631}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1617 ( .a ({signal_4655, signal_4654, signal_4653, signal_4652, signal_1499}), .b ({signal_5187, signal_5186, signal_5185, signal_5184, signal_1632}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1618 ( .a ({signal_4659, signal_4658, signal_4657, signal_4656, signal_1500}), .b ({signal_5191, signal_5190, signal_5189, signal_5188, signal_1633}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1619 ( .a ({signal_4663, signal_4662, signal_4661, signal_4660, signal_1501}), .b ({signal_5195, signal_5194, signal_5193, signal_5192, signal_1634}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1620 ( .a ({signal_4667, signal_4666, signal_4665, signal_4664, signal_1502}), .b ({signal_5199, signal_5198, signal_5197, signal_5196, signal_1635}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1621 ( .a ({signal_4671, signal_4670, signal_4669, signal_4668, signal_1503}), .b ({signal_5203, signal_5202, signal_5201, signal_5200, signal_1636}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1622 ( .a ({signal_4675, signal_4674, signal_4673, signal_4672, signal_1504}), .b ({signal_5207, signal_5206, signal_5205, signal_5204, signal_1637}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1623 ( .a ({signal_17687, signal_17685, signal_17683, signal_17681, signal_17679}), .b ({signal_3579, signal_3578, signal_3577, signal_3576, signal_1230}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680]}), .c ({signal_5211, signal_5210, signal_5209, signal_5208, signal_1638}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1624 ( .a ({signal_17727, signal_17725, signal_17723, signal_17721, signal_17719}), .b ({signal_3583, signal_3582, signal_3581, signal_3580, signal_1231}), .clk ( clk ), .r ({Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_5215, signal_5214, signal_5213, signal_5212, signal_1639}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1625 ( .a ({signal_17547, signal_17545, signal_17543, signal_17541, signal_17539}), .b ({signal_3603, signal_3602, signal_3601, signal_3600, signal_1236}), .clk ( clk ), .r ({Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700]}), .c ({signal_5219, signal_5218, signal_5217, signal_5216, signal_1640}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1626 ( .a ({signal_3599, signal_3598, signal_3597, signal_3596, signal_1235}), .b ({signal_3683, signal_3682, signal_3681, signal_3680, signal_1256}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710]}), .c ({signal_5223, signal_5222, signal_5221, signal_5220, signal_1641}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1627 ( .a ({signal_17737, signal_17735, signal_17733, signal_17731, signal_17729}), .b ({signal_3687, signal_3686, signal_3685, signal_3684, signal_1257}), .clk ( clk ), .r ({Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_5227, signal_5226, signal_5225, signal_5224, signal_1642}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1628 ( .a ({signal_17707, signal_17705, signal_17703, signal_17701, signal_17699}), .b ({signal_3711, signal_3710, signal_3709, signal_3708, signal_1263}), .clk ( clk ), .r ({Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730]}), .c ({signal_5231, signal_5230, signal_5229, signal_5228, signal_1643}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1629 ( .a ({signal_3659, signal_3658, signal_3657, signal_3656, signal_1250}), .b ({signal_3671, signal_3670, signal_3669, signal_3668, signal_1253}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740]}), .c ({signal_5235, signal_5234, signal_5233, signal_5232, signal_1644}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1630 ( .a ({signal_3727, signal_3726, signal_3725, signal_3724, signal_1267}), .b ({signal_3731, signal_3730, signal_3729, signal_3728, signal_1268}), .clk ( clk ), .r ({Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_5239, signal_5238, signal_5237, signal_5236, signal_1645}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1631 ( .a ({signal_17747, signal_17745, signal_17743, signal_17741, signal_17739}), .b ({signal_3619, signal_3618, signal_3617, signal_3616, signal_1240}), .clk ( clk ), .r ({Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760]}), .c ({signal_5243, signal_5242, signal_5241, signal_5240, signal_1646}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1632 ( .a ({signal_3735, signal_3734, signal_3733, signal_3732, signal_1269}), .b ({signal_3739, signal_3738, signal_3737, signal_3736, signal_1270}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770]}), .c ({signal_5247, signal_5246, signal_5245, signal_5244, signal_1647}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1633 ( .a ({signal_3599, signal_3598, signal_3597, signal_3596, signal_1235}), .b ({signal_3679, signal_3678, signal_3677, signal_3676, signal_1255}), .clk ( clk ), .r ({Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_5251, signal_5250, signal_5249, signal_5248, signal_1648}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1634 ( .a ({signal_3751, signal_3750, signal_3749, signal_3748, signal_1273}), .b ({signal_3755, signal_3754, signal_3753, signal_3752, signal_1274}), .clk ( clk ), .r ({Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790]}), .c ({signal_5255, signal_5254, signal_5253, signal_5252, signal_1649}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1635 ( .a ({signal_2879, signal_2878, signal_2877, signal_2876, signal_1055}), .b ({signal_3675, signal_3674, signal_3673, signal_3672, signal_1254}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800]}), .c ({signal_5259, signal_5258, signal_5257, signal_5256, signal_1650}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1636 ( .a ({signal_17717, signal_17715, signal_17713, signal_17711, signal_17709}), .b ({signal_3623, signal_3622, signal_3621, signal_3620, signal_1241}), .clk ( clk ), .r ({Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_5263, signal_5262, signal_5261, signal_5260, signal_1651}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1637 ( .a ({signal_3603, signal_3602, signal_3601, signal_3600, signal_1236}), .b ({signal_2895, signal_2894, signal_2893, signal_2892, signal_1059}), .clk ( clk ), .r ({Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820]}), .c ({signal_5267, signal_5266, signal_5265, signal_5264, signal_1652}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1638 ( .a ({signal_3779, signal_3778, signal_3777, signal_3776, signal_1280}), .b ({signal_3783, signal_3782, signal_3781, signal_3780, signal_1281}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830]}), .c ({signal_5271, signal_5270, signal_5269, signal_5268, signal_1653}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1639 ( .a ({signal_3791, signal_3790, signal_3789, signal_3788, signal_1283}), .b ({signal_3795, signal_3794, signal_3793, signal_3792, signal_1284}), .clk ( clk ), .r ({Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_5275, signal_5274, signal_5273, signal_5272, signal_1654}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1640 ( .a ({signal_3591, signal_3590, signal_3589, signal_3588, signal_1233}), .b ({signal_3803, signal_3802, signal_3801, signal_3800, signal_1286}), .clk ( clk ), .r ({Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850]}), .c ({signal_5279, signal_5278, signal_5277, signal_5276, signal_1655}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1641 ( .a ({signal_3607, signal_3606, signal_3605, signal_3604, signal_1237}), .b ({signal_3811, signal_3810, signal_3809, signal_3808, signal_1288}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860]}), .c ({signal_5283, signal_5282, signal_5281, signal_5280, signal_1656}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1642 ( .a ({signal_2895, signal_2894, signal_2893, signal_2892, signal_1059}), .b ({signal_3611, signal_3610, signal_3609, signal_3608, signal_1238}), .clk ( clk ), .r ({Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_5287, signal_5286, signal_5285, signal_5284, signal_1657}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1643 ( .a ({signal_3627, signal_3626, signal_3625, signal_3624, signal_1242}), .b ({signal_3631, signal_3630, signal_3629, signal_3628, signal_1243}), .clk ( clk ), .r ({Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880]}), .c ({signal_5291, signal_5290, signal_5289, signal_5288, signal_1658}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1645 ( .a ({signal_3835, signal_3834, signal_3833, signal_3832, signal_1294}), .b ({signal_3839, signal_3838, signal_3837, signal_3836, signal_1295}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890]}), .c ({signal_5299, signal_5298, signal_5297, signal_5296, signal_1660}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1646 ( .a ({signal_3611, signal_3610, signal_3609, signal_3608, signal_1238}), .b ({signal_3867, signal_3866, signal_3865, signal_3864, signal_1302}), .clk ( clk ), .r ({Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_5303, signal_5302, signal_5301, signal_5300, signal_1661}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1647 ( .a ({signal_17757, signal_17755, signal_17753, signal_17751, signal_17749}), .b ({signal_3883, signal_3882, signal_3881, signal_3880, signal_1306}), .clk ( clk ), .r ({Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910]}), .c ({signal_5307, signal_5306, signal_5305, signal_5304, signal_1662}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1648 ( .a ({signal_3667, signal_3666, signal_3665, signal_3664, signal_1252}), .b ({signal_3899, signal_3898, signal_3897, signal_3896, signal_1310}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920]}), .c ({signal_5311, signal_5310, signal_5309, signal_5308, signal_1663}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1649 ( .a ({signal_17767, signal_17765, signal_17763, signal_17761, signal_17759}), .b ({signal_4191, signal_4190, signal_4189, signal_4188, signal_1383}), .clk ( clk ), .r ({Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_5315, signal_5314, signal_5313, signal_5312, signal_1664}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1650 ( .a ({signal_17227, signal_17223, signal_17219, signal_17215, signal_17211}), .b ({signal_3847, signal_3846, signal_3845, signal_3844, signal_1297}), .clk ( clk ), .r ({Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940]}), .c ({signal_5319, signal_5318, signal_5317, signal_5316, signal_1665}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1651 ( .a ({signal_3635, signal_3634, signal_3633, signal_3632, signal_1244}), .b ({signal_3903, signal_3902, signal_3901, signal_3900, signal_1311}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950]}), .c ({signal_5323, signal_5322, signal_5321, signal_5320, signal_1666}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1653 ( .a ({signal_4163, signal_4162, signal_4161, signal_4160, signal_1376}), .b ({signal_3927, signal_3926, signal_3925, signal_3924, signal_1317}), .clk ( clk ), .r ({Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_5331, signal_5330, signal_5329, signal_5328, signal_1668}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1654 ( .a ({signal_3599, signal_3598, signal_3597, signal_3596, signal_1235}), .b ({signal_3935, signal_3934, signal_3933, signal_3932, signal_1319}), .clk ( clk ), .r ({Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970]}), .c ({signal_5335, signal_5334, signal_5333, signal_5332, signal_1669}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1655 ( .a ({signal_4219, signal_4218, signal_4217, signal_4216, signal_1390}), .b ({signal_2919, signal_2918, signal_2917, signal_2916, signal_1065}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980]}), .c ({signal_5339, signal_5338, signal_5337, signal_5336, signal_1670}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1656 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_3939, signal_3938, signal_3937, signal_3936, signal_1320}), .clk ( clk ), .r ({Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_5343, signal_5342, signal_5341, signal_5340, signal_1671}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1657 ( .a ({signal_3699, signal_3698, signal_3697, signal_3696, signal_1260}), .b ({signal_3859, signal_3858, signal_3857, signal_3856, signal_1300}), .clk ( clk ), .r ({Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000]}), .c ({signal_5347, signal_5346, signal_5345, signal_5344, signal_1672}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1658 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_3943, signal_3942, signal_3941, signal_3940, signal_1321}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010]}), .c ({signal_5351, signal_5350, signal_5349, signal_5348, signal_1673}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1659 ( .a ({signal_3923, signal_3922, signal_3921, signal_3920, signal_1316}), .b ({signal_3947, signal_3946, signal_3945, signal_3944, signal_1322}), .clk ( clk ), .r ({Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_5355, signal_5354, signal_5353, signal_5352, signal_1674}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1660 ( .a ({signal_2911, signal_2910, signal_2909, signal_2908, signal_1063}), .b ({signal_3951, signal_3950, signal_3949, signal_3948, signal_1323}), .clk ( clk ), .r ({Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030]}), .c ({signal_5359, signal_5358, signal_5357, signal_5356, signal_1675}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1661 ( .a ({signal_3955, signal_3954, signal_3953, signal_3952, signal_1324}), .b ({signal_3959, signal_3958, signal_3957, signal_3956, signal_1325}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040]}), .c ({signal_5363, signal_5362, signal_5361, signal_5360, signal_1676}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1663 ( .a ({signal_3619, signal_3618, signal_3617, signal_3616, signal_1240}), .b ({signal_3847, signal_3846, signal_3845, signal_3844, signal_1297}), .clk ( clk ), .r ({Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_5371, signal_5370, signal_5369, signal_5368, signal_1678}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1664 ( .a ({signal_3715, signal_3714, signal_3713, signal_3712, signal_1264}), .b ({signal_3983, signal_3982, signal_3981, signal_3980, signal_1331}), .clk ( clk ), .r ({Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060]}), .c ({signal_5375, signal_5374, signal_5373, signal_5372, signal_1679}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1665 ( .a ({signal_3627, signal_3626, signal_3625, signal_3624, signal_1242}), .b ({signal_3987, signal_3986, signal_3985, signal_3984, signal_1332}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070]}), .c ({signal_5379, signal_5378, signal_5377, signal_5376, signal_1680}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1666 ( .a ({signal_3723, signal_3722, signal_3721, signal_3720, signal_1266}), .b ({signal_3995, signal_3994, signal_3993, signal_3992, signal_1334}), .clk ( clk ), .r ({Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_5383, signal_5382, signal_5381, signal_5380, signal_1681}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1667 ( .a ({signal_3847, signal_3846, signal_3845, signal_3844, signal_1297}), .b ({signal_4007, signal_4006, signal_4005, signal_4004, signal_1337}), .clk ( clk ), .r ({Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090]}), .c ({signal_5387, signal_5386, signal_5385, signal_5384, signal_1682}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1668 ( .a ({signal_3743, signal_3742, signal_3741, signal_3740, signal_1271}), .b ({signal_3983, signal_3982, signal_3981, signal_3980, signal_1331}), .clk ( clk ), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100]}), .c ({signal_5391, signal_5390, signal_5389, signal_5388, signal_1683}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1669 ( .a ({signal_17337, signal_17335, signal_17333, signal_17331, signal_17329}), .b ({signal_3939, signal_3938, signal_3937, signal_3936, signal_1320}), .clk ( clk ), .r ({Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({signal_5395, signal_5394, signal_5393, signal_5392, signal_1684}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1670 ( .a ({signal_3815, signal_3814, signal_3813, signal_3812, signal_1289}), .b ({signal_4019, signal_4018, signal_4017, signal_4016, signal_1340}), .clk ( clk ), .r ({Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120]}), .c ({signal_5399, signal_5398, signal_5397, signal_5396, signal_1685}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1671 ( .a ({signal_17777, signal_17775, signal_17773, signal_17771, signal_17769}), .b ({signal_4023, signal_4022, signal_4021, signal_4020, signal_1341}), .clk ( clk ), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130]}), .c ({signal_5403, signal_5402, signal_5401, signal_5400, signal_1686}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1673 ( .a ({signal_3763, signal_3762, signal_3761, signal_3760, signal_1276}), .b ({signal_3979, signal_3978, signal_3977, signal_3976, signal_1330}), .clk ( clk ), .r ({Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({signal_5411, signal_5410, signal_5409, signal_5408, signal_1688}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1674 ( .a ({signal_3931, signal_3930, signal_3929, signal_3928, signal_1318}), .b ({signal_4331, signal_4330, signal_4329, signal_4328, signal_1418}), .clk ( clk ), .r ({Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150]}), .c ({signal_5415, signal_5414, signal_5413, signal_5412, signal_1689}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1675 ( .a ({signal_3695, signal_3694, signal_3693, signal_3692, signal_1259}), .b ({signal_3955, signal_3954, signal_3953, signal_3952, signal_1324}), .clk ( clk ), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160]}), .c ({signal_5419, signal_5418, signal_5417, signal_5416, signal_1690}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1676 ( .a ({signal_3767, signal_3766, signal_3765, signal_3764, signal_1277}), .b ({signal_4043, signal_4042, signal_4041, signal_4040, signal_1346}), .clk ( clk ), .r ({Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({signal_5423, signal_5422, signal_5421, signal_5420, signal_1691}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1677 ( .a ({signal_4047, signal_4046, signal_4045, signal_4044, signal_1347}), .b ({signal_4051, signal_4050, signal_4049, signal_4048, signal_1348}), .clk ( clk ), .r ({Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180]}), .c ({signal_5427, signal_5426, signal_5425, signal_5424, signal_1692}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1678 ( .a ({signal_3659, signal_3658, signal_3657, signal_3656, signal_1250}), .b ({signal_4055, signal_4054, signal_4053, signal_4052, signal_1349}), .clk ( clk ), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190]}), .c ({signal_5431, signal_5430, signal_5429, signal_5428, signal_1693}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1679 ( .a ({signal_4063, signal_4062, signal_4061, signal_4060, signal_1351}), .b ({signal_4067, signal_4066, signal_4065, signal_4064, signal_1352}), .clk ( clk ), .r ({Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({signal_5435, signal_5434, signal_5433, signal_5432, signal_1694}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1680 ( .a ({signal_3599, signal_3598, signal_3597, signal_3596, signal_1235}), .b ({signal_3895, signal_3894, signal_3893, signal_3892, signal_1309}), .clk ( clk ), .r ({Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210]}), .c ({signal_5439, signal_5438, signal_5437, signal_5436, signal_1695}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1681 ( .a ({signal_4079, signal_4078, signal_4077, signal_4076, signal_1355}), .b ({signal_4083, signal_4082, signal_4081, signal_4080, signal_1356}), .clk ( clk ), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220]}), .c ({signal_5443, signal_5442, signal_5441, signal_5440, signal_1696}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1682 ( .a ({signal_3919, signal_3918, signal_3917, signal_3916, signal_1315}), .b ({signal_4087, signal_4086, signal_4085, signal_4084, signal_1357}), .clk ( clk ), .r ({Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({signal_5447, signal_5446, signal_5445, signal_5444, signal_1697}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1684 ( .a ({signal_3815, signal_3814, signal_3813, signal_3812, signal_1289}), .b ({signal_3819, signal_3818, signal_3817, signal_3816, signal_1290}), .clk ( clk ), .r ({Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240]}), .c ({signal_5455, signal_5454, signal_5453, signal_5452, signal_1699}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1687 ( .a ({signal_3631, signal_3630, signal_3629, signal_3628, signal_1243}), .b ({signal_3819, signal_3818, signal_3817, signal_3816, signal_1290}), .clk ( clk ), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250]}), .c ({signal_5467, signal_5466, signal_5465, signal_5464, signal_1702}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1693 ( .a ({signal_3819, signal_3818, signal_3817, signal_3816, signal_1290}), .b ({signal_3879, signal_3878, signal_3877, signal_3876, signal_1305}), .clk ( clk ), .r ({Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({signal_5491, signal_5490, signal_5489, signal_5488, signal_1708}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1698 ( .a ({signal_3831, signal_3830, signal_3829, signal_3828, signal_1293}), .b ({signal_4115, signal_4114, signal_4113, signal_4112, signal_1364}), .clk ( clk ), .r ({Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270]}), .c ({signal_5511, signal_5510, signal_5509, signal_5508, signal_1713}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1700 ( .a ({signal_5211, signal_5210, signal_5209, signal_5208, signal_1638}), .b ({signal_5519, signal_5518, signal_5517, signal_5516, signal_1715}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1701 ( .a ({signal_5215, signal_5214, signal_5213, signal_5212, signal_1639}), .b ({signal_5523, signal_5522, signal_5521, signal_5520, signal_1716}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1702 ( .a ({signal_5223, signal_5222, signal_5221, signal_5220, signal_1641}), .b ({signal_5527, signal_5526, signal_5525, signal_5524, signal_1717}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1703 ( .a ({signal_5227, signal_5226, signal_5225, signal_5224, signal_1642}), .b ({signal_5531, signal_5530, signal_5529, signal_5528, signal_1718}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1704 ( .a ({signal_5231, signal_5230, signal_5229, signal_5228, signal_1643}), .b ({signal_5535, signal_5534, signal_5533, signal_5532, signal_1719}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1705 ( .a ({signal_5235, signal_5234, signal_5233, signal_5232, signal_1644}), .b ({signal_5539, signal_5538, signal_5537, signal_5536, signal_1720}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1706 ( .a ({signal_5243, signal_5242, signal_5241, signal_5240, signal_1646}), .b ({signal_5543, signal_5542, signal_5541, signal_5540, signal_1721}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1707 ( .a ({signal_5247, signal_5246, signal_5245, signal_5244, signal_1647}), .b ({signal_5547, signal_5546, signal_5545, signal_5544, signal_1722}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1708 ( .a ({signal_5251, signal_5250, signal_5249, signal_5248, signal_1648}), .b ({signal_5551, signal_5550, signal_5549, signal_5548, signal_1723}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1709 ( .a ({signal_5259, signal_5258, signal_5257, signal_5256, signal_1650}), .b ({signal_5555, signal_5554, signal_5553, signal_5552, signal_1724}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1710 ( .a ({signal_5263, signal_5262, signal_5261, signal_5260, signal_1651}), .b ({signal_5559, signal_5558, signal_5557, signal_5556, signal_1725}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1711 ( .a ({signal_5267, signal_5266, signal_5265, signal_5264, signal_1652}), .b ({signal_5563, signal_5562, signal_5561, signal_5560, signal_1726}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1712 ( .a ({signal_5283, signal_5282, signal_5281, signal_5280, signal_1656}), .b ({signal_5567, signal_5566, signal_5565, signal_5564, signal_1727}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1713 ( .a ({signal_5287, signal_5286, signal_5285, signal_5284, signal_1657}), .b ({signal_5571, signal_5570, signal_5569, signal_5568, signal_1728}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1714 ( .a ({signal_5291, signal_5290, signal_5289, signal_5288, signal_1658}), .b ({signal_5575, signal_5574, signal_5573, signal_5572, signal_1729}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1716 ( .a ({signal_5307, signal_5306, signal_5305, signal_5304, signal_1662}), .b ({signal_5583, signal_5582, signal_5581, signal_5580, signal_1731}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1717 ( .a ({signal_5311, signal_5310, signal_5309, signal_5308, signal_1663}), .b ({signal_5587, signal_5586, signal_5585, signal_5584, signal_1732}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1718 ( .a ({signal_5315, signal_5314, signal_5313, signal_5312, signal_1664}), .b ({signal_5591, signal_5590, signal_5589, signal_5588, signal_1733}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1719 ( .a ({signal_5319, signal_5318, signal_5317, signal_5316, signal_1665}), .b ({signal_5595, signal_5594, signal_5593, signal_5592, signal_1734}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1720 ( .a ({signal_5323, signal_5322, signal_5321, signal_5320, signal_1666}), .b ({signal_5599, signal_5598, signal_5597, signal_5596, signal_1735}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1722 ( .a ({signal_5335, signal_5334, signal_5333, signal_5332, signal_1669}), .b ({signal_5607, signal_5606, signal_5605, signal_5604, signal_1737}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1723 ( .a ({signal_5351, signal_5350, signal_5349, signal_5348, signal_1673}), .b ({signal_5611, signal_5610, signal_5609, signal_5608, signal_1738}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1724 ( .a ({signal_5363, signal_5362, signal_5361, signal_5360, signal_1676}), .b ({signal_5615, signal_5614, signal_5613, signal_5612, signal_1739}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1726 ( .a ({signal_5371, signal_5370, signal_5369, signal_5368, signal_1678}), .b ({signal_5623, signal_5622, signal_5621, signal_5620, signal_1741}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1727 ( .a ({signal_5375, signal_5374, signal_5373, signal_5372, signal_1679}), .b ({signal_5627, signal_5626, signal_5625, signal_5624, signal_1742}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1728 ( .a ({signal_5379, signal_5378, signal_5377, signal_5376, signal_1680}), .b ({signal_5631, signal_5630, signal_5629, signal_5628, signal_1743}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1729 ( .a ({signal_5383, signal_5382, signal_5381, signal_5380, signal_1681}), .b ({signal_5635, signal_5634, signal_5633, signal_5632, signal_1744}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1730 ( .a ({signal_5387, signal_5386, signal_5385, signal_5384, signal_1682}), .b ({signal_5639, signal_5638, signal_5637, signal_5636, signal_1745}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1731 ( .a ({signal_5403, signal_5402, signal_5401, signal_5400, signal_1686}), .b ({signal_5643, signal_5642, signal_5641, signal_5640, signal_1746}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1732 ( .a ({signal_5415, signal_5414, signal_5413, signal_5412, signal_1689}), .b ({signal_5647, signal_5646, signal_5645, signal_5644, signal_1747}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1733 ( .a ({signal_5431, signal_5430, signal_5429, signal_5428, signal_1693}), .b ({signal_5651, signal_5650, signal_5649, signal_5648, signal_1748}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1734 ( .a ({signal_5443, signal_5442, signal_5441, signal_5440, signal_1696}), .b ({signal_5655, signal_5654, signal_5653, signal_5652, signal_1749}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1735 ( .a ({signal_5447, signal_5446, signal_5445, signal_5444, signal_1697}), .b ({signal_5659, signal_5658, signal_5657, signal_5656, signal_1750}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1736 ( .a ({signal_5455, signal_5454, signal_5453, signal_5452, signal_1699}), .b ({signal_5663, signal_5662, signal_5661, signal_5660, signal_1751}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1739 ( .a ({signal_5467, signal_5466, signal_5465, signal_5464, signal_1702}), .b ({signal_5675, signal_5674, signal_5673, signal_5672, signal_1754}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1745 ( .a ({signal_5491, signal_5490, signal_5489, signal_5488, signal_1708}), .b ({signal_5699, signal_5698, signal_5697, signal_5696, signal_1760}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1749 ( .a ({signal_5511, signal_5510, signal_5509, signal_5508, signal_1713}), .b ({signal_5715, signal_5714, signal_5713, signal_5712, signal_1764}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1751 ( .a ({signal_3067, signal_3066, signal_3065, signal_3064, signal_1102}), .b ({signal_4687, signal_4686, signal_4685, signal_4684, signal_1507}), .clk ( clk ), .r ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280]}), .c ({signal_5723, signal_5722, signal_5721, signal_5720, signal_1766}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1753 ( .a ({signal_17587, signal_17583, signal_17579, signal_17575, signal_17571}), .b ({signal_4691, signal_4690, signal_4689, signal_4688, signal_1508}), .clk ( clk ), .r ({Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .c ({signal_5731, signal_5730, signal_5729, signal_5728, signal_1768}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1754 ( .a ({signal_17467, signal_17465, signal_17463, signal_17461, signal_17459}), .b ({signal_4695, signal_4694, signal_4693, signal_4692, signal_1509}), .clk ( clk ), .r ({Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300]}), .c ({signal_5735, signal_5734, signal_5733, signal_5732, signal_1769}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1755 ( .a ({signal_2991, signal_2990, signal_2989, signal_2988, signal_1083}), .b ({signal_4699, signal_4698, signal_4697, signal_4696, signal_1510}), .clk ( clk ), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310]}), .c ({signal_5739, signal_5738, signal_5737, signal_5736, signal_1770}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1756 ( .a ({signal_17567, signal_17565, signal_17563, signal_17561, signal_17559}), .b ({signal_4687, signal_4686, signal_4685, signal_4684, signal_1507}), .clk ( clk ), .r ({Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({signal_5743, signal_5742, signal_5741, signal_5740, signal_1771}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1757 ( .a ({signal_3187, signal_3186, signal_3185, signal_3184, signal_1132}), .b ({signal_4703, signal_4702, signal_4701, signal_4700, signal_1511}), .clk ( clk ), .r ({Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330]}), .c ({signal_5747, signal_5746, signal_5745, signal_5744, signal_1772}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1758 ( .a ({signal_17697, signal_17695, signal_17693, signal_17691, signal_17689}), .b ({signal_4703, signal_4702, signal_4701, signal_4700, signal_1511}), .clk ( clk ), .r ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340]}), .c ({signal_5751, signal_5750, signal_5749, signal_5748, signal_1773}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1760 ( .a ({signal_17787, signal_17785, signal_17783, signal_17781, signal_17779}), .b ({signal_4715, signal_4714, signal_4713, signal_4712, signal_1514}), .clk ( clk ), .r ({Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .c ({signal_5759, signal_5758, signal_5757, signal_5756, signal_1775}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1761 ( .a ({signal_17797, signal_17795, signal_17793, signal_17791, signal_17789}), .b ({signal_4719, signal_4718, signal_4717, signal_4716, signal_1515}), .clk ( clk ), .r ({Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360]}), .c ({signal_5763, signal_5762, signal_5761, signal_5760, signal_1776}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1762 ( .a ({signal_17267, signal_17265, signal_17263, signal_17261, signal_17259}), .b ({signal_4723, signal_4722, signal_4721, signal_4720, signal_1516}), .clk ( clk ), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370]}), .c ({signal_5767, signal_5766, signal_5765, signal_5764, signal_1777}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1764 ( .a ({signal_17517, signal_17515, signal_17513, signal_17511, signal_17509}), .b ({signal_4735, signal_4734, signal_4733, signal_4732, signal_1519}), .clk ( clk ), .r ({Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({signal_5775, signal_5774, signal_5773, signal_5772, signal_1779}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1765 ( .a ({signal_17757, signal_17755, signal_17753, signal_17751, signal_17749}), .b ({signal_4739, signal_4738, signal_4737, signal_4736, signal_1520}), .clk ( clk ), .r ({Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390]}), .c ({signal_5779, signal_5778, signal_5777, signal_5776, signal_1780}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1766 ( .a ({signal_17297, signal_17295, signal_17293, signal_17291, signal_17289}), .b ({signal_4743, signal_4742, signal_4741, signal_4740, signal_1521}), .clk ( clk ), .r ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400]}), .c ({signal_5783, signal_5782, signal_5781, signal_5780, signal_1781}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1767 ( .a ({signal_17397, signal_17395, signal_17393, signal_17391, signal_17389}), .b ({signal_4747, signal_4746, signal_4745, signal_4744, signal_1522}), .clk ( clk ), .r ({Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .c ({signal_5787, signal_5786, signal_5785, signal_5784, signal_1782}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1769 ( .a ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1078}), .b ({signal_4747, signal_4746, signal_4745, signal_4744, signal_1522}), .clk ( clk ), .r ({Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420]}), .c ({signal_5795, signal_5794, signal_5793, signal_5792, signal_1784}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1770 ( .a ({signal_2999, signal_2998, signal_2997, signal_2996, signal_1085}), .b ({signal_4771, signal_4770, signal_4769, signal_4768, signal_1528}), .clk ( clk ), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430]}), .c ({signal_5799, signal_5798, signal_5797, signal_5796, signal_1785}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1772 ( .a ({signal_17347, signal_17345, signal_17343, signal_17341, signal_17339}), .b ({signal_4743, signal_4742, signal_4741, signal_4740, signal_1521}), .clk ( clk ), .r ({Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({signal_5807, signal_5806, signal_5805, signal_5804, signal_1787}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1773 ( .a ({signal_3271, signal_3270, signal_3269, signal_3268, signal_1153}), .b ({signal_4799, signal_4798, signal_4797, signal_4796, signal_1535}), .clk ( clk ), .r ({Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450]}), .c ({signal_5811, signal_5810, signal_5809, signal_5808, signal_1788}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1776 ( .a ({signal_17637, signal_17635, signal_17633, signal_17631, signal_17629}), .b ({signal_4739, signal_4738, signal_4737, signal_4736, signal_1520}), .clk ( clk ), .r ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460]}), .c ({signal_5823, signal_5822, signal_5821, signal_5820, signal_1791}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1778 ( .a ({signal_17807, signal_17805, signal_17803, signal_17801, signal_17799}), .b ({signal_4847, signal_4846, signal_4845, signal_4844, signal_1547}), .clk ( clk ), .r ({Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .c ({signal_5831, signal_5830, signal_5829, signal_5828, signal_1793}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1779 ( .a ({signal_3003, signal_3002, signal_3001, signal_3000, signal_1086}), .b ({signal_4851, signal_4850, signal_4849, signal_4848, signal_1548}), .clk ( clk ), .r ({Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480]}), .c ({signal_5835, signal_5834, signal_5833, signal_5832, signal_1794}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1782 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_4871, signal_4870, signal_4869, signal_4868, signal_1553}), .clk ( clk ), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490]}), .c ({signal_5847, signal_5846, signal_5845, signal_5844, signal_1797}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1783 ( .a ({signal_17287, signal_17285, signal_17283, signal_17281, signal_17279}), .b ({signal_4875, signal_4874, signal_4873, signal_4872, signal_1554}), .clk ( clk ), .r ({Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({signal_5851, signal_5850, signal_5849, signal_5848, signal_1798}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1784 ( .a ({signal_2987, signal_2986, signal_2985, signal_2984, signal_1082}), .b ({signal_4719, signal_4718, signal_4717, signal_4716, signal_1515}), .clk ( clk ), .r ({Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510]}), .c ({signal_5855, signal_5854, signal_5853, signal_5852, signal_1799}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1785 ( .a ({signal_17617, signal_17615, signal_17613, signal_17611, signal_17609}), .b ({signal_4891, signal_4890, signal_4889, signal_4888, signal_1558}), .clk ( clk ), .r ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520]}), .c ({signal_5859, signal_5858, signal_5857, signal_5856, signal_1800}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1786 ( .a ({signal_17497, signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_4895, signal_4894, signal_4893, signal_4892, signal_1559}), .clk ( clk ), .r ({Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .c ({signal_5863, signal_5862, signal_5861, signal_5860, signal_1801}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1835 ( .a ({signal_5723, signal_5722, signal_5721, signal_5720, signal_1766}), .b ({signal_6059, signal_6058, signal_6057, signal_6056, signal_1850}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1836 ( .a ({signal_5739, signal_5738, signal_5737, signal_5736, signal_1770}), .b ({signal_6063, signal_6062, signal_6061, signal_6060, signal_1851}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1837 ( .a ({signal_5747, signal_5746, signal_5745, signal_5744, signal_1772}), .b ({signal_6067, signal_6066, signal_6065, signal_6064, signal_1852}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1838 ( .a ({signal_5751, signal_5750, signal_5749, signal_5748, signal_1773}), .b ({signal_6071, signal_6070, signal_6069, signal_6068, signal_1853}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1839 ( .a ({signal_5759, signal_5758, signal_5757, signal_5756, signal_1775}), .b ({signal_6075, signal_6074, signal_6073, signal_6072, signal_1854}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1840 ( .a ({signal_5763, signal_5762, signal_5761, signal_5760, signal_1776}), .b ({signal_6079, signal_6078, signal_6077, signal_6076, signal_1855}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1841 ( .a ({signal_5767, signal_5766, signal_5765, signal_5764, signal_1777}), .b ({signal_6083, signal_6082, signal_6081, signal_6080, signal_1856}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1843 ( .a ({signal_5775, signal_5774, signal_5773, signal_5772, signal_1779}), .b ({signal_6091, signal_6090, signal_6089, signal_6088, signal_1858}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1844 ( .a ({signal_5779, signal_5778, signal_5777, signal_5776, signal_1780}), .b ({signal_6095, signal_6094, signal_6093, signal_6092, signal_1859}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1845 ( .a ({signal_5783, signal_5782, signal_5781, signal_5780, signal_1781}), .b ({signal_6099, signal_6098, signal_6097, signal_6096, signal_1860}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1846 ( .a ({signal_5795, signal_5794, signal_5793, signal_5792, signal_1784}), .b ({signal_6103, signal_6102, signal_6101, signal_6100, signal_1861}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1847 ( .a ({signal_5799, signal_5798, signal_5797, signal_5796, signal_1785}), .b ({signal_6107, signal_6106, signal_6105, signal_6104, signal_1862}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1848 ( .a ({signal_5807, signal_5806, signal_5805, signal_5804, signal_1787}), .b ({signal_6111, signal_6110, signal_6109, signal_6108, signal_1863}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1849 ( .a ({signal_5811, signal_5810, signal_5809, signal_5808, signal_1788}), .b ({signal_6115, signal_6114, signal_6113, signal_6112, signal_1864}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1850 ( .a ({signal_5823, signal_5822, signal_5821, signal_5820, signal_1791}), .b ({signal_6119, signal_6118, signal_6117, signal_6116, signal_1865}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1851 ( .a ({signal_5831, signal_5830, signal_5829, signal_5828, signal_1793}), .b ({signal_6123, signal_6122, signal_6121, signal_6120, signal_1866}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1852 ( .a ({signal_5835, signal_5834, signal_5833, signal_5832, signal_1794}), .b ({signal_6127, signal_6126, signal_6125, signal_6124, signal_1867}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1854 ( .a ({signal_5847, signal_5846, signal_5845, signal_5844, signal_1797}), .b ({signal_6135, signal_6134, signal_6133, signal_6132, signal_1869}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1855 ( .a ({signal_5851, signal_5850, signal_5849, signal_5848, signal_1798}), .b ({signal_6139, signal_6138, signal_6137, signal_6136, signal_1870}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1856 ( .a ({signal_5855, signal_5854, signal_5853, signal_5852, signal_1799}), .b ({signal_6143, signal_6142, signal_6141, signal_6140, signal_1871}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1857 ( .a ({signal_5859, signal_5858, signal_5857, signal_5856, signal_1800}), .b ({signal_6147, signal_6146, signal_6145, signal_6144, signal_1872}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1858 ( .a ({signal_5863, signal_5862, signal_5861, signal_5860, signal_1801}), .b ({signal_6151, signal_6150, signal_6149, signal_6148, signal_1873}) ) ;
    buf_clk cell_3116 ( .C ( clk ), .D ( signal_17808 ), .Q ( signal_17809 ) ) ;
    buf_clk cell_3118 ( .C ( clk ), .D ( signal_17810 ), .Q ( signal_17811 ) ) ;
    buf_clk cell_3120 ( .C ( clk ), .D ( signal_17812 ), .Q ( signal_17813 ) ) ;
    buf_clk cell_3122 ( .C ( clk ), .D ( signal_17814 ), .Q ( signal_17815 ) ) ;
    buf_clk cell_3124 ( .C ( clk ), .D ( signal_17816 ), .Q ( signal_17817 ) ) ;
    buf_clk cell_3126 ( .C ( clk ), .D ( signal_17818 ), .Q ( signal_17819 ) ) ;
    buf_clk cell_3128 ( .C ( clk ), .D ( signal_17820 ), .Q ( signal_17821 ) ) ;
    buf_clk cell_3130 ( .C ( clk ), .D ( signal_17822 ), .Q ( signal_17823 ) ) ;
    buf_clk cell_3132 ( .C ( clk ), .D ( signal_17824 ), .Q ( signal_17825 ) ) ;
    buf_clk cell_3134 ( .C ( clk ), .D ( signal_17826 ), .Q ( signal_17827 ) ) ;
    buf_clk cell_3136 ( .C ( clk ), .D ( signal_17828 ), .Q ( signal_17829 ) ) ;
    buf_clk cell_3138 ( .C ( clk ), .D ( signal_17830 ), .Q ( signal_17831 ) ) ;
    buf_clk cell_3140 ( .C ( clk ), .D ( signal_17832 ), .Q ( signal_17833 ) ) ;
    buf_clk cell_3142 ( .C ( clk ), .D ( signal_17834 ), .Q ( signal_17835 ) ) ;
    buf_clk cell_3144 ( .C ( clk ), .D ( signal_17836 ), .Q ( signal_17837 ) ) ;
    buf_clk cell_3146 ( .C ( clk ), .D ( signal_17838 ), .Q ( signal_17839 ) ) ;
    buf_clk cell_3148 ( .C ( clk ), .D ( signal_17840 ), .Q ( signal_17841 ) ) ;
    buf_clk cell_3150 ( .C ( clk ), .D ( signal_17842 ), .Q ( signal_17843 ) ) ;
    buf_clk cell_3152 ( .C ( clk ), .D ( signal_17844 ), .Q ( signal_17845 ) ) ;
    buf_clk cell_3154 ( .C ( clk ), .D ( signal_17846 ), .Q ( signal_17847 ) ) ;
    buf_clk cell_3156 ( .C ( clk ), .D ( signal_17848 ), .Q ( signal_17849 ) ) ;
    buf_clk cell_3158 ( .C ( clk ), .D ( signal_17850 ), .Q ( signal_17851 ) ) ;
    buf_clk cell_3160 ( .C ( clk ), .D ( signal_17852 ), .Q ( signal_17853 ) ) ;
    buf_clk cell_3162 ( .C ( clk ), .D ( signal_17854 ), .Q ( signal_17855 ) ) ;
    buf_clk cell_3164 ( .C ( clk ), .D ( signal_17856 ), .Q ( signal_17857 ) ) ;
    buf_clk cell_3166 ( .C ( clk ), .D ( signal_17858 ), .Q ( signal_17859 ) ) ;
    buf_clk cell_3168 ( .C ( clk ), .D ( signal_17860 ), .Q ( signal_17861 ) ) ;
    buf_clk cell_3170 ( .C ( clk ), .D ( signal_17862 ), .Q ( signal_17863 ) ) ;
    buf_clk cell_3172 ( .C ( clk ), .D ( signal_17864 ), .Q ( signal_17865 ) ) ;
    buf_clk cell_3174 ( .C ( clk ), .D ( signal_17866 ), .Q ( signal_17867 ) ) ;
    buf_clk cell_3176 ( .C ( clk ), .D ( signal_17868 ), .Q ( signal_17869 ) ) ;
    buf_clk cell_3178 ( .C ( clk ), .D ( signal_17870 ), .Q ( signal_17871 ) ) ;
    buf_clk cell_3180 ( .C ( clk ), .D ( signal_17872 ), .Q ( signal_17873 ) ) ;
    buf_clk cell_3182 ( .C ( clk ), .D ( signal_17874 ), .Q ( signal_17875 ) ) ;
    buf_clk cell_3184 ( .C ( clk ), .D ( signal_17876 ), .Q ( signal_17877 ) ) ;
    buf_clk cell_3186 ( .C ( clk ), .D ( signal_17878 ), .Q ( signal_17879 ) ) ;
    buf_clk cell_3188 ( .C ( clk ), .D ( signal_17880 ), .Q ( signal_17881 ) ) ;
    buf_clk cell_3190 ( .C ( clk ), .D ( signal_17882 ), .Q ( signal_17883 ) ) ;
    buf_clk cell_3192 ( .C ( clk ), .D ( signal_17884 ), .Q ( signal_17885 ) ) ;
    buf_clk cell_3194 ( .C ( clk ), .D ( signal_17886 ), .Q ( signal_17887 ) ) ;
    buf_clk cell_3196 ( .C ( clk ), .D ( signal_17888 ), .Q ( signal_17889 ) ) ;
    buf_clk cell_3198 ( .C ( clk ), .D ( signal_17890 ), .Q ( signal_17891 ) ) ;
    buf_clk cell_3200 ( .C ( clk ), .D ( signal_17892 ), .Q ( signal_17893 ) ) ;
    buf_clk cell_3202 ( .C ( clk ), .D ( signal_17894 ), .Q ( signal_17895 ) ) ;
    buf_clk cell_3204 ( .C ( clk ), .D ( signal_17896 ), .Q ( signal_17897 ) ) ;
    buf_clk cell_3206 ( .C ( clk ), .D ( signal_17898 ), .Q ( signal_17899 ) ) ;
    buf_clk cell_3208 ( .C ( clk ), .D ( signal_17900 ), .Q ( signal_17901 ) ) ;
    buf_clk cell_3210 ( .C ( clk ), .D ( signal_17902 ), .Q ( signal_17903 ) ) ;
    buf_clk cell_3212 ( .C ( clk ), .D ( signal_17904 ), .Q ( signal_17905 ) ) ;
    buf_clk cell_3214 ( .C ( clk ), .D ( signal_17906 ), .Q ( signal_17907 ) ) ;
    buf_clk cell_3216 ( .C ( clk ), .D ( signal_17908 ), .Q ( signal_17909 ) ) ;
    buf_clk cell_3218 ( .C ( clk ), .D ( signal_17910 ), .Q ( signal_17911 ) ) ;
    buf_clk cell_3220 ( .C ( clk ), .D ( signal_17912 ), .Q ( signal_17913 ) ) ;
    buf_clk cell_3222 ( .C ( clk ), .D ( signal_17914 ), .Q ( signal_17915 ) ) ;
    buf_clk cell_3224 ( .C ( clk ), .D ( signal_17916 ), .Q ( signal_17917 ) ) ;
    buf_clk cell_3230 ( .C ( clk ), .D ( signal_17922 ), .Q ( signal_17923 ) ) ;
    buf_clk cell_3236 ( .C ( clk ), .D ( signal_17928 ), .Q ( signal_17929 ) ) ;
    buf_clk cell_3242 ( .C ( clk ), .D ( signal_17934 ), .Q ( signal_17935 ) ) ;
    buf_clk cell_3248 ( .C ( clk ), .D ( signal_17940 ), .Q ( signal_17941 ) ) ;
    buf_clk cell_3254 ( .C ( clk ), .D ( signal_17946 ), .Q ( signal_17947 ) ) ;
    buf_clk cell_3256 ( .C ( clk ), .D ( signal_17948 ), .Q ( signal_17949 ) ) ;
    buf_clk cell_3258 ( .C ( clk ), .D ( signal_17950 ), .Q ( signal_17951 ) ) ;
    buf_clk cell_3260 ( .C ( clk ), .D ( signal_17952 ), .Q ( signal_17953 ) ) ;
    buf_clk cell_3262 ( .C ( clk ), .D ( signal_17954 ), .Q ( signal_17955 ) ) ;
    buf_clk cell_3264 ( .C ( clk ), .D ( signal_17956 ), .Q ( signal_17957 ) ) ;
    buf_clk cell_3266 ( .C ( clk ), .D ( signal_17958 ), .Q ( signal_17959 ) ) ;
    buf_clk cell_3268 ( .C ( clk ), .D ( signal_17960 ), .Q ( signal_17961 ) ) ;
    buf_clk cell_3270 ( .C ( clk ), .D ( signal_17962 ), .Q ( signal_17963 ) ) ;
    buf_clk cell_3272 ( .C ( clk ), .D ( signal_17964 ), .Q ( signal_17965 ) ) ;
    buf_clk cell_3274 ( .C ( clk ), .D ( signal_17966 ), .Q ( signal_17967 ) ) ;
    buf_clk cell_3276 ( .C ( clk ), .D ( signal_17968 ), .Q ( signal_17969 ) ) ;
    buf_clk cell_3278 ( .C ( clk ), .D ( signal_17970 ), .Q ( signal_17971 ) ) ;
    buf_clk cell_3280 ( .C ( clk ), .D ( signal_17972 ), .Q ( signal_17973 ) ) ;
    buf_clk cell_3282 ( .C ( clk ), .D ( signal_17974 ), .Q ( signal_17975 ) ) ;
    buf_clk cell_3284 ( .C ( clk ), .D ( signal_17976 ), .Q ( signal_17977 ) ) ;
    buf_clk cell_3286 ( .C ( clk ), .D ( signal_17978 ), .Q ( signal_17979 ) ) ;
    buf_clk cell_3288 ( .C ( clk ), .D ( signal_17980 ), .Q ( signal_17981 ) ) ;
    buf_clk cell_3290 ( .C ( clk ), .D ( signal_17982 ), .Q ( signal_17983 ) ) ;
    buf_clk cell_3292 ( .C ( clk ), .D ( signal_17984 ), .Q ( signal_17985 ) ) ;
    buf_clk cell_3294 ( .C ( clk ), .D ( signal_17986 ), .Q ( signal_17987 ) ) ;
    buf_clk cell_3296 ( .C ( clk ), .D ( signal_17988 ), .Q ( signal_17989 ) ) ;
    buf_clk cell_3298 ( .C ( clk ), .D ( signal_17990 ), .Q ( signal_17991 ) ) ;
    buf_clk cell_3300 ( .C ( clk ), .D ( signal_17992 ), .Q ( signal_17993 ) ) ;
    buf_clk cell_3302 ( .C ( clk ), .D ( signal_17994 ), .Q ( signal_17995 ) ) ;
    buf_clk cell_3304 ( .C ( clk ), .D ( signal_17996 ), .Q ( signal_17997 ) ) ;
    buf_clk cell_3306 ( .C ( clk ), .D ( signal_17998 ), .Q ( signal_17999 ) ) ;
    buf_clk cell_3308 ( .C ( clk ), .D ( signal_18000 ), .Q ( signal_18001 ) ) ;
    buf_clk cell_3310 ( .C ( clk ), .D ( signal_18002 ), .Q ( signal_18003 ) ) ;
    buf_clk cell_3312 ( .C ( clk ), .D ( signal_18004 ), .Q ( signal_18005 ) ) ;
    buf_clk cell_3314 ( .C ( clk ), .D ( signal_18006 ), .Q ( signal_18007 ) ) ;
    buf_clk cell_3316 ( .C ( clk ), .D ( signal_18008 ), .Q ( signal_18009 ) ) ;
    buf_clk cell_3318 ( .C ( clk ), .D ( signal_18010 ), .Q ( signal_18011 ) ) ;
    buf_clk cell_3320 ( .C ( clk ), .D ( signal_18012 ), .Q ( signal_18013 ) ) ;
    buf_clk cell_3322 ( .C ( clk ), .D ( signal_18014 ), .Q ( signal_18015 ) ) ;
    buf_clk cell_3324 ( .C ( clk ), .D ( signal_18016 ), .Q ( signal_18017 ) ) ;
    buf_clk cell_3326 ( .C ( clk ), .D ( signal_18018 ), .Q ( signal_18019 ) ) ;
    buf_clk cell_3328 ( .C ( clk ), .D ( signal_18020 ), .Q ( signal_18021 ) ) ;
    buf_clk cell_3330 ( .C ( clk ), .D ( signal_18022 ), .Q ( signal_18023 ) ) ;
    buf_clk cell_3332 ( .C ( clk ), .D ( signal_18024 ), .Q ( signal_18025 ) ) ;
    buf_clk cell_3334 ( .C ( clk ), .D ( signal_18026 ), .Q ( signal_18027 ) ) ;
    buf_clk cell_3336 ( .C ( clk ), .D ( signal_18028 ), .Q ( signal_18029 ) ) ;
    buf_clk cell_3338 ( .C ( clk ), .D ( signal_18030 ), .Q ( signal_18031 ) ) ;
    buf_clk cell_3340 ( .C ( clk ), .D ( signal_18032 ), .Q ( signal_18033 ) ) ;
    buf_clk cell_3342 ( .C ( clk ), .D ( signal_18034 ), .Q ( signal_18035 ) ) ;
    buf_clk cell_3344 ( .C ( clk ), .D ( signal_18036 ), .Q ( signal_18037 ) ) ;
    buf_clk cell_3346 ( .C ( clk ), .D ( signal_18038 ), .Q ( signal_18039 ) ) ;
    buf_clk cell_3348 ( .C ( clk ), .D ( signal_18040 ), .Q ( signal_18041 ) ) ;
    buf_clk cell_3350 ( .C ( clk ), .D ( signal_18042 ), .Q ( signal_18043 ) ) ;
    buf_clk cell_3352 ( .C ( clk ), .D ( signal_18044 ), .Q ( signal_18045 ) ) ;
    buf_clk cell_3354 ( .C ( clk ), .D ( signal_18046 ), .Q ( signal_18047 ) ) ;
    buf_clk cell_3356 ( .C ( clk ), .D ( signal_18048 ), .Q ( signal_18049 ) ) ;
    buf_clk cell_3358 ( .C ( clk ), .D ( signal_18050 ), .Q ( signal_18051 ) ) ;
    buf_clk cell_3360 ( .C ( clk ), .D ( signal_18052 ), .Q ( signal_18053 ) ) ;
    buf_clk cell_3362 ( .C ( clk ), .D ( signal_18054 ), .Q ( signal_18055 ) ) ;
    buf_clk cell_3364 ( .C ( clk ), .D ( signal_18056 ), .Q ( signal_18057 ) ) ;
    buf_clk cell_3366 ( .C ( clk ), .D ( signal_18058 ), .Q ( signal_18059 ) ) ;
    buf_clk cell_3368 ( .C ( clk ), .D ( signal_18060 ), .Q ( signal_18061 ) ) ;
    buf_clk cell_3370 ( .C ( clk ), .D ( signal_18062 ), .Q ( signal_18063 ) ) ;
    buf_clk cell_3372 ( .C ( clk ), .D ( signal_18064 ), .Q ( signal_18065 ) ) ;
    buf_clk cell_3374 ( .C ( clk ), .D ( signal_18066 ), .Q ( signal_18067 ) ) ;
    buf_clk cell_3376 ( .C ( clk ), .D ( signal_18068 ), .Q ( signal_18069 ) ) ;
    buf_clk cell_3378 ( .C ( clk ), .D ( signal_18070 ), .Q ( signal_18071 ) ) ;
    buf_clk cell_3380 ( .C ( clk ), .D ( signal_18072 ), .Q ( signal_18073 ) ) ;
    buf_clk cell_3382 ( .C ( clk ), .D ( signal_18074 ), .Q ( signal_18075 ) ) ;
    buf_clk cell_3384 ( .C ( clk ), .D ( signal_18076 ), .Q ( signal_18077 ) ) ;
    buf_clk cell_3386 ( .C ( clk ), .D ( signal_18078 ), .Q ( signal_18079 ) ) ;
    buf_clk cell_3388 ( .C ( clk ), .D ( signal_18080 ), .Q ( signal_18081 ) ) ;
    buf_clk cell_3390 ( .C ( clk ), .D ( signal_18082 ), .Q ( signal_18083 ) ) ;
    buf_clk cell_3392 ( .C ( clk ), .D ( signal_18084 ), .Q ( signal_18085 ) ) ;
    buf_clk cell_3394 ( .C ( clk ), .D ( signal_18086 ), .Q ( signal_18087 ) ) ;
    buf_clk cell_3396 ( .C ( clk ), .D ( signal_18088 ), .Q ( signal_18089 ) ) ;
    buf_clk cell_3398 ( .C ( clk ), .D ( signal_18090 ), .Q ( signal_18091 ) ) ;
    buf_clk cell_3400 ( .C ( clk ), .D ( signal_18092 ), .Q ( signal_18093 ) ) ;
    buf_clk cell_3402 ( .C ( clk ), .D ( signal_18094 ), .Q ( signal_18095 ) ) ;
    buf_clk cell_3404 ( .C ( clk ), .D ( signal_18096 ), .Q ( signal_18097 ) ) ;
    buf_clk cell_3406 ( .C ( clk ), .D ( signal_18098 ), .Q ( signal_18099 ) ) ;
    buf_clk cell_3408 ( .C ( clk ), .D ( signal_18100 ), .Q ( signal_18101 ) ) ;
    buf_clk cell_3410 ( .C ( clk ), .D ( signal_18102 ), .Q ( signal_18103 ) ) ;
    buf_clk cell_3412 ( .C ( clk ), .D ( signal_18104 ), .Q ( signal_18105 ) ) ;
    buf_clk cell_3414 ( .C ( clk ), .D ( signal_18106 ), .Q ( signal_18107 ) ) ;
    buf_clk cell_3416 ( .C ( clk ), .D ( signal_18108 ), .Q ( signal_18109 ) ) ;
    buf_clk cell_3418 ( .C ( clk ), .D ( signal_18110 ), .Q ( signal_18111 ) ) ;
    buf_clk cell_3420 ( .C ( clk ), .D ( signal_18112 ), .Q ( signal_18113 ) ) ;
    buf_clk cell_3422 ( .C ( clk ), .D ( signal_18114 ), .Q ( signal_18115 ) ) ;
    buf_clk cell_3424 ( .C ( clk ), .D ( signal_18116 ), .Q ( signal_18117 ) ) ;
    buf_clk cell_3426 ( .C ( clk ), .D ( signal_18118 ), .Q ( signal_18119 ) ) ;
    buf_clk cell_3428 ( .C ( clk ), .D ( signal_18120 ), .Q ( signal_18121 ) ) ;
    buf_clk cell_3430 ( .C ( clk ), .D ( signal_18122 ), .Q ( signal_18123 ) ) ;
    buf_clk cell_3432 ( .C ( clk ), .D ( signal_18124 ), .Q ( signal_18125 ) ) ;
    buf_clk cell_3434 ( .C ( clk ), .D ( signal_18126 ), .Q ( signal_18127 ) ) ;
    buf_clk cell_3436 ( .C ( clk ), .D ( signal_18128 ), .Q ( signal_18129 ) ) ;
    buf_clk cell_3438 ( .C ( clk ), .D ( signal_18130 ), .Q ( signal_18131 ) ) ;
    buf_clk cell_3440 ( .C ( clk ), .D ( signal_18132 ), .Q ( signal_18133 ) ) ;
    buf_clk cell_3442 ( .C ( clk ), .D ( signal_18134 ), .Q ( signal_18135 ) ) ;
    buf_clk cell_3444 ( .C ( clk ), .D ( signal_18136 ), .Q ( signal_18137 ) ) ;
    buf_clk cell_3446 ( .C ( clk ), .D ( signal_18138 ), .Q ( signal_18139 ) ) ;
    buf_clk cell_3448 ( .C ( clk ), .D ( signal_18140 ), .Q ( signal_18141 ) ) ;
    buf_clk cell_3450 ( .C ( clk ), .D ( signal_18142 ), .Q ( signal_18143 ) ) ;
    buf_clk cell_3452 ( .C ( clk ), .D ( signal_18144 ), .Q ( signal_18145 ) ) ;
    buf_clk cell_3454 ( .C ( clk ), .D ( signal_18146 ), .Q ( signal_18147 ) ) ;
    buf_clk cell_3458 ( .C ( clk ), .D ( signal_18150 ), .Q ( signal_18151 ) ) ;
    buf_clk cell_3462 ( .C ( clk ), .D ( signal_18154 ), .Q ( signal_18155 ) ) ;
    buf_clk cell_3466 ( .C ( clk ), .D ( signal_18158 ), .Q ( signal_18159 ) ) ;
    buf_clk cell_3470 ( .C ( clk ), .D ( signal_18162 ), .Q ( signal_18163 ) ) ;
    buf_clk cell_3474 ( .C ( clk ), .D ( signal_18166 ), .Q ( signal_18167 ) ) ;
    buf_clk cell_3476 ( .C ( clk ), .D ( signal_18168 ), .Q ( signal_18169 ) ) ;
    buf_clk cell_3478 ( .C ( clk ), .D ( signal_18170 ), .Q ( signal_18171 ) ) ;
    buf_clk cell_3480 ( .C ( clk ), .D ( signal_18172 ), .Q ( signal_18173 ) ) ;
    buf_clk cell_3482 ( .C ( clk ), .D ( signal_18174 ), .Q ( signal_18175 ) ) ;
    buf_clk cell_3484 ( .C ( clk ), .D ( signal_18176 ), .Q ( signal_18177 ) ) ;
    buf_clk cell_3486 ( .C ( clk ), .D ( signal_18178 ), .Q ( signal_18179 ) ) ;
    buf_clk cell_3488 ( .C ( clk ), .D ( signal_18180 ), .Q ( signal_18181 ) ) ;
    buf_clk cell_3490 ( .C ( clk ), .D ( signal_18182 ), .Q ( signal_18183 ) ) ;
    buf_clk cell_3492 ( .C ( clk ), .D ( signal_18184 ), .Q ( signal_18185 ) ) ;
    buf_clk cell_3494 ( .C ( clk ), .D ( signal_18186 ), .Q ( signal_18187 ) ) ;
    buf_clk cell_3498 ( .C ( clk ), .D ( signal_18190 ), .Q ( signal_18191 ) ) ;
    buf_clk cell_3502 ( .C ( clk ), .D ( signal_18194 ), .Q ( signal_18195 ) ) ;
    buf_clk cell_3506 ( .C ( clk ), .D ( signal_18198 ), .Q ( signal_18199 ) ) ;
    buf_clk cell_3510 ( .C ( clk ), .D ( signal_18202 ), .Q ( signal_18203 ) ) ;
    buf_clk cell_3514 ( .C ( clk ), .D ( signal_18206 ), .Q ( signal_18207 ) ) ;
    buf_clk cell_3516 ( .C ( clk ), .D ( signal_18208 ), .Q ( signal_18209 ) ) ;
    buf_clk cell_3518 ( .C ( clk ), .D ( signal_18210 ), .Q ( signal_18211 ) ) ;
    buf_clk cell_3520 ( .C ( clk ), .D ( signal_18212 ), .Q ( signal_18213 ) ) ;
    buf_clk cell_3522 ( .C ( clk ), .D ( signal_18214 ), .Q ( signal_18215 ) ) ;
    buf_clk cell_3524 ( .C ( clk ), .D ( signal_18216 ), .Q ( signal_18217 ) ) ;
    buf_clk cell_3526 ( .C ( clk ), .D ( signal_18218 ), .Q ( signal_18219 ) ) ;
    buf_clk cell_3528 ( .C ( clk ), .D ( signal_18220 ), .Q ( signal_18221 ) ) ;
    buf_clk cell_3530 ( .C ( clk ), .D ( signal_18222 ), .Q ( signal_18223 ) ) ;
    buf_clk cell_3532 ( .C ( clk ), .D ( signal_18224 ), .Q ( signal_18225 ) ) ;
    buf_clk cell_3534 ( .C ( clk ), .D ( signal_18226 ), .Q ( signal_18227 ) ) ;
    buf_clk cell_3536 ( .C ( clk ), .D ( signal_18228 ), .Q ( signal_18229 ) ) ;
    buf_clk cell_3538 ( .C ( clk ), .D ( signal_18230 ), .Q ( signal_18231 ) ) ;
    buf_clk cell_3540 ( .C ( clk ), .D ( signal_18232 ), .Q ( signal_18233 ) ) ;
    buf_clk cell_3542 ( .C ( clk ), .D ( signal_18234 ), .Q ( signal_18235 ) ) ;
    buf_clk cell_3544 ( .C ( clk ), .D ( signal_18236 ), .Q ( signal_18237 ) ) ;
    buf_clk cell_3546 ( .C ( clk ), .D ( signal_18238 ), .Q ( signal_18239 ) ) ;
    buf_clk cell_3548 ( .C ( clk ), .D ( signal_18240 ), .Q ( signal_18241 ) ) ;
    buf_clk cell_3550 ( .C ( clk ), .D ( signal_18242 ), .Q ( signal_18243 ) ) ;
    buf_clk cell_3552 ( .C ( clk ), .D ( signal_18244 ), .Q ( signal_18245 ) ) ;
    buf_clk cell_3554 ( .C ( clk ), .D ( signal_18246 ), .Q ( signal_18247 ) ) ;
    buf_clk cell_3556 ( .C ( clk ), .D ( signal_18248 ), .Q ( signal_18249 ) ) ;
    buf_clk cell_3558 ( .C ( clk ), .D ( signal_18250 ), .Q ( signal_18251 ) ) ;
    buf_clk cell_3560 ( .C ( clk ), .D ( signal_18252 ), .Q ( signal_18253 ) ) ;
    buf_clk cell_3562 ( .C ( clk ), .D ( signal_18254 ), .Q ( signal_18255 ) ) ;
    buf_clk cell_3564 ( .C ( clk ), .D ( signal_18256 ), .Q ( signal_18257 ) ) ;
    buf_clk cell_3566 ( .C ( clk ), .D ( signal_18258 ), .Q ( signal_18259 ) ) ;
    buf_clk cell_3568 ( .C ( clk ), .D ( signal_18260 ), .Q ( signal_18261 ) ) ;
    buf_clk cell_3570 ( .C ( clk ), .D ( signal_18262 ), .Q ( signal_18263 ) ) ;
    buf_clk cell_3572 ( .C ( clk ), .D ( signal_18264 ), .Q ( signal_18265 ) ) ;
    buf_clk cell_3574 ( .C ( clk ), .D ( signal_18266 ), .Q ( signal_18267 ) ) ;
    buf_clk cell_3576 ( .C ( clk ), .D ( signal_18268 ), .Q ( signal_18269 ) ) ;
    buf_clk cell_3578 ( .C ( clk ), .D ( signal_18270 ), .Q ( signal_18271 ) ) ;
    buf_clk cell_3580 ( .C ( clk ), .D ( signal_18272 ), .Q ( signal_18273 ) ) ;
    buf_clk cell_3582 ( .C ( clk ), .D ( signal_18274 ), .Q ( signal_18275 ) ) ;
    buf_clk cell_3584 ( .C ( clk ), .D ( signal_18276 ), .Q ( signal_18277 ) ) ;
    buf_clk cell_3586 ( .C ( clk ), .D ( signal_18278 ), .Q ( signal_18279 ) ) ;
    buf_clk cell_3588 ( .C ( clk ), .D ( signal_18280 ), .Q ( signal_18281 ) ) ;
    buf_clk cell_3590 ( .C ( clk ), .D ( signal_18282 ), .Q ( signal_18283 ) ) ;
    buf_clk cell_3592 ( .C ( clk ), .D ( signal_18284 ), .Q ( signal_18285 ) ) ;
    buf_clk cell_3594 ( .C ( clk ), .D ( signal_18286 ), .Q ( signal_18287 ) ) ;
    buf_clk cell_3596 ( .C ( clk ), .D ( signal_18288 ), .Q ( signal_18289 ) ) ;
    buf_clk cell_3598 ( .C ( clk ), .D ( signal_18290 ), .Q ( signal_18291 ) ) ;
    buf_clk cell_3600 ( .C ( clk ), .D ( signal_18292 ), .Q ( signal_18293 ) ) ;
    buf_clk cell_3602 ( .C ( clk ), .D ( signal_18294 ), .Q ( signal_18295 ) ) ;
    buf_clk cell_3604 ( .C ( clk ), .D ( signal_18296 ), .Q ( signal_18297 ) ) ;
    buf_clk cell_3606 ( .C ( clk ), .D ( signal_18298 ), .Q ( signal_18299 ) ) ;
    buf_clk cell_3608 ( .C ( clk ), .D ( signal_18300 ), .Q ( signal_18301 ) ) ;
    buf_clk cell_3610 ( .C ( clk ), .D ( signal_18302 ), .Q ( signal_18303 ) ) ;
    buf_clk cell_3612 ( .C ( clk ), .D ( signal_18304 ), .Q ( signal_18305 ) ) ;
    buf_clk cell_3614 ( .C ( clk ), .D ( signal_18306 ), .Q ( signal_18307 ) ) ;
    buf_clk cell_3616 ( .C ( clk ), .D ( signal_18308 ), .Q ( signal_18309 ) ) ;
    buf_clk cell_3618 ( .C ( clk ), .D ( signal_18310 ), .Q ( signal_18311 ) ) ;
    buf_clk cell_3620 ( .C ( clk ), .D ( signal_18312 ), .Q ( signal_18313 ) ) ;
    buf_clk cell_3622 ( .C ( clk ), .D ( signal_18314 ), .Q ( signal_18315 ) ) ;
    buf_clk cell_3624 ( .C ( clk ), .D ( signal_18316 ), .Q ( signal_18317 ) ) ;
    buf_clk cell_3628 ( .C ( clk ), .D ( signal_18320 ), .Q ( signal_18321 ) ) ;
    buf_clk cell_3632 ( .C ( clk ), .D ( signal_18324 ), .Q ( signal_18325 ) ) ;
    buf_clk cell_3636 ( .C ( clk ), .D ( signal_18328 ), .Q ( signal_18329 ) ) ;
    buf_clk cell_3640 ( .C ( clk ), .D ( signal_18332 ), .Q ( signal_18333 ) ) ;
    buf_clk cell_3644 ( .C ( clk ), .D ( signal_18336 ), .Q ( signal_18337 ) ) ;
    buf_clk cell_3646 ( .C ( clk ), .D ( signal_18338 ), .Q ( signal_18339 ) ) ;
    buf_clk cell_3648 ( .C ( clk ), .D ( signal_18340 ), .Q ( signal_18341 ) ) ;
    buf_clk cell_3650 ( .C ( clk ), .D ( signal_18342 ), .Q ( signal_18343 ) ) ;
    buf_clk cell_3652 ( .C ( clk ), .D ( signal_18344 ), .Q ( signal_18345 ) ) ;
    buf_clk cell_3654 ( .C ( clk ), .D ( signal_18346 ), .Q ( signal_18347 ) ) ;
    buf_clk cell_3658 ( .C ( clk ), .D ( signal_18350 ), .Q ( signal_18351 ) ) ;
    buf_clk cell_3662 ( .C ( clk ), .D ( signal_18354 ), .Q ( signal_18355 ) ) ;
    buf_clk cell_3666 ( .C ( clk ), .D ( signal_18358 ), .Q ( signal_18359 ) ) ;
    buf_clk cell_3670 ( .C ( clk ), .D ( signal_18362 ), .Q ( signal_18363 ) ) ;
    buf_clk cell_3674 ( .C ( clk ), .D ( signal_18366 ), .Q ( signal_18367 ) ) ;
    buf_clk cell_3676 ( .C ( clk ), .D ( signal_18368 ), .Q ( signal_18369 ) ) ;
    buf_clk cell_3678 ( .C ( clk ), .D ( signal_18370 ), .Q ( signal_18371 ) ) ;
    buf_clk cell_3680 ( .C ( clk ), .D ( signal_18372 ), .Q ( signal_18373 ) ) ;
    buf_clk cell_3682 ( .C ( clk ), .D ( signal_18374 ), .Q ( signal_18375 ) ) ;
    buf_clk cell_3684 ( .C ( clk ), .D ( signal_18376 ), .Q ( signal_18377 ) ) ;
    buf_clk cell_3686 ( .C ( clk ), .D ( signal_18378 ), .Q ( signal_18379 ) ) ;
    buf_clk cell_3688 ( .C ( clk ), .D ( signal_18380 ), .Q ( signal_18381 ) ) ;
    buf_clk cell_3690 ( .C ( clk ), .D ( signal_18382 ), .Q ( signal_18383 ) ) ;
    buf_clk cell_3692 ( .C ( clk ), .D ( signal_18384 ), .Q ( signal_18385 ) ) ;
    buf_clk cell_3694 ( .C ( clk ), .D ( signal_18386 ), .Q ( signal_18387 ) ) ;
    buf_clk cell_3696 ( .C ( clk ), .D ( signal_18388 ), .Q ( signal_18389 ) ) ;
    buf_clk cell_3698 ( .C ( clk ), .D ( signal_18390 ), .Q ( signal_18391 ) ) ;
    buf_clk cell_3700 ( .C ( clk ), .D ( signal_18392 ), .Q ( signal_18393 ) ) ;
    buf_clk cell_3702 ( .C ( clk ), .D ( signal_18394 ), .Q ( signal_18395 ) ) ;
    buf_clk cell_3704 ( .C ( clk ), .D ( signal_18396 ), .Q ( signal_18397 ) ) ;
    buf_clk cell_3710 ( .C ( clk ), .D ( signal_18402 ), .Q ( signal_18403 ) ) ;
    buf_clk cell_3716 ( .C ( clk ), .D ( signal_18408 ), .Q ( signal_18409 ) ) ;
    buf_clk cell_3722 ( .C ( clk ), .D ( signal_18414 ), .Q ( signal_18415 ) ) ;
    buf_clk cell_3728 ( .C ( clk ), .D ( signal_18420 ), .Q ( signal_18421 ) ) ;
    buf_clk cell_3734 ( .C ( clk ), .D ( signal_18426 ), .Q ( signal_18427 ) ) ;
    buf_clk cell_3736 ( .C ( clk ), .D ( signal_18428 ), .Q ( signal_18429 ) ) ;
    buf_clk cell_3738 ( .C ( clk ), .D ( signal_18430 ), .Q ( signal_18431 ) ) ;
    buf_clk cell_3740 ( .C ( clk ), .D ( signal_18432 ), .Q ( signal_18433 ) ) ;
    buf_clk cell_3742 ( .C ( clk ), .D ( signal_18434 ), .Q ( signal_18435 ) ) ;
    buf_clk cell_3744 ( .C ( clk ), .D ( signal_18436 ), .Q ( signal_18437 ) ) ;
    buf_clk cell_3746 ( .C ( clk ), .D ( signal_18438 ), .Q ( signal_18439 ) ) ;
    buf_clk cell_3748 ( .C ( clk ), .D ( signal_18440 ), .Q ( signal_18441 ) ) ;
    buf_clk cell_3750 ( .C ( clk ), .D ( signal_18442 ), .Q ( signal_18443 ) ) ;
    buf_clk cell_3752 ( .C ( clk ), .D ( signal_18444 ), .Q ( signal_18445 ) ) ;
    buf_clk cell_3754 ( .C ( clk ), .D ( signal_18446 ), .Q ( signal_18447 ) ) ;
    buf_clk cell_3756 ( .C ( clk ), .D ( signal_18448 ), .Q ( signal_18449 ) ) ;
    buf_clk cell_3758 ( .C ( clk ), .D ( signal_18450 ), .Q ( signal_18451 ) ) ;
    buf_clk cell_3760 ( .C ( clk ), .D ( signal_18452 ), .Q ( signal_18453 ) ) ;
    buf_clk cell_3762 ( .C ( clk ), .D ( signal_18454 ), .Q ( signal_18455 ) ) ;
    buf_clk cell_3764 ( .C ( clk ), .D ( signal_18456 ), .Q ( signal_18457 ) ) ;
    buf_clk cell_3766 ( .C ( clk ), .D ( signal_18458 ), .Q ( signal_18459 ) ) ;
    buf_clk cell_3768 ( .C ( clk ), .D ( signal_18460 ), .Q ( signal_18461 ) ) ;
    buf_clk cell_3770 ( .C ( clk ), .D ( signal_18462 ), .Q ( signal_18463 ) ) ;
    buf_clk cell_3772 ( .C ( clk ), .D ( signal_18464 ), .Q ( signal_18465 ) ) ;
    buf_clk cell_3774 ( .C ( clk ), .D ( signal_18466 ), .Q ( signal_18467 ) ) ;
    buf_clk cell_3778 ( .C ( clk ), .D ( signal_18470 ), .Q ( signal_18471 ) ) ;
    buf_clk cell_3782 ( .C ( clk ), .D ( signal_18474 ), .Q ( signal_18475 ) ) ;
    buf_clk cell_3786 ( .C ( clk ), .D ( signal_18478 ), .Q ( signal_18479 ) ) ;
    buf_clk cell_3790 ( .C ( clk ), .D ( signal_18482 ), .Q ( signal_18483 ) ) ;
    buf_clk cell_3794 ( .C ( clk ), .D ( signal_18486 ), .Q ( signal_18487 ) ) ;
    buf_clk cell_3796 ( .C ( clk ), .D ( signal_18488 ), .Q ( signal_18489 ) ) ;
    buf_clk cell_3798 ( .C ( clk ), .D ( signal_18490 ), .Q ( signal_18491 ) ) ;
    buf_clk cell_3800 ( .C ( clk ), .D ( signal_18492 ), .Q ( signal_18493 ) ) ;
    buf_clk cell_3802 ( .C ( clk ), .D ( signal_18494 ), .Q ( signal_18495 ) ) ;
    buf_clk cell_3804 ( .C ( clk ), .D ( signal_18496 ), .Q ( signal_18497 ) ) ;
    buf_clk cell_3806 ( .C ( clk ), .D ( signal_18498 ), .Q ( signal_18499 ) ) ;
    buf_clk cell_3808 ( .C ( clk ), .D ( signal_18500 ), .Q ( signal_18501 ) ) ;
    buf_clk cell_3810 ( .C ( clk ), .D ( signal_18502 ), .Q ( signal_18503 ) ) ;
    buf_clk cell_3812 ( .C ( clk ), .D ( signal_18504 ), .Q ( signal_18505 ) ) ;
    buf_clk cell_3814 ( .C ( clk ), .D ( signal_18506 ), .Q ( signal_18507 ) ) ;
    buf_clk cell_3816 ( .C ( clk ), .D ( signal_18508 ), .Q ( signal_18509 ) ) ;
    buf_clk cell_3818 ( .C ( clk ), .D ( signal_18510 ), .Q ( signal_18511 ) ) ;
    buf_clk cell_3820 ( .C ( clk ), .D ( signal_18512 ), .Q ( signal_18513 ) ) ;
    buf_clk cell_3822 ( .C ( clk ), .D ( signal_18514 ), .Q ( signal_18515 ) ) ;
    buf_clk cell_3824 ( .C ( clk ), .D ( signal_18516 ), .Q ( signal_18517 ) ) ;
    buf_clk cell_3826 ( .C ( clk ), .D ( signal_18518 ), .Q ( signal_18519 ) ) ;
    buf_clk cell_3828 ( .C ( clk ), .D ( signal_18520 ), .Q ( signal_18521 ) ) ;
    buf_clk cell_3830 ( .C ( clk ), .D ( signal_18522 ), .Q ( signal_18523 ) ) ;
    buf_clk cell_3832 ( .C ( clk ), .D ( signal_18524 ), .Q ( signal_18525 ) ) ;
    buf_clk cell_3834 ( .C ( clk ), .D ( signal_18526 ), .Q ( signal_18527 ) ) ;
    buf_clk cell_3836 ( .C ( clk ), .D ( signal_18528 ), .Q ( signal_18529 ) ) ;
    buf_clk cell_3838 ( .C ( clk ), .D ( signal_18530 ), .Q ( signal_18531 ) ) ;
    buf_clk cell_3840 ( .C ( clk ), .D ( signal_18532 ), .Q ( signal_18533 ) ) ;
    buf_clk cell_3842 ( .C ( clk ), .D ( signal_18534 ), .Q ( signal_18535 ) ) ;
    buf_clk cell_3844 ( .C ( clk ), .D ( signal_18536 ), .Q ( signal_18537 ) ) ;
    buf_clk cell_3846 ( .C ( clk ), .D ( signal_18538 ), .Q ( signal_18539 ) ) ;
    buf_clk cell_3848 ( .C ( clk ), .D ( signal_18540 ), .Q ( signal_18541 ) ) ;
    buf_clk cell_3850 ( .C ( clk ), .D ( signal_18542 ), .Q ( signal_18543 ) ) ;
    buf_clk cell_3852 ( .C ( clk ), .D ( signal_18544 ), .Q ( signal_18545 ) ) ;
    buf_clk cell_3854 ( .C ( clk ), .D ( signal_18546 ), .Q ( signal_18547 ) ) ;
    buf_clk cell_3856 ( .C ( clk ), .D ( signal_18548 ), .Q ( signal_18549 ) ) ;
    buf_clk cell_3858 ( .C ( clk ), .D ( signal_18550 ), .Q ( signal_18551 ) ) ;
    buf_clk cell_3860 ( .C ( clk ), .D ( signal_18552 ), .Q ( signal_18553 ) ) ;
    buf_clk cell_3862 ( .C ( clk ), .D ( signal_18554 ), .Q ( signal_18555 ) ) ;
    buf_clk cell_3864 ( .C ( clk ), .D ( signal_18556 ), .Q ( signal_18557 ) ) ;
    buf_clk cell_3866 ( .C ( clk ), .D ( signal_18558 ), .Q ( signal_18559 ) ) ;
    buf_clk cell_3868 ( .C ( clk ), .D ( signal_18560 ), .Q ( signal_18561 ) ) ;
    buf_clk cell_3870 ( .C ( clk ), .D ( signal_18562 ), .Q ( signal_18563 ) ) ;
    buf_clk cell_3872 ( .C ( clk ), .D ( signal_18564 ), .Q ( signal_18565 ) ) ;
    buf_clk cell_3874 ( .C ( clk ), .D ( signal_18566 ), .Q ( signal_18567 ) ) ;
    buf_clk cell_3876 ( .C ( clk ), .D ( signal_18568 ), .Q ( signal_18569 ) ) ;
    buf_clk cell_3878 ( .C ( clk ), .D ( signal_18570 ), .Q ( signal_18571 ) ) ;
    buf_clk cell_3880 ( .C ( clk ), .D ( signal_18572 ), .Q ( signal_18573 ) ) ;
    buf_clk cell_3882 ( .C ( clk ), .D ( signal_18574 ), .Q ( signal_18575 ) ) ;
    buf_clk cell_3884 ( .C ( clk ), .D ( signal_18576 ), .Q ( signal_18577 ) ) ;
    buf_clk cell_3888 ( .C ( clk ), .D ( signal_18580 ), .Q ( signal_18581 ) ) ;
    buf_clk cell_3892 ( .C ( clk ), .D ( signal_18584 ), .Q ( signal_18585 ) ) ;
    buf_clk cell_3896 ( .C ( clk ), .D ( signal_18588 ), .Q ( signal_18589 ) ) ;
    buf_clk cell_3900 ( .C ( clk ), .D ( signal_18592 ), .Q ( signal_18593 ) ) ;
    buf_clk cell_3904 ( .C ( clk ), .D ( signal_18596 ), .Q ( signal_18597 ) ) ;
    buf_clk cell_3906 ( .C ( clk ), .D ( signal_18598 ), .Q ( signal_18599 ) ) ;
    buf_clk cell_3908 ( .C ( clk ), .D ( signal_18600 ), .Q ( signal_18601 ) ) ;
    buf_clk cell_3910 ( .C ( clk ), .D ( signal_18602 ), .Q ( signal_18603 ) ) ;
    buf_clk cell_3912 ( .C ( clk ), .D ( signal_18604 ), .Q ( signal_18605 ) ) ;
    buf_clk cell_3914 ( .C ( clk ), .D ( signal_18606 ), .Q ( signal_18607 ) ) ;
    buf_clk cell_3916 ( .C ( clk ), .D ( signal_18608 ), .Q ( signal_18609 ) ) ;
    buf_clk cell_3918 ( .C ( clk ), .D ( signal_18610 ), .Q ( signal_18611 ) ) ;
    buf_clk cell_3920 ( .C ( clk ), .D ( signal_18612 ), .Q ( signal_18613 ) ) ;
    buf_clk cell_3922 ( .C ( clk ), .D ( signal_18614 ), .Q ( signal_18615 ) ) ;
    buf_clk cell_3924 ( .C ( clk ), .D ( signal_18616 ), .Q ( signal_18617 ) ) ;
    buf_clk cell_3926 ( .C ( clk ), .D ( signal_18618 ), .Q ( signal_18619 ) ) ;
    buf_clk cell_3928 ( .C ( clk ), .D ( signal_18620 ), .Q ( signal_18621 ) ) ;
    buf_clk cell_3930 ( .C ( clk ), .D ( signal_18622 ), .Q ( signal_18623 ) ) ;
    buf_clk cell_3932 ( .C ( clk ), .D ( signal_18624 ), .Q ( signal_18625 ) ) ;
    buf_clk cell_3934 ( .C ( clk ), .D ( signal_18626 ), .Q ( signal_18627 ) ) ;
    buf_clk cell_3936 ( .C ( clk ), .D ( signal_18628 ), .Q ( signal_18629 ) ) ;
    buf_clk cell_3938 ( .C ( clk ), .D ( signal_18630 ), .Q ( signal_18631 ) ) ;
    buf_clk cell_3940 ( .C ( clk ), .D ( signal_18632 ), .Q ( signal_18633 ) ) ;
    buf_clk cell_3942 ( .C ( clk ), .D ( signal_18634 ), .Q ( signal_18635 ) ) ;
    buf_clk cell_3944 ( .C ( clk ), .D ( signal_18636 ), .Q ( signal_18637 ) ) ;
    buf_clk cell_3946 ( .C ( clk ), .D ( signal_18638 ), .Q ( signal_18639 ) ) ;
    buf_clk cell_3948 ( .C ( clk ), .D ( signal_18640 ), .Q ( signal_18641 ) ) ;
    buf_clk cell_3950 ( .C ( clk ), .D ( signal_18642 ), .Q ( signal_18643 ) ) ;
    buf_clk cell_3952 ( .C ( clk ), .D ( signal_18644 ), .Q ( signal_18645 ) ) ;
    buf_clk cell_3954 ( .C ( clk ), .D ( signal_18646 ), .Q ( signal_18647 ) ) ;
    buf_clk cell_3956 ( .C ( clk ), .D ( signal_18648 ), .Q ( signal_18649 ) ) ;
    buf_clk cell_3958 ( .C ( clk ), .D ( signal_18650 ), .Q ( signal_18651 ) ) ;
    buf_clk cell_3960 ( .C ( clk ), .D ( signal_18652 ), .Q ( signal_18653 ) ) ;
    buf_clk cell_3962 ( .C ( clk ), .D ( signal_18654 ), .Q ( signal_18655 ) ) ;
    buf_clk cell_3964 ( .C ( clk ), .D ( signal_18656 ), .Q ( signal_18657 ) ) ;
    buf_clk cell_3986 ( .C ( clk ), .D ( signal_18678 ), .Q ( signal_18679 ) ) ;
    buf_clk cell_3990 ( .C ( clk ), .D ( signal_18682 ), .Q ( signal_18683 ) ) ;
    buf_clk cell_3994 ( .C ( clk ), .D ( signal_18686 ), .Q ( signal_18687 ) ) ;
    buf_clk cell_3998 ( .C ( clk ), .D ( signal_18690 ), .Q ( signal_18691 ) ) ;
    buf_clk cell_4002 ( .C ( clk ), .D ( signal_18694 ), .Q ( signal_18695 ) ) ;
    buf_clk cell_4016 ( .C ( clk ), .D ( signal_18708 ), .Q ( signal_18709 ) ) ;
    buf_clk cell_4020 ( .C ( clk ), .D ( signal_18712 ), .Q ( signal_18713 ) ) ;
    buf_clk cell_4024 ( .C ( clk ), .D ( signal_18716 ), .Q ( signal_18717 ) ) ;
    buf_clk cell_4028 ( .C ( clk ), .D ( signal_18720 ), .Q ( signal_18721 ) ) ;
    buf_clk cell_4032 ( .C ( clk ), .D ( signal_18724 ), .Q ( signal_18725 ) ) ;
    buf_clk cell_4036 ( .C ( clk ), .D ( signal_18728 ), .Q ( signal_18729 ) ) ;
    buf_clk cell_4040 ( .C ( clk ), .D ( signal_18732 ), .Q ( signal_18733 ) ) ;
    buf_clk cell_4044 ( .C ( clk ), .D ( signal_18736 ), .Q ( signal_18737 ) ) ;
    buf_clk cell_4048 ( .C ( clk ), .D ( signal_18740 ), .Q ( signal_18741 ) ) ;
    buf_clk cell_4052 ( .C ( clk ), .D ( signal_18744 ), .Q ( signal_18745 ) ) ;
    buf_clk cell_4056 ( .C ( clk ), .D ( signal_18748 ), .Q ( signal_18749 ) ) ;
    buf_clk cell_4060 ( .C ( clk ), .D ( signal_18752 ), .Q ( signal_18753 ) ) ;
    buf_clk cell_4064 ( .C ( clk ), .D ( signal_18756 ), .Q ( signal_18757 ) ) ;
    buf_clk cell_4068 ( .C ( clk ), .D ( signal_18760 ), .Q ( signal_18761 ) ) ;
    buf_clk cell_4072 ( .C ( clk ), .D ( signal_18764 ), .Q ( signal_18765 ) ) ;
    buf_clk cell_4080 ( .C ( clk ), .D ( signal_18772 ), .Q ( signal_18773 ) ) ;
    buf_clk cell_4088 ( .C ( clk ), .D ( signal_18780 ), .Q ( signal_18781 ) ) ;
    buf_clk cell_4096 ( .C ( clk ), .D ( signal_18788 ), .Q ( signal_18789 ) ) ;
    buf_clk cell_4104 ( .C ( clk ), .D ( signal_18796 ), .Q ( signal_18797 ) ) ;
    buf_clk cell_4112 ( .C ( clk ), .D ( signal_18804 ), .Q ( signal_18805 ) ) ;
    buf_clk cell_4136 ( .C ( clk ), .D ( signal_18828 ), .Q ( signal_18829 ) ) ;
    buf_clk cell_4140 ( .C ( clk ), .D ( signal_18832 ), .Q ( signal_18833 ) ) ;
    buf_clk cell_4144 ( .C ( clk ), .D ( signal_18836 ), .Q ( signal_18837 ) ) ;
    buf_clk cell_4148 ( .C ( clk ), .D ( signal_18840 ), .Q ( signal_18841 ) ) ;
    buf_clk cell_4152 ( .C ( clk ), .D ( signal_18844 ), .Q ( signal_18845 ) ) ;
    buf_clk cell_4176 ( .C ( clk ), .D ( signal_18868 ), .Q ( signal_18869 ) ) ;
    buf_clk cell_4180 ( .C ( clk ), .D ( signal_18872 ), .Q ( signal_18873 ) ) ;
    buf_clk cell_4184 ( .C ( clk ), .D ( signal_18876 ), .Q ( signal_18877 ) ) ;
    buf_clk cell_4188 ( .C ( clk ), .D ( signal_18880 ), .Q ( signal_18881 ) ) ;
    buf_clk cell_4192 ( .C ( clk ), .D ( signal_18884 ), .Q ( signal_18885 ) ) ;
    buf_clk cell_4246 ( .C ( clk ), .D ( signal_18938 ), .Q ( signal_18939 ) ) ;
    buf_clk cell_4250 ( .C ( clk ), .D ( signal_18942 ), .Q ( signal_18943 ) ) ;
    buf_clk cell_4254 ( .C ( clk ), .D ( signal_18946 ), .Q ( signal_18947 ) ) ;
    buf_clk cell_4258 ( .C ( clk ), .D ( signal_18950 ), .Q ( signal_18951 ) ) ;
    buf_clk cell_4262 ( .C ( clk ), .D ( signal_18954 ), .Q ( signal_18955 ) ) ;
    buf_clk cell_4306 ( .C ( clk ), .D ( signal_18998 ), .Q ( signal_18999 ) ) ;
    buf_clk cell_4310 ( .C ( clk ), .D ( signal_19002 ), .Q ( signal_19003 ) ) ;
    buf_clk cell_4314 ( .C ( clk ), .D ( signal_19006 ), .Q ( signal_19007 ) ) ;
    buf_clk cell_4318 ( .C ( clk ), .D ( signal_19010 ), .Q ( signal_19011 ) ) ;
    buf_clk cell_4322 ( .C ( clk ), .D ( signal_19014 ), .Q ( signal_19015 ) ) ;
    buf_clk cell_4346 ( .C ( clk ), .D ( signal_19038 ), .Q ( signal_19039 ) ) ;
    buf_clk cell_4350 ( .C ( clk ), .D ( signal_19042 ), .Q ( signal_19043 ) ) ;
    buf_clk cell_4354 ( .C ( clk ), .D ( signal_19046 ), .Q ( signal_19047 ) ) ;
    buf_clk cell_4358 ( .C ( clk ), .D ( signal_19050 ), .Q ( signal_19051 ) ) ;
    buf_clk cell_4362 ( .C ( clk ), .D ( signal_19054 ), .Q ( signal_19055 ) ) ;
    buf_clk cell_4366 ( .C ( clk ), .D ( signal_19058 ), .Q ( signal_19059 ) ) ;
    buf_clk cell_4370 ( .C ( clk ), .D ( signal_19062 ), .Q ( signal_19063 ) ) ;
    buf_clk cell_4374 ( .C ( clk ), .D ( signal_19066 ), .Q ( signal_19067 ) ) ;
    buf_clk cell_4378 ( .C ( clk ), .D ( signal_19070 ), .Q ( signal_19071 ) ) ;
    buf_clk cell_4382 ( .C ( clk ), .D ( signal_19074 ), .Q ( signal_19075 ) ) ;
    buf_clk cell_4386 ( .C ( clk ), .D ( signal_19078 ), .Q ( signal_19079 ) ) ;
    buf_clk cell_4390 ( .C ( clk ), .D ( signal_19082 ), .Q ( signal_19083 ) ) ;
    buf_clk cell_4394 ( .C ( clk ), .D ( signal_19086 ), .Q ( signal_19087 ) ) ;
    buf_clk cell_4398 ( .C ( clk ), .D ( signal_19090 ), .Q ( signal_19091 ) ) ;
    buf_clk cell_4402 ( .C ( clk ), .D ( signal_19094 ), .Q ( signal_19095 ) ) ;
    buf_clk cell_4406 ( .C ( clk ), .D ( signal_19098 ), .Q ( signal_19099 ) ) ;
    buf_clk cell_4410 ( .C ( clk ), .D ( signal_19102 ), .Q ( signal_19103 ) ) ;
    buf_clk cell_4414 ( .C ( clk ), .D ( signal_19106 ), .Q ( signal_19107 ) ) ;
    buf_clk cell_4418 ( .C ( clk ), .D ( signal_19110 ), .Q ( signal_19111 ) ) ;
    buf_clk cell_4422 ( .C ( clk ), .D ( signal_19114 ), .Q ( signal_19115 ) ) ;
    buf_clk cell_4476 ( .C ( clk ), .D ( signal_19168 ), .Q ( signal_19169 ) ) ;
    buf_clk cell_4480 ( .C ( clk ), .D ( signal_19172 ), .Q ( signal_19173 ) ) ;
    buf_clk cell_4484 ( .C ( clk ), .D ( signal_19176 ), .Q ( signal_19177 ) ) ;
    buf_clk cell_4488 ( .C ( clk ), .D ( signal_19180 ), .Q ( signal_19181 ) ) ;
    buf_clk cell_4492 ( .C ( clk ), .D ( signal_19184 ), .Q ( signal_19185 ) ) ;
    buf_clk cell_4496 ( .C ( clk ), .D ( signal_19188 ), .Q ( signal_19189 ) ) ;
    buf_clk cell_4500 ( .C ( clk ), .D ( signal_19192 ), .Q ( signal_19193 ) ) ;
    buf_clk cell_4504 ( .C ( clk ), .D ( signal_19196 ), .Q ( signal_19197 ) ) ;
    buf_clk cell_4508 ( .C ( clk ), .D ( signal_19200 ), .Q ( signal_19201 ) ) ;
    buf_clk cell_4512 ( .C ( clk ), .D ( signal_19204 ), .Q ( signal_19205 ) ) ;
    buf_clk cell_4516 ( .C ( clk ), .D ( signal_19208 ), .Q ( signal_19209 ) ) ;
    buf_clk cell_4520 ( .C ( clk ), .D ( signal_19212 ), .Q ( signal_19213 ) ) ;
    buf_clk cell_4524 ( .C ( clk ), .D ( signal_19216 ), .Q ( signal_19217 ) ) ;
    buf_clk cell_4528 ( .C ( clk ), .D ( signal_19220 ), .Q ( signal_19221 ) ) ;
    buf_clk cell_4532 ( .C ( clk ), .D ( signal_19224 ), .Q ( signal_19225 ) ) ;
    buf_clk cell_4546 ( .C ( clk ), .D ( signal_19238 ), .Q ( signal_19239 ) ) ;
    buf_clk cell_4550 ( .C ( clk ), .D ( signal_19242 ), .Q ( signal_19243 ) ) ;
    buf_clk cell_4554 ( .C ( clk ), .D ( signal_19246 ), .Q ( signal_19247 ) ) ;
    buf_clk cell_4558 ( .C ( clk ), .D ( signal_19250 ), .Q ( signal_19251 ) ) ;
    buf_clk cell_4562 ( .C ( clk ), .D ( signal_19254 ), .Q ( signal_19255 ) ) ;
    buf_clk cell_4616 ( .C ( clk ), .D ( signal_19308 ), .Q ( signal_19309 ) ) ;
    buf_clk cell_4620 ( .C ( clk ), .D ( signal_19312 ), .Q ( signal_19313 ) ) ;
    buf_clk cell_4624 ( .C ( clk ), .D ( signal_19316 ), .Q ( signal_19317 ) ) ;
    buf_clk cell_4628 ( .C ( clk ), .D ( signal_19320 ), .Q ( signal_19321 ) ) ;
    buf_clk cell_4632 ( .C ( clk ), .D ( signal_19324 ), .Q ( signal_19325 ) ) ;
    buf_clk cell_4636 ( .C ( clk ), .D ( signal_19328 ), .Q ( signal_19329 ) ) ;
    buf_clk cell_4640 ( .C ( clk ), .D ( signal_19332 ), .Q ( signal_19333 ) ) ;
    buf_clk cell_4644 ( .C ( clk ), .D ( signal_19336 ), .Q ( signal_19337 ) ) ;
    buf_clk cell_4648 ( .C ( clk ), .D ( signal_19340 ), .Q ( signal_19341 ) ) ;
    buf_clk cell_4652 ( .C ( clk ), .D ( signal_19344 ), .Q ( signal_19345 ) ) ;
    buf_clk cell_4666 ( .C ( clk ), .D ( signal_19358 ), .Q ( signal_19359 ) ) ;
    buf_clk cell_4670 ( .C ( clk ), .D ( signal_19362 ), .Q ( signal_19363 ) ) ;
    buf_clk cell_4674 ( .C ( clk ), .D ( signal_19366 ), .Q ( signal_19367 ) ) ;
    buf_clk cell_4678 ( .C ( clk ), .D ( signal_19370 ), .Q ( signal_19371 ) ) ;
    buf_clk cell_4682 ( .C ( clk ), .D ( signal_19374 ), .Q ( signal_19375 ) ) ;
    buf_clk cell_4706 ( .C ( clk ), .D ( signal_19398 ), .Q ( signal_19399 ) ) ;
    buf_clk cell_4710 ( .C ( clk ), .D ( signal_19402 ), .Q ( signal_19403 ) ) ;
    buf_clk cell_4714 ( .C ( clk ), .D ( signal_19406 ), .Q ( signal_19407 ) ) ;
    buf_clk cell_4718 ( .C ( clk ), .D ( signal_19410 ), .Q ( signal_19411 ) ) ;
    buf_clk cell_4722 ( .C ( clk ), .D ( signal_19414 ), .Q ( signal_19415 ) ) ;
    buf_clk cell_4726 ( .C ( clk ), .D ( signal_19418 ), .Q ( signal_19419 ) ) ;
    buf_clk cell_4730 ( .C ( clk ), .D ( signal_19422 ), .Q ( signal_19423 ) ) ;
    buf_clk cell_4734 ( .C ( clk ), .D ( signal_19426 ), .Q ( signal_19427 ) ) ;
    buf_clk cell_4738 ( .C ( clk ), .D ( signal_19430 ), .Q ( signal_19431 ) ) ;
    buf_clk cell_4742 ( .C ( clk ), .D ( signal_19434 ), .Q ( signal_19435 ) ) ;
    buf_clk cell_4746 ( .C ( clk ), .D ( signal_19438 ), .Q ( signal_19439 ) ) ;
    buf_clk cell_4750 ( .C ( clk ), .D ( signal_19442 ), .Q ( signal_19443 ) ) ;
    buf_clk cell_4754 ( .C ( clk ), .D ( signal_19446 ), .Q ( signal_19447 ) ) ;
    buf_clk cell_4758 ( .C ( clk ), .D ( signal_19450 ), .Q ( signal_19451 ) ) ;
    buf_clk cell_4762 ( .C ( clk ), .D ( signal_19454 ), .Q ( signal_19455 ) ) ;
    buf_clk cell_4776 ( .C ( clk ), .D ( signal_19468 ), .Q ( signal_19469 ) ) ;
    buf_clk cell_4780 ( .C ( clk ), .D ( signal_19472 ), .Q ( signal_19473 ) ) ;
    buf_clk cell_4784 ( .C ( clk ), .D ( signal_19476 ), .Q ( signal_19477 ) ) ;
    buf_clk cell_4788 ( .C ( clk ), .D ( signal_19480 ), .Q ( signal_19481 ) ) ;
    buf_clk cell_4792 ( .C ( clk ), .D ( signal_19484 ), .Q ( signal_19485 ) ) ;
    buf_clk cell_4796 ( .C ( clk ), .D ( signal_19488 ), .Q ( signal_19489 ) ) ;
    buf_clk cell_4800 ( .C ( clk ), .D ( signal_19492 ), .Q ( signal_19493 ) ) ;
    buf_clk cell_4804 ( .C ( clk ), .D ( signal_19496 ), .Q ( signal_19497 ) ) ;
    buf_clk cell_4808 ( .C ( clk ), .D ( signal_19500 ), .Q ( signal_19501 ) ) ;
    buf_clk cell_4812 ( .C ( clk ), .D ( signal_19504 ), .Q ( signal_19505 ) ) ;
    buf_clk cell_4826 ( .C ( clk ), .D ( signal_19518 ), .Q ( signal_19519 ) ) ;
    buf_clk cell_4830 ( .C ( clk ), .D ( signal_19522 ), .Q ( signal_19523 ) ) ;
    buf_clk cell_4834 ( .C ( clk ), .D ( signal_19526 ), .Q ( signal_19527 ) ) ;
    buf_clk cell_4838 ( .C ( clk ), .D ( signal_19530 ), .Q ( signal_19531 ) ) ;
    buf_clk cell_4842 ( .C ( clk ), .D ( signal_19534 ), .Q ( signal_19535 ) ) ;
    buf_clk cell_4876 ( .C ( clk ), .D ( signal_19568 ), .Q ( signal_19569 ) ) ;
    buf_clk cell_4880 ( .C ( clk ), .D ( signal_19572 ), .Q ( signal_19573 ) ) ;
    buf_clk cell_4884 ( .C ( clk ), .D ( signal_19576 ), .Q ( signal_19577 ) ) ;
    buf_clk cell_4888 ( .C ( clk ), .D ( signal_19580 ), .Q ( signal_19581 ) ) ;
    buf_clk cell_4892 ( .C ( clk ), .D ( signal_19584 ), .Q ( signal_19585 ) ) ;
    buf_clk cell_4906 ( .C ( clk ), .D ( signal_19598 ), .Q ( signal_19599 ) ) ;
    buf_clk cell_4912 ( .C ( clk ), .D ( signal_19604 ), .Q ( signal_19605 ) ) ;
    buf_clk cell_4918 ( .C ( clk ), .D ( signal_19610 ), .Q ( signal_19611 ) ) ;
    buf_clk cell_4924 ( .C ( clk ), .D ( signal_19616 ), .Q ( signal_19617 ) ) ;
    buf_clk cell_4930 ( .C ( clk ), .D ( signal_19622 ), .Q ( signal_19623 ) ) ;
    buf_clk cell_4936 ( .C ( clk ), .D ( signal_19628 ), .Q ( signal_19629 ) ) ;
    buf_clk cell_4942 ( .C ( clk ), .D ( signal_19634 ), .Q ( signal_19635 ) ) ;
    buf_clk cell_4948 ( .C ( clk ), .D ( signal_19640 ), .Q ( signal_19641 ) ) ;
    buf_clk cell_4954 ( .C ( clk ), .D ( signal_19646 ), .Q ( signal_19647 ) ) ;
    buf_clk cell_4960 ( .C ( clk ), .D ( signal_19652 ), .Q ( signal_19653 ) ) ;
    buf_clk cell_4966 ( .C ( clk ), .D ( signal_19658 ), .Q ( signal_19659 ) ) ;
    buf_clk cell_4972 ( .C ( clk ), .D ( signal_19664 ), .Q ( signal_19665 ) ) ;
    buf_clk cell_4978 ( .C ( clk ), .D ( signal_19670 ), .Q ( signal_19671 ) ) ;
    buf_clk cell_4984 ( .C ( clk ), .D ( signal_19676 ), .Q ( signal_19677 ) ) ;
    buf_clk cell_4990 ( .C ( clk ), .D ( signal_19682 ), .Q ( signal_19683 ) ) ;
    buf_clk cell_5016 ( .C ( clk ), .D ( signal_19708 ), .Q ( signal_19709 ) ) ;
    buf_clk cell_5022 ( .C ( clk ), .D ( signal_19714 ), .Q ( signal_19715 ) ) ;
    buf_clk cell_5028 ( .C ( clk ), .D ( signal_19720 ), .Q ( signal_19721 ) ) ;
    buf_clk cell_5034 ( .C ( clk ), .D ( signal_19726 ), .Q ( signal_19727 ) ) ;
    buf_clk cell_5040 ( .C ( clk ), .D ( signal_19732 ), .Q ( signal_19733 ) ) ;
    buf_clk cell_5146 ( .C ( clk ), .D ( signal_19838 ), .Q ( signal_19839 ) ) ;
    buf_clk cell_5152 ( .C ( clk ), .D ( signal_19844 ), .Q ( signal_19845 ) ) ;
    buf_clk cell_5158 ( .C ( clk ), .D ( signal_19850 ), .Q ( signal_19851 ) ) ;
    buf_clk cell_5164 ( .C ( clk ), .D ( signal_19856 ), .Q ( signal_19857 ) ) ;
    buf_clk cell_5170 ( .C ( clk ), .D ( signal_19862 ), .Q ( signal_19863 ) ) ;
    buf_clk cell_5296 ( .C ( clk ), .D ( signal_19988 ), .Q ( signal_19989 ) ) ;
    buf_clk cell_5302 ( .C ( clk ), .D ( signal_19994 ), .Q ( signal_19995 ) ) ;
    buf_clk cell_5308 ( .C ( clk ), .D ( signal_20000 ), .Q ( signal_20001 ) ) ;
    buf_clk cell_5314 ( .C ( clk ), .D ( signal_20006 ), .Q ( signal_20007 ) ) ;
    buf_clk cell_5320 ( .C ( clk ), .D ( signal_20012 ), .Q ( signal_20013 ) ) ;
    buf_clk cell_5376 ( .C ( clk ), .D ( signal_20068 ), .Q ( signal_20069 ) ) ;
    buf_clk cell_5382 ( .C ( clk ), .D ( signal_20074 ), .Q ( signal_20075 ) ) ;
    buf_clk cell_5388 ( .C ( clk ), .D ( signal_20080 ), .Q ( signal_20081 ) ) ;
    buf_clk cell_5394 ( .C ( clk ), .D ( signal_20086 ), .Q ( signal_20087 ) ) ;
    buf_clk cell_5400 ( .C ( clk ), .D ( signal_20092 ), .Q ( signal_20093 ) ) ;
    buf_clk cell_5516 ( .C ( clk ), .D ( signal_20208 ), .Q ( signal_20209 ) ) ;
    buf_clk cell_5522 ( .C ( clk ), .D ( signal_20214 ), .Q ( signal_20215 ) ) ;
    buf_clk cell_5528 ( .C ( clk ), .D ( signal_20220 ), .Q ( signal_20221 ) ) ;
    buf_clk cell_5534 ( .C ( clk ), .D ( signal_20226 ), .Q ( signal_20227 ) ) ;
    buf_clk cell_5540 ( .C ( clk ), .D ( signal_20232 ), .Q ( signal_20233 ) ) ;
    buf_clk cell_5566 ( .C ( clk ), .D ( signal_20258 ), .Q ( signal_20259 ) ) ;
    buf_clk cell_5572 ( .C ( clk ), .D ( signal_20264 ), .Q ( signal_20265 ) ) ;
    buf_clk cell_5578 ( .C ( clk ), .D ( signal_20270 ), .Q ( signal_20271 ) ) ;
    buf_clk cell_5584 ( .C ( clk ), .D ( signal_20276 ), .Q ( signal_20277 ) ) ;
    buf_clk cell_5590 ( .C ( clk ), .D ( signal_20282 ), .Q ( signal_20283 ) ) ;
    buf_clk cell_5706 ( .C ( clk ), .D ( signal_20398 ), .Q ( signal_20399 ) ) ;
    buf_clk cell_5712 ( .C ( clk ), .D ( signal_20404 ), .Q ( signal_20405 ) ) ;
    buf_clk cell_5718 ( .C ( clk ), .D ( signal_20410 ), .Q ( signal_20411 ) ) ;
    buf_clk cell_5724 ( .C ( clk ), .D ( signal_20416 ), .Q ( signal_20417 ) ) ;
    buf_clk cell_5730 ( .C ( clk ), .D ( signal_20422 ), .Q ( signal_20423 ) ) ;
    buf_clk cell_5776 ( .C ( clk ), .D ( signal_20468 ), .Q ( signal_20469 ) ) ;
    buf_clk cell_5782 ( .C ( clk ), .D ( signal_20474 ), .Q ( signal_20475 ) ) ;
    buf_clk cell_5788 ( .C ( clk ), .D ( signal_20480 ), .Q ( signal_20481 ) ) ;
    buf_clk cell_5794 ( .C ( clk ), .D ( signal_20486 ), .Q ( signal_20487 ) ) ;
    buf_clk cell_5800 ( .C ( clk ), .D ( signal_20492 ), .Q ( signal_20493 ) ) ;
    buf_clk cell_5806 ( .C ( clk ), .D ( signal_20498 ), .Q ( signal_20499 ) ) ;
    buf_clk cell_5812 ( .C ( clk ), .D ( signal_20504 ), .Q ( signal_20505 ) ) ;
    buf_clk cell_5818 ( .C ( clk ), .D ( signal_20510 ), .Q ( signal_20511 ) ) ;
    buf_clk cell_5824 ( .C ( clk ), .D ( signal_20516 ), .Q ( signal_20517 ) ) ;
    buf_clk cell_5830 ( .C ( clk ), .D ( signal_20522 ), .Q ( signal_20523 ) ) ;
    buf_clk cell_5836 ( .C ( clk ), .D ( signal_20528 ), .Q ( signal_20529 ) ) ;
    buf_clk cell_5842 ( .C ( clk ), .D ( signal_20534 ), .Q ( signal_20535 ) ) ;
    buf_clk cell_5848 ( .C ( clk ), .D ( signal_20540 ), .Q ( signal_20541 ) ) ;
    buf_clk cell_5854 ( .C ( clk ), .D ( signal_20546 ), .Q ( signal_20547 ) ) ;
    buf_clk cell_5860 ( .C ( clk ), .D ( signal_20552 ), .Q ( signal_20553 ) ) ;
    buf_clk cell_5906 ( .C ( clk ), .D ( signal_20598 ), .Q ( signal_20599 ) ) ;
    buf_clk cell_5914 ( .C ( clk ), .D ( signal_20606 ), .Q ( signal_20607 ) ) ;
    buf_clk cell_5922 ( .C ( clk ), .D ( signal_20614 ), .Q ( signal_20615 ) ) ;
    buf_clk cell_5930 ( .C ( clk ), .D ( signal_20622 ), .Q ( signal_20623 ) ) ;
    buf_clk cell_5938 ( .C ( clk ), .D ( signal_20630 ), .Q ( signal_20631 ) ) ;
    buf_clk cell_6336 ( .C ( clk ), .D ( signal_21028 ), .Q ( signal_21029 ) ) ;
    buf_clk cell_6344 ( .C ( clk ), .D ( signal_21036 ), .Q ( signal_21037 ) ) ;
    buf_clk cell_6352 ( .C ( clk ), .D ( signal_21044 ), .Q ( signal_21045 ) ) ;
    buf_clk cell_6360 ( .C ( clk ), .D ( signal_21052 ), .Q ( signal_21053 ) ) ;
    buf_clk cell_6368 ( .C ( clk ), .D ( signal_21060 ), .Q ( signal_21061 ) ) ;
    buf_clk cell_6496 ( .C ( clk ), .D ( signal_21188 ), .Q ( signal_21189 ) ) ;
    buf_clk cell_6504 ( .C ( clk ), .D ( signal_21196 ), .Q ( signal_21197 ) ) ;
    buf_clk cell_6512 ( .C ( clk ), .D ( signal_21204 ), .Q ( signal_21205 ) ) ;
    buf_clk cell_6520 ( .C ( clk ), .D ( signal_21212 ), .Q ( signal_21213 ) ) ;
    buf_clk cell_6528 ( .C ( clk ), .D ( signal_21220 ), .Q ( signal_21221 ) ) ;
    buf_clk cell_6746 ( .C ( clk ), .D ( signal_21438 ), .Q ( signal_21439 ) ) ;
    buf_clk cell_6756 ( .C ( clk ), .D ( signal_21448 ), .Q ( signal_21449 ) ) ;
    buf_clk cell_6766 ( .C ( clk ), .D ( signal_21458 ), .Q ( signal_21459 ) ) ;
    buf_clk cell_6776 ( .C ( clk ), .D ( signal_21468 ), .Q ( signal_21469 ) ) ;
    buf_clk cell_6786 ( .C ( clk ), .D ( signal_21478 ), .Q ( signal_21479 ) ) ;
    buf_clk cell_6986 ( .C ( clk ), .D ( signal_21678 ), .Q ( signal_21679 ) ) ;
    buf_clk cell_6996 ( .C ( clk ), .D ( signal_21688 ), .Q ( signal_21689 ) ) ;
    buf_clk cell_7006 ( .C ( clk ), .D ( signal_21698 ), .Q ( signal_21699 ) ) ;
    buf_clk cell_7016 ( .C ( clk ), .D ( signal_21708 ), .Q ( signal_21709 ) ) ;
    buf_clk cell_7026 ( .C ( clk ), .D ( signal_21718 ), .Q ( signal_21719 ) ) ;
    buf_clk cell_7266 ( .C ( clk ), .D ( signal_21958 ), .Q ( signal_21959 ) ) ;
    buf_clk cell_7276 ( .C ( clk ), .D ( signal_21968 ), .Q ( signal_21969 ) ) ;
    buf_clk cell_7286 ( .C ( clk ), .D ( signal_21978 ), .Q ( signal_21979 ) ) ;
    buf_clk cell_7296 ( .C ( clk ), .D ( signal_21988 ), .Q ( signal_21989 ) ) ;
    buf_clk cell_7306 ( .C ( clk ), .D ( signal_21998 ), .Q ( signal_21999 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_3965 ( .C ( clk ), .D ( signal_1550 ), .Q ( signal_18658 ) ) ;
    buf_clk cell_3967 ( .C ( clk ), .D ( signal_4856 ), .Q ( signal_18660 ) ) ;
    buf_clk cell_3969 ( .C ( clk ), .D ( signal_4857 ), .Q ( signal_18662 ) ) ;
    buf_clk cell_3971 ( .C ( clk ), .D ( signal_4858 ), .Q ( signal_18664 ) ) ;
    buf_clk cell_3973 ( .C ( clk ), .D ( signal_4859 ), .Q ( signal_18666 ) ) ;
    buf_clk cell_3975 ( .C ( clk ), .D ( signal_1566 ), .Q ( signal_18668 ) ) ;
    buf_clk cell_3977 ( .C ( clk ), .D ( signal_4920 ), .Q ( signal_18670 ) ) ;
    buf_clk cell_3979 ( .C ( clk ), .D ( signal_4921 ), .Q ( signal_18672 ) ) ;
    buf_clk cell_3981 ( .C ( clk ), .D ( signal_4922 ), .Q ( signal_18674 ) ) ;
    buf_clk cell_3983 ( .C ( clk ), .D ( signal_4923 ), .Q ( signal_18676 ) ) ;
    buf_clk cell_3987 ( .C ( clk ), .D ( signal_18679 ), .Q ( signal_18680 ) ) ;
    buf_clk cell_3991 ( .C ( clk ), .D ( signal_18683 ), .Q ( signal_18684 ) ) ;
    buf_clk cell_3995 ( .C ( clk ), .D ( signal_18687 ), .Q ( signal_18688 ) ) ;
    buf_clk cell_3999 ( .C ( clk ), .D ( signal_18691 ), .Q ( signal_18692 ) ) ;
    buf_clk cell_4003 ( .C ( clk ), .D ( signal_18695 ), .Q ( signal_18696 ) ) ;
    buf_clk cell_4005 ( .C ( clk ), .D ( signal_1604 ), .Q ( signal_18698 ) ) ;
    buf_clk cell_4007 ( .C ( clk ), .D ( signal_5072 ), .Q ( signal_18700 ) ) ;
    buf_clk cell_4009 ( .C ( clk ), .D ( signal_5073 ), .Q ( signal_18702 ) ) ;
    buf_clk cell_4011 ( .C ( clk ), .D ( signal_5074 ), .Q ( signal_18704 ) ) ;
    buf_clk cell_4013 ( .C ( clk ), .D ( signal_5075 ), .Q ( signal_18706 ) ) ;
    buf_clk cell_4017 ( .C ( clk ), .D ( signal_18709 ), .Q ( signal_18710 ) ) ;
    buf_clk cell_4021 ( .C ( clk ), .D ( signal_18713 ), .Q ( signal_18714 ) ) ;
    buf_clk cell_4025 ( .C ( clk ), .D ( signal_18717 ), .Q ( signal_18718 ) ) ;
    buf_clk cell_4029 ( .C ( clk ), .D ( signal_18721 ), .Q ( signal_18722 ) ) ;
    buf_clk cell_4033 ( .C ( clk ), .D ( signal_18725 ), .Q ( signal_18726 ) ) ;
    buf_clk cell_4037 ( .C ( clk ), .D ( signal_18729 ), .Q ( signal_18730 ) ) ;
    buf_clk cell_4041 ( .C ( clk ), .D ( signal_18733 ), .Q ( signal_18734 ) ) ;
    buf_clk cell_4045 ( .C ( clk ), .D ( signal_18737 ), .Q ( signal_18738 ) ) ;
    buf_clk cell_4049 ( .C ( clk ), .D ( signal_18741 ), .Q ( signal_18742 ) ) ;
    buf_clk cell_4053 ( .C ( clk ), .D ( signal_18745 ), .Q ( signal_18746 ) ) ;
    buf_clk cell_4057 ( .C ( clk ), .D ( signal_18749 ), .Q ( signal_18750 ) ) ;
    buf_clk cell_4061 ( .C ( clk ), .D ( signal_18753 ), .Q ( signal_18754 ) ) ;
    buf_clk cell_4065 ( .C ( clk ), .D ( signal_18757 ), .Q ( signal_18758 ) ) ;
    buf_clk cell_4069 ( .C ( clk ), .D ( signal_18761 ), .Q ( signal_18762 ) ) ;
    buf_clk cell_4073 ( .C ( clk ), .D ( signal_18765 ), .Q ( signal_18766 ) ) ;
    buf_clk cell_4081 ( .C ( clk ), .D ( signal_18773 ), .Q ( signal_18774 ) ) ;
    buf_clk cell_4089 ( .C ( clk ), .D ( signal_18781 ), .Q ( signal_18782 ) ) ;
    buf_clk cell_4097 ( .C ( clk ), .D ( signal_18789 ), .Q ( signal_18790 ) ) ;
    buf_clk cell_4105 ( .C ( clk ), .D ( signal_18797 ), .Q ( signal_18798 ) ) ;
    buf_clk cell_4113 ( .C ( clk ), .D ( signal_18805 ), .Q ( signal_18806 ) ) ;
    buf_clk cell_4115 ( .C ( clk ), .D ( signal_1576 ), .Q ( signal_18808 ) ) ;
    buf_clk cell_4117 ( .C ( clk ), .D ( signal_4960 ), .Q ( signal_18810 ) ) ;
    buf_clk cell_4119 ( .C ( clk ), .D ( signal_4961 ), .Q ( signal_18812 ) ) ;
    buf_clk cell_4121 ( .C ( clk ), .D ( signal_4962 ), .Q ( signal_18814 ) ) ;
    buf_clk cell_4123 ( .C ( clk ), .D ( signal_4963 ), .Q ( signal_18816 ) ) ;
    buf_clk cell_4125 ( .C ( clk ), .D ( signal_1582 ), .Q ( signal_18818 ) ) ;
    buf_clk cell_4127 ( .C ( clk ), .D ( signal_4984 ), .Q ( signal_18820 ) ) ;
    buf_clk cell_4129 ( .C ( clk ), .D ( signal_4985 ), .Q ( signal_18822 ) ) ;
    buf_clk cell_4131 ( .C ( clk ), .D ( signal_4986 ), .Q ( signal_18824 ) ) ;
    buf_clk cell_4133 ( .C ( clk ), .D ( signal_4987 ), .Q ( signal_18826 ) ) ;
    buf_clk cell_4137 ( .C ( clk ), .D ( signal_18829 ), .Q ( signal_18830 ) ) ;
    buf_clk cell_4141 ( .C ( clk ), .D ( signal_18833 ), .Q ( signal_18834 ) ) ;
    buf_clk cell_4145 ( .C ( clk ), .D ( signal_18837 ), .Q ( signal_18838 ) ) ;
    buf_clk cell_4149 ( .C ( clk ), .D ( signal_18841 ), .Q ( signal_18842 ) ) ;
    buf_clk cell_4153 ( .C ( clk ), .D ( signal_18845 ), .Q ( signal_18846 ) ) ;
    buf_clk cell_4155 ( .C ( clk ), .D ( signal_1632 ), .Q ( signal_18848 ) ) ;
    buf_clk cell_4157 ( .C ( clk ), .D ( signal_5184 ), .Q ( signal_18850 ) ) ;
    buf_clk cell_4159 ( .C ( clk ), .D ( signal_5185 ), .Q ( signal_18852 ) ) ;
    buf_clk cell_4161 ( .C ( clk ), .D ( signal_5186 ), .Q ( signal_18854 ) ) ;
    buf_clk cell_4163 ( .C ( clk ), .D ( signal_5187 ), .Q ( signal_18856 ) ) ;
    buf_clk cell_4165 ( .C ( clk ), .D ( signal_1597 ), .Q ( signal_18858 ) ) ;
    buf_clk cell_4167 ( .C ( clk ), .D ( signal_5044 ), .Q ( signal_18860 ) ) ;
    buf_clk cell_4169 ( .C ( clk ), .D ( signal_5045 ), .Q ( signal_18862 ) ) ;
    buf_clk cell_4171 ( .C ( clk ), .D ( signal_5046 ), .Q ( signal_18864 ) ) ;
    buf_clk cell_4173 ( .C ( clk ), .D ( signal_5047 ), .Q ( signal_18866 ) ) ;
    buf_clk cell_4177 ( .C ( clk ), .D ( signal_18869 ), .Q ( signal_18870 ) ) ;
    buf_clk cell_4181 ( .C ( clk ), .D ( signal_18873 ), .Q ( signal_18874 ) ) ;
    buf_clk cell_4185 ( .C ( clk ), .D ( signal_18877 ), .Q ( signal_18878 ) ) ;
    buf_clk cell_4189 ( .C ( clk ), .D ( signal_18881 ), .Q ( signal_18882 ) ) ;
    buf_clk cell_4193 ( .C ( clk ), .D ( signal_18885 ), .Q ( signal_18886 ) ) ;
    buf_clk cell_4195 ( .C ( clk ), .D ( signal_1595 ), .Q ( signal_18888 ) ) ;
    buf_clk cell_4197 ( .C ( clk ), .D ( signal_5036 ), .Q ( signal_18890 ) ) ;
    buf_clk cell_4199 ( .C ( clk ), .D ( signal_5037 ), .Q ( signal_18892 ) ) ;
    buf_clk cell_4201 ( .C ( clk ), .D ( signal_5038 ), .Q ( signal_18894 ) ) ;
    buf_clk cell_4203 ( .C ( clk ), .D ( signal_5039 ), .Q ( signal_18896 ) ) ;
    buf_clk cell_4205 ( .C ( clk ), .D ( signal_1551 ), .Q ( signal_18898 ) ) ;
    buf_clk cell_4207 ( .C ( clk ), .D ( signal_4860 ), .Q ( signal_18900 ) ) ;
    buf_clk cell_4209 ( .C ( clk ), .D ( signal_4861 ), .Q ( signal_18902 ) ) ;
    buf_clk cell_4211 ( .C ( clk ), .D ( signal_4862 ), .Q ( signal_18904 ) ) ;
    buf_clk cell_4213 ( .C ( clk ), .D ( signal_4863 ), .Q ( signal_18906 ) ) ;
    buf_clk cell_4215 ( .C ( clk ), .D ( signal_1613 ), .Q ( signal_18908 ) ) ;
    buf_clk cell_4217 ( .C ( clk ), .D ( signal_5108 ), .Q ( signal_18910 ) ) ;
    buf_clk cell_4219 ( .C ( clk ), .D ( signal_5109 ), .Q ( signal_18912 ) ) ;
    buf_clk cell_4221 ( .C ( clk ), .D ( signal_5110 ), .Q ( signal_18914 ) ) ;
    buf_clk cell_4223 ( .C ( clk ), .D ( signal_5111 ), .Q ( signal_18916 ) ) ;
    buf_clk cell_4225 ( .C ( clk ), .D ( signal_1690 ), .Q ( signal_18918 ) ) ;
    buf_clk cell_4227 ( .C ( clk ), .D ( signal_5416 ), .Q ( signal_18920 ) ) ;
    buf_clk cell_4229 ( .C ( clk ), .D ( signal_5417 ), .Q ( signal_18922 ) ) ;
    buf_clk cell_4231 ( .C ( clk ), .D ( signal_5418 ), .Q ( signal_18924 ) ) ;
    buf_clk cell_4233 ( .C ( clk ), .D ( signal_5419 ), .Q ( signal_18926 ) ) ;
    buf_clk cell_4235 ( .C ( clk ), .D ( signal_1555 ), .Q ( signal_18928 ) ) ;
    buf_clk cell_4237 ( .C ( clk ), .D ( signal_4876 ), .Q ( signal_18930 ) ) ;
    buf_clk cell_4239 ( .C ( clk ), .D ( signal_4877 ), .Q ( signal_18932 ) ) ;
    buf_clk cell_4241 ( .C ( clk ), .D ( signal_4878 ), .Q ( signal_18934 ) ) ;
    buf_clk cell_4243 ( .C ( clk ), .D ( signal_4879 ), .Q ( signal_18936 ) ) ;
    buf_clk cell_4247 ( .C ( clk ), .D ( signal_18939 ), .Q ( signal_18940 ) ) ;
    buf_clk cell_4251 ( .C ( clk ), .D ( signal_18943 ), .Q ( signal_18944 ) ) ;
    buf_clk cell_4255 ( .C ( clk ), .D ( signal_18947 ), .Q ( signal_18948 ) ) ;
    buf_clk cell_4259 ( .C ( clk ), .D ( signal_18951 ), .Q ( signal_18952 ) ) ;
    buf_clk cell_4263 ( .C ( clk ), .D ( signal_18955 ), .Q ( signal_18956 ) ) ;
    buf_clk cell_4265 ( .C ( clk ), .D ( signal_1562 ), .Q ( signal_18958 ) ) ;
    buf_clk cell_4267 ( .C ( clk ), .D ( signal_4904 ), .Q ( signal_18960 ) ) ;
    buf_clk cell_4269 ( .C ( clk ), .D ( signal_4905 ), .Q ( signal_18962 ) ) ;
    buf_clk cell_4271 ( .C ( clk ), .D ( signal_4906 ), .Q ( signal_18964 ) ) ;
    buf_clk cell_4273 ( .C ( clk ), .D ( signal_4907 ), .Q ( signal_18966 ) ) ;
    buf_clk cell_4275 ( .C ( clk ), .D ( signal_1694 ), .Q ( signal_18968 ) ) ;
    buf_clk cell_4277 ( .C ( clk ), .D ( signal_5432 ), .Q ( signal_18970 ) ) ;
    buf_clk cell_4279 ( .C ( clk ), .D ( signal_5433 ), .Q ( signal_18972 ) ) ;
    buf_clk cell_4281 ( .C ( clk ), .D ( signal_5434 ), .Q ( signal_18974 ) ) ;
    buf_clk cell_4283 ( .C ( clk ), .D ( signal_5435 ), .Q ( signal_18976 ) ) ;
    buf_clk cell_4285 ( .C ( clk ), .D ( signal_1636 ), .Q ( signal_18978 ) ) ;
    buf_clk cell_4287 ( .C ( clk ), .D ( signal_5200 ), .Q ( signal_18980 ) ) ;
    buf_clk cell_4289 ( .C ( clk ), .D ( signal_5201 ), .Q ( signal_18982 ) ) ;
    buf_clk cell_4291 ( .C ( clk ), .D ( signal_5202 ), .Q ( signal_18984 ) ) ;
    buf_clk cell_4293 ( .C ( clk ), .D ( signal_5203 ), .Q ( signal_18986 ) ) ;
    buf_clk cell_4295 ( .C ( clk ), .D ( signal_1568 ), .Q ( signal_18988 ) ) ;
    buf_clk cell_4297 ( .C ( clk ), .D ( signal_4928 ), .Q ( signal_18990 ) ) ;
    buf_clk cell_4299 ( .C ( clk ), .D ( signal_4929 ), .Q ( signal_18992 ) ) ;
    buf_clk cell_4301 ( .C ( clk ), .D ( signal_4930 ), .Q ( signal_18994 ) ) ;
    buf_clk cell_4303 ( .C ( clk ), .D ( signal_4931 ), .Q ( signal_18996 ) ) ;
    buf_clk cell_4307 ( .C ( clk ), .D ( signal_18999 ), .Q ( signal_19000 ) ) ;
    buf_clk cell_4311 ( .C ( clk ), .D ( signal_19003 ), .Q ( signal_19004 ) ) ;
    buf_clk cell_4315 ( .C ( clk ), .D ( signal_19007 ), .Q ( signal_19008 ) ) ;
    buf_clk cell_4319 ( .C ( clk ), .D ( signal_19011 ), .Q ( signal_19012 ) ) ;
    buf_clk cell_4323 ( .C ( clk ), .D ( signal_19015 ), .Q ( signal_19016 ) ) ;
    buf_clk cell_4325 ( .C ( clk ), .D ( signal_1853 ), .Q ( signal_19018 ) ) ;
    buf_clk cell_4327 ( .C ( clk ), .D ( signal_6068 ), .Q ( signal_19020 ) ) ;
    buf_clk cell_4329 ( .C ( clk ), .D ( signal_6069 ), .Q ( signal_19022 ) ) ;
    buf_clk cell_4331 ( .C ( clk ), .D ( signal_6070 ), .Q ( signal_19024 ) ) ;
    buf_clk cell_4333 ( .C ( clk ), .D ( signal_6071 ), .Q ( signal_19026 ) ) ;
    buf_clk cell_4335 ( .C ( clk ), .D ( signal_18549 ), .Q ( signal_19028 ) ) ;
    buf_clk cell_4337 ( .C ( clk ), .D ( signal_18551 ), .Q ( signal_19030 ) ) ;
    buf_clk cell_4339 ( .C ( clk ), .D ( signal_18553 ), .Q ( signal_19032 ) ) ;
    buf_clk cell_4341 ( .C ( clk ), .D ( signal_18555 ), .Q ( signal_19034 ) ) ;
    buf_clk cell_4343 ( .C ( clk ), .D ( signal_18557 ), .Q ( signal_19036 ) ) ;
    buf_clk cell_4347 ( .C ( clk ), .D ( signal_19039 ), .Q ( signal_19040 ) ) ;
    buf_clk cell_4351 ( .C ( clk ), .D ( signal_19043 ), .Q ( signal_19044 ) ) ;
    buf_clk cell_4355 ( .C ( clk ), .D ( signal_19047 ), .Q ( signal_19048 ) ) ;
    buf_clk cell_4359 ( .C ( clk ), .D ( signal_19051 ), .Q ( signal_19052 ) ) ;
    buf_clk cell_4363 ( .C ( clk ), .D ( signal_19055 ), .Q ( signal_19056 ) ) ;
    buf_clk cell_4367 ( .C ( clk ), .D ( signal_19059 ), .Q ( signal_19060 ) ) ;
    buf_clk cell_4371 ( .C ( clk ), .D ( signal_19063 ), .Q ( signal_19064 ) ) ;
    buf_clk cell_4375 ( .C ( clk ), .D ( signal_19067 ), .Q ( signal_19068 ) ) ;
    buf_clk cell_4379 ( .C ( clk ), .D ( signal_19071 ), .Q ( signal_19072 ) ) ;
    buf_clk cell_4383 ( .C ( clk ), .D ( signal_19075 ), .Q ( signal_19076 ) ) ;
    buf_clk cell_4387 ( .C ( clk ), .D ( signal_19079 ), .Q ( signal_19080 ) ) ;
    buf_clk cell_4391 ( .C ( clk ), .D ( signal_19083 ), .Q ( signal_19084 ) ) ;
    buf_clk cell_4395 ( .C ( clk ), .D ( signal_19087 ), .Q ( signal_19088 ) ) ;
    buf_clk cell_4399 ( .C ( clk ), .D ( signal_19091 ), .Q ( signal_19092 ) ) ;
    buf_clk cell_4403 ( .C ( clk ), .D ( signal_19095 ), .Q ( signal_19096 ) ) ;
    buf_clk cell_4407 ( .C ( clk ), .D ( signal_19099 ), .Q ( signal_19100 ) ) ;
    buf_clk cell_4411 ( .C ( clk ), .D ( signal_19103 ), .Q ( signal_19104 ) ) ;
    buf_clk cell_4415 ( .C ( clk ), .D ( signal_19107 ), .Q ( signal_19108 ) ) ;
    buf_clk cell_4419 ( .C ( clk ), .D ( signal_19111 ), .Q ( signal_19112 ) ) ;
    buf_clk cell_4423 ( .C ( clk ), .D ( signal_19115 ), .Q ( signal_19116 ) ) ;
    buf_clk cell_4425 ( .C ( clk ), .D ( signal_18429 ), .Q ( signal_19118 ) ) ;
    buf_clk cell_4427 ( .C ( clk ), .D ( signal_18431 ), .Q ( signal_19120 ) ) ;
    buf_clk cell_4429 ( .C ( clk ), .D ( signal_18433 ), .Q ( signal_19122 ) ) ;
    buf_clk cell_4431 ( .C ( clk ), .D ( signal_18435 ), .Q ( signal_19124 ) ) ;
    buf_clk cell_4433 ( .C ( clk ), .D ( signal_18437 ), .Q ( signal_19126 ) ) ;
    buf_clk cell_4435 ( .C ( clk ), .D ( signal_18219 ), .Q ( signal_19128 ) ) ;
    buf_clk cell_4437 ( .C ( clk ), .D ( signal_18221 ), .Q ( signal_19130 ) ) ;
    buf_clk cell_4439 ( .C ( clk ), .D ( signal_18223 ), .Q ( signal_19132 ) ) ;
    buf_clk cell_4441 ( .C ( clk ), .D ( signal_18225 ), .Q ( signal_19134 ) ) ;
    buf_clk cell_4443 ( .C ( clk ), .D ( signal_18227 ), .Q ( signal_19136 ) ) ;
    buf_clk cell_4445 ( .C ( clk ), .D ( signal_1854 ), .Q ( signal_19138 ) ) ;
    buf_clk cell_4447 ( .C ( clk ), .D ( signal_6072 ), .Q ( signal_19140 ) ) ;
    buf_clk cell_4449 ( .C ( clk ), .D ( signal_6073 ), .Q ( signal_19142 ) ) ;
    buf_clk cell_4451 ( .C ( clk ), .D ( signal_6074 ), .Q ( signal_19144 ) ) ;
    buf_clk cell_4453 ( .C ( clk ), .D ( signal_6075 ), .Q ( signal_19146 ) ) ;
    buf_clk cell_4455 ( .C ( clk ), .D ( signal_17869 ), .Q ( signal_19148 ) ) ;
    buf_clk cell_4457 ( .C ( clk ), .D ( signal_17871 ), .Q ( signal_19150 ) ) ;
    buf_clk cell_4459 ( .C ( clk ), .D ( signal_17873 ), .Q ( signal_19152 ) ) ;
    buf_clk cell_4461 ( .C ( clk ), .D ( signal_17875 ), .Q ( signal_19154 ) ) ;
    buf_clk cell_4463 ( .C ( clk ), .D ( signal_17877 ), .Q ( signal_19156 ) ) ;
    buf_clk cell_4465 ( .C ( clk ), .D ( signal_18609 ), .Q ( signal_19158 ) ) ;
    buf_clk cell_4467 ( .C ( clk ), .D ( signal_18611 ), .Q ( signal_19160 ) ) ;
    buf_clk cell_4469 ( .C ( clk ), .D ( signal_18613 ), .Q ( signal_19162 ) ) ;
    buf_clk cell_4471 ( .C ( clk ), .D ( signal_18615 ), .Q ( signal_19164 ) ) ;
    buf_clk cell_4473 ( .C ( clk ), .D ( signal_18617 ), .Q ( signal_19166 ) ) ;
    buf_clk cell_4477 ( .C ( clk ), .D ( signal_19169 ), .Q ( signal_19170 ) ) ;
    buf_clk cell_4481 ( .C ( clk ), .D ( signal_19173 ), .Q ( signal_19174 ) ) ;
    buf_clk cell_4485 ( .C ( clk ), .D ( signal_19177 ), .Q ( signal_19178 ) ) ;
    buf_clk cell_4489 ( .C ( clk ), .D ( signal_19181 ), .Q ( signal_19182 ) ) ;
    buf_clk cell_4493 ( .C ( clk ), .D ( signal_19185 ), .Q ( signal_19186 ) ) ;
    buf_clk cell_4497 ( .C ( clk ), .D ( signal_19189 ), .Q ( signal_19190 ) ) ;
    buf_clk cell_4501 ( .C ( clk ), .D ( signal_19193 ), .Q ( signal_19194 ) ) ;
    buf_clk cell_4505 ( .C ( clk ), .D ( signal_19197 ), .Q ( signal_19198 ) ) ;
    buf_clk cell_4509 ( .C ( clk ), .D ( signal_19201 ), .Q ( signal_19202 ) ) ;
    buf_clk cell_4513 ( .C ( clk ), .D ( signal_19205 ), .Q ( signal_19206 ) ) ;
    buf_clk cell_4517 ( .C ( clk ), .D ( signal_19209 ), .Q ( signal_19210 ) ) ;
    buf_clk cell_4521 ( .C ( clk ), .D ( signal_19213 ), .Q ( signal_19214 ) ) ;
    buf_clk cell_4525 ( .C ( clk ), .D ( signal_19217 ), .Q ( signal_19218 ) ) ;
    buf_clk cell_4529 ( .C ( clk ), .D ( signal_19221 ), .Q ( signal_19222 ) ) ;
    buf_clk cell_4533 ( .C ( clk ), .D ( signal_19225 ), .Q ( signal_19226 ) ) ;
    buf_clk cell_4535 ( .C ( clk ), .D ( signal_1862 ), .Q ( signal_19228 ) ) ;
    buf_clk cell_4537 ( .C ( clk ), .D ( signal_6104 ), .Q ( signal_19230 ) ) ;
    buf_clk cell_4539 ( .C ( clk ), .D ( signal_6105 ), .Q ( signal_19232 ) ) ;
    buf_clk cell_4541 ( .C ( clk ), .D ( signal_6106 ), .Q ( signal_19234 ) ) ;
    buf_clk cell_4543 ( .C ( clk ), .D ( signal_6107 ), .Q ( signal_19236 ) ) ;
    buf_clk cell_4547 ( .C ( clk ), .D ( signal_19239 ), .Q ( signal_19240 ) ) ;
    buf_clk cell_4551 ( .C ( clk ), .D ( signal_19243 ), .Q ( signal_19244 ) ) ;
    buf_clk cell_4555 ( .C ( clk ), .D ( signal_19247 ), .Q ( signal_19248 ) ) ;
    buf_clk cell_4559 ( .C ( clk ), .D ( signal_19251 ), .Q ( signal_19252 ) ) ;
    buf_clk cell_4563 ( .C ( clk ), .D ( signal_19255 ), .Q ( signal_19256 ) ) ;
    buf_clk cell_4565 ( .C ( clk ), .D ( signal_17949 ), .Q ( signal_19258 ) ) ;
    buf_clk cell_4567 ( .C ( clk ), .D ( signal_17951 ), .Q ( signal_19260 ) ) ;
    buf_clk cell_4569 ( .C ( clk ), .D ( signal_17953 ), .Q ( signal_19262 ) ) ;
    buf_clk cell_4571 ( .C ( clk ), .D ( signal_17955 ), .Q ( signal_19264 ) ) ;
    buf_clk cell_4573 ( .C ( clk ), .D ( signal_17957 ), .Q ( signal_19266 ) ) ;
    buf_clk cell_4575 ( .C ( clk ), .D ( signal_1866 ), .Q ( signal_19268 ) ) ;
    buf_clk cell_4577 ( .C ( clk ), .D ( signal_6120 ), .Q ( signal_19270 ) ) ;
    buf_clk cell_4579 ( .C ( clk ), .D ( signal_6121 ), .Q ( signal_19272 ) ) ;
    buf_clk cell_4581 ( .C ( clk ), .D ( signal_6122 ), .Q ( signal_19274 ) ) ;
    buf_clk cell_4583 ( .C ( clk ), .D ( signal_6123 ), .Q ( signal_19276 ) ) ;
    buf_clk cell_4585 ( .C ( clk ), .D ( signal_17819 ), .Q ( signal_19278 ) ) ;
    buf_clk cell_4587 ( .C ( clk ), .D ( signal_17821 ), .Q ( signal_19280 ) ) ;
    buf_clk cell_4589 ( .C ( clk ), .D ( signal_17823 ), .Q ( signal_19282 ) ) ;
    buf_clk cell_4591 ( .C ( clk ), .D ( signal_17825 ), .Q ( signal_19284 ) ) ;
    buf_clk cell_4593 ( .C ( clk ), .D ( signal_17827 ), .Q ( signal_19286 ) ) ;
    buf_clk cell_4595 ( .C ( clk ), .D ( signal_1873 ), .Q ( signal_19288 ) ) ;
    buf_clk cell_4597 ( .C ( clk ), .D ( signal_6148 ), .Q ( signal_19290 ) ) ;
    buf_clk cell_4599 ( .C ( clk ), .D ( signal_6149 ), .Q ( signal_19292 ) ) ;
    buf_clk cell_4601 ( .C ( clk ), .D ( signal_6150 ), .Q ( signal_19294 ) ) ;
    buf_clk cell_4603 ( .C ( clk ), .D ( signal_6151 ), .Q ( signal_19296 ) ) ;
    buf_clk cell_4605 ( .C ( clk ), .D ( signal_1851 ), .Q ( signal_19298 ) ) ;
    buf_clk cell_4607 ( .C ( clk ), .D ( signal_6060 ), .Q ( signal_19300 ) ) ;
    buf_clk cell_4609 ( .C ( clk ), .D ( signal_6061 ), .Q ( signal_19302 ) ) ;
    buf_clk cell_4611 ( .C ( clk ), .D ( signal_6062 ), .Q ( signal_19304 ) ) ;
    buf_clk cell_4613 ( .C ( clk ), .D ( signal_6063 ), .Q ( signal_19306 ) ) ;
    buf_clk cell_4617 ( .C ( clk ), .D ( signal_19309 ), .Q ( signal_19310 ) ) ;
    buf_clk cell_4621 ( .C ( clk ), .D ( signal_19313 ), .Q ( signal_19314 ) ) ;
    buf_clk cell_4625 ( .C ( clk ), .D ( signal_19317 ), .Q ( signal_19318 ) ) ;
    buf_clk cell_4629 ( .C ( clk ), .D ( signal_19321 ), .Q ( signal_19322 ) ) ;
    buf_clk cell_4633 ( .C ( clk ), .D ( signal_19325 ), .Q ( signal_19326 ) ) ;
    buf_clk cell_4637 ( .C ( clk ), .D ( signal_19329 ), .Q ( signal_19330 ) ) ;
    buf_clk cell_4641 ( .C ( clk ), .D ( signal_19333 ), .Q ( signal_19334 ) ) ;
    buf_clk cell_4645 ( .C ( clk ), .D ( signal_19337 ), .Q ( signal_19338 ) ) ;
    buf_clk cell_4649 ( .C ( clk ), .D ( signal_19341 ), .Q ( signal_19342 ) ) ;
    buf_clk cell_4653 ( .C ( clk ), .D ( signal_19345 ), .Q ( signal_19346 ) ) ;
    buf_clk cell_4655 ( .C ( clk ), .D ( signal_1571 ), .Q ( signal_19348 ) ) ;
    buf_clk cell_4657 ( .C ( clk ), .D ( signal_4940 ), .Q ( signal_19350 ) ) ;
    buf_clk cell_4659 ( .C ( clk ), .D ( signal_4941 ), .Q ( signal_19352 ) ) ;
    buf_clk cell_4661 ( .C ( clk ), .D ( signal_4942 ), .Q ( signal_19354 ) ) ;
    buf_clk cell_4663 ( .C ( clk ), .D ( signal_4943 ), .Q ( signal_19356 ) ) ;
    buf_clk cell_4667 ( .C ( clk ), .D ( signal_19359 ), .Q ( signal_19360 ) ) ;
    buf_clk cell_4671 ( .C ( clk ), .D ( signal_19363 ), .Q ( signal_19364 ) ) ;
    buf_clk cell_4675 ( .C ( clk ), .D ( signal_19367 ), .Q ( signal_19368 ) ) ;
    buf_clk cell_4679 ( .C ( clk ), .D ( signal_19371 ), .Q ( signal_19372 ) ) ;
    buf_clk cell_4683 ( .C ( clk ), .D ( signal_19375 ), .Q ( signal_19376 ) ) ;
    buf_clk cell_4685 ( .C ( clk ), .D ( signal_1540 ), .Q ( signal_19378 ) ) ;
    buf_clk cell_4687 ( .C ( clk ), .D ( signal_4816 ), .Q ( signal_19380 ) ) ;
    buf_clk cell_4689 ( .C ( clk ), .D ( signal_4817 ), .Q ( signal_19382 ) ) ;
    buf_clk cell_4691 ( .C ( clk ), .D ( signal_4818 ), .Q ( signal_19384 ) ) ;
    buf_clk cell_4693 ( .C ( clk ), .D ( signal_4819 ), .Q ( signal_19386 ) ) ;
    buf_clk cell_4695 ( .C ( clk ), .D ( signal_1872 ), .Q ( signal_19388 ) ) ;
    buf_clk cell_4697 ( .C ( clk ), .D ( signal_6144 ), .Q ( signal_19390 ) ) ;
    buf_clk cell_4699 ( .C ( clk ), .D ( signal_6145 ), .Q ( signal_19392 ) ) ;
    buf_clk cell_4701 ( .C ( clk ), .D ( signal_6146 ), .Q ( signal_19394 ) ) ;
    buf_clk cell_4703 ( .C ( clk ), .D ( signal_6147 ), .Q ( signal_19396 ) ) ;
    buf_clk cell_4707 ( .C ( clk ), .D ( signal_19399 ), .Q ( signal_19400 ) ) ;
    buf_clk cell_4711 ( .C ( clk ), .D ( signal_19403 ), .Q ( signal_19404 ) ) ;
    buf_clk cell_4715 ( .C ( clk ), .D ( signal_19407 ), .Q ( signal_19408 ) ) ;
    buf_clk cell_4719 ( .C ( clk ), .D ( signal_19411 ), .Q ( signal_19412 ) ) ;
    buf_clk cell_4723 ( .C ( clk ), .D ( signal_19415 ), .Q ( signal_19416 ) ) ;
    buf_clk cell_4727 ( .C ( clk ), .D ( signal_19419 ), .Q ( signal_19420 ) ) ;
    buf_clk cell_4731 ( .C ( clk ), .D ( signal_19423 ), .Q ( signal_19424 ) ) ;
    buf_clk cell_4735 ( .C ( clk ), .D ( signal_19427 ), .Q ( signal_19428 ) ) ;
    buf_clk cell_4739 ( .C ( clk ), .D ( signal_19431 ), .Q ( signal_19432 ) ) ;
    buf_clk cell_4743 ( .C ( clk ), .D ( signal_19435 ), .Q ( signal_19436 ) ) ;
    buf_clk cell_4747 ( .C ( clk ), .D ( signal_19439 ), .Q ( signal_19440 ) ) ;
    buf_clk cell_4751 ( .C ( clk ), .D ( signal_19443 ), .Q ( signal_19444 ) ) ;
    buf_clk cell_4755 ( .C ( clk ), .D ( signal_19447 ), .Q ( signal_19448 ) ) ;
    buf_clk cell_4759 ( .C ( clk ), .D ( signal_19451 ), .Q ( signal_19452 ) ) ;
    buf_clk cell_4763 ( .C ( clk ), .D ( signal_19455 ), .Q ( signal_19456 ) ) ;
    buf_clk cell_4765 ( .C ( clk ), .D ( signal_1583 ), .Q ( signal_19458 ) ) ;
    buf_clk cell_4767 ( .C ( clk ), .D ( signal_4988 ), .Q ( signal_19460 ) ) ;
    buf_clk cell_4769 ( .C ( clk ), .D ( signal_4989 ), .Q ( signal_19462 ) ) ;
    buf_clk cell_4771 ( .C ( clk ), .D ( signal_4990 ), .Q ( signal_19464 ) ) ;
    buf_clk cell_4773 ( .C ( clk ), .D ( signal_4991 ), .Q ( signal_19466 ) ) ;
    buf_clk cell_4777 ( .C ( clk ), .D ( signal_19469 ), .Q ( signal_19470 ) ) ;
    buf_clk cell_4781 ( .C ( clk ), .D ( signal_19473 ), .Q ( signal_19474 ) ) ;
    buf_clk cell_4785 ( .C ( clk ), .D ( signal_19477 ), .Q ( signal_19478 ) ) ;
    buf_clk cell_4789 ( .C ( clk ), .D ( signal_19481 ), .Q ( signal_19482 ) ) ;
    buf_clk cell_4793 ( .C ( clk ), .D ( signal_19485 ), .Q ( signal_19486 ) ) ;
    buf_clk cell_4797 ( .C ( clk ), .D ( signal_19489 ), .Q ( signal_19490 ) ) ;
    buf_clk cell_4801 ( .C ( clk ), .D ( signal_19493 ), .Q ( signal_19494 ) ) ;
    buf_clk cell_4805 ( .C ( clk ), .D ( signal_19497 ), .Q ( signal_19498 ) ) ;
    buf_clk cell_4809 ( .C ( clk ), .D ( signal_19501 ), .Q ( signal_19502 ) ) ;
    buf_clk cell_4813 ( .C ( clk ), .D ( signal_19505 ), .Q ( signal_19506 ) ) ;
    buf_clk cell_4815 ( .C ( clk ), .D ( signal_1600 ), .Q ( signal_19508 ) ) ;
    buf_clk cell_4817 ( .C ( clk ), .D ( signal_5056 ), .Q ( signal_19510 ) ) ;
    buf_clk cell_4819 ( .C ( clk ), .D ( signal_5057 ), .Q ( signal_19512 ) ) ;
    buf_clk cell_4821 ( .C ( clk ), .D ( signal_5058 ), .Q ( signal_19514 ) ) ;
    buf_clk cell_4823 ( .C ( clk ), .D ( signal_5059 ), .Q ( signal_19516 ) ) ;
    buf_clk cell_4827 ( .C ( clk ), .D ( signal_19519 ), .Q ( signal_19520 ) ) ;
    buf_clk cell_4831 ( .C ( clk ), .D ( signal_19523 ), .Q ( signal_19524 ) ) ;
    buf_clk cell_4835 ( .C ( clk ), .D ( signal_19527 ), .Q ( signal_19528 ) ) ;
    buf_clk cell_4839 ( .C ( clk ), .D ( signal_19531 ), .Q ( signal_19532 ) ) ;
    buf_clk cell_4843 ( .C ( clk ), .D ( signal_19535 ), .Q ( signal_19536 ) ) ;
    buf_clk cell_4845 ( .C ( clk ), .D ( signal_1870 ), .Q ( signal_19538 ) ) ;
    buf_clk cell_4847 ( .C ( clk ), .D ( signal_6136 ), .Q ( signal_19540 ) ) ;
    buf_clk cell_4849 ( .C ( clk ), .D ( signal_6137 ), .Q ( signal_19542 ) ) ;
    buf_clk cell_4851 ( .C ( clk ), .D ( signal_6138 ), .Q ( signal_19544 ) ) ;
    buf_clk cell_4853 ( .C ( clk ), .D ( signal_6139 ), .Q ( signal_19546 ) ) ;
    buf_clk cell_4855 ( .C ( clk ), .D ( signal_1312 ), .Q ( signal_19548 ) ) ;
    buf_clk cell_4857 ( .C ( clk ), .D ( signal_3904 ), .Q ( signal_19550 ) ) ;
    buf_clk cell_4859 ( .C ( clk ), .D ( signal_3905 ), .Q ( signal_19552 ) ) ;
    buf_clk cell_4861 ( .C ( clk ), .D ( signal_3906 ), .Q ( signal_19554 ) ) ;
    buf_clk cell_4863 ( .C ( clk ), .D ( signal_3907 ), .Q ( signal_19556 ) ) ;
    buf_clk cell_4865 ( .C ( clk ), .D ( signal_17909 ), .Q ( signal_19558 ) ) ;
    buf_clk cell_4867 ( .C ( clk ), .D ( signal_17911 ), .Q ( signal_19560 ) ) ;
    buf_clk cell_4869 ( .C ( clk ), .D ( signal_17913 ), .Q ( signal_19562 ) ) ;
    buf_clk cell_4871 ( .C ( clk ), .D ( signal_17915 ), .Q ( signal_19564 ) ) ;
    buf_clk cell_4873 ( .C ( clk ), .D ( signal_17917 ), .Q ( signal_19566 ) ) ;
    buf_clk cell_4877 ( .C ( clk ), .D ( signal_19569 ), .Q ( signal_19570 ) ) ;
    buf_clk cell_4881 ( .C ( clk ), .D ( signal_19573 ), .Q ( signal_19574 ) ) ;
    buf_clk cell_4885 ( .C ( clk ), .D ( signal_19577 ), .Q ( signal_19578 ) ) ;
    buf_clk cell_4889 ( .C ( clk ), .D ( signal_19581 ), .Q ( signal_19582 ) ) ;
    buf_clk cell_4893 ( .C ( clk ), .D ( signal_19585 ), .Q ( signal_19586 ) ) ;
    buf_clk cell_4907 ( .C ( clk ), .D ( signal_19599 ), .Q ( signal_19600 ) ) ;
    buf_clk cell_4913 ( .C ( clk ), .D ( signal_19605 ), .Q ( signal_19606 ) ) ;
    buf_clk cell_4919 ( .C ( clk ), .D ( signal_19611 ), .Q ( signal_19612 ) ) ;
    buf_clk cell_4925 ( .C ( clk ), .D ( signal_19617 ), .Q ( signal_19618 ) ) ;
    buf_clk cell_4931 ( .C ( clk ), .D ( signal_19623 ), .Q ( signal_19624 ) ) ;
    buf_clk cell_4937 ( .C ( clk ), .D ( signal_19629 ), .Q ( signal_19630 ) ) ;
    buf_clk cell_4943 ( .C ( clk ), .D ( signal_19635 ), .Q ( signal_19636 ) ) ;
    buf_clk cell_4949 ( .C ( clk ), .D ( signal_19641 ), .Q ( signal_19642 ) ) ;
    buf_clk cell_4955 ( .C ( clk ), .D ( signal_19647 ), .Q ( signal_19648 ) ) ;
    buf_clk cell_4961 ( .C ( clk ), .D ( signal_19653 ), .Q ( signal_19654 ) ) ;
    buf_clk cell_4967 ( .C ( clk ), .D ( signal_19659 ), .Q ( signal_19660 ) ) ;
    buf_clk cell_4973 ( .C ( clk ), .D ( signal_19665 ), .Q ( signal_19666 ) ) ;
    buf_clk cell_4979 ( .C ( clk ), .D ( signal_19671 ), .Q ( signal_19672 ) ) ;
    buf_clk cell_4985 ( .C ( clk ), .D ( signal_19677 ), .Q ( signal_19678 ) ) ;
    buf_clk cell_4991 ( .C ( clk ), .D ( signal_19683 ), .Q ( signal_19684 ) ) ;
    buf_clk cell_4995 ( .C ( clk ), .D ( signal_1537 ), .Q ( signal_19688 ) ) ;
    buf_clk cell_4999 ( .C ( clk ), .D ( signal_4804 ), .Q ( signal_19692 ) ) ;
    buf_clk cell_5003 ( .C ( clk ), .D ( signal_4805 ), .Q ( signal_19696 ) ) ;
    buf_clk cell_5007 ( .C ( clk ), .D ( signal_4806 ), .Q ( signal_19700 ) ) ;
    buf_clk cell_5011 ( .C ( clk ), .D ( signal_4807 ), .Q ( signal_19704 ) ) ;
    buf_clk cell_5017 ( .C ( clk ), .D ( signal_19709 ), .Q ( signal_19710 ) ) ;
    buf_clk cell_5023 ( .C ( clk ), .D ( signal_19715 ), .Q ( signal_19716 ) ) ;
    buf_clk cell_5029 ( .C ( clk ), .D ( signal_19721 ), .Q ( signal_19722 ) ) ;
    buf_clk cell_5035 ( .C ( clk ), .D ( signal_19727 ), .Q ( signal_19728 ) ) ;
    buf_clk cell_5041 ( .C ( clk ), .D ( signal_19733 ), .Q ( signal_19734 ) ) ;
    buf_clk cell_5045 ( .C ( clk ), .D ( signal_1552 ), .Q ( signal_19738 ) ) ;
    buf_clk cell_5049 ( .C ( clk ), .D ( signal_4864 ), .Q ( signal_19742 ) ) ;
    buf_clk cell_5053 ( .C ( clk ), .D ( signal_4865 ), .Q ( signal_19746 ) ) ;
    buf_clk cell_5057 ( .C ( clk ), .D ( signal_4866 ), .Q ( signal_19750 ) ) ;
    buf_clk cell_5061 ( .C ( clk ), .D ( signal_4867 ), .Q ( signal_19754 ) ) ;
    buf_clk cell_5065 ( .C ( clk ), .D ( signal_1618 ), .Q ( signal_19758 ) ) ;
    buf_clk cell_5069 ( .C ( clk ), .D ( signal_5128 ), .Q ( signal_19762 ) ) ;
    buf_clk cell_5073 ( .C ( clk ), .D ( signal_5129 ), .Q ( signal_19766 ) ) ;
    buf_clk cell_5077 ( .C ( clk ), .D ( signal_5130 ), .Q ( signal_19770 ) ) ;
    buf_clk cell_5081 ( .C ( clk ), .D ( signal_5131 ), .Q ( signal_19774 ) ) ;
    buf_clk cell_5085 ( .C ( clk ), .D ( signal_1560 ), .Q ( signal_19778 ) ) ;
    buf_clk cell_5089 ( .C ( clk ), .D ( signal_4896 ), .Q ( signal_19782 ) ) ;
    buf_clk cell_5093 ( .C ( clk ), .D ( signal_4897 ), .Q ( signal_19786 ) ) ;
    buf_clk cell_5097 ( .C ( clk ), .D ( signal_4898 ), .Q ( signal_19790 ) ) ;
    buf_clk cell_5101 ( .C ( clk ), .D ( signal_4899 ), .Q ( signal_19794 ) ) ;
    buf_clk cell_5105 ( .C ( clk ), .D ( signal_1622 ), .Q ( signal_19798 ) ) ;
    buf_clk cell_5109 ( .C ( clk ), .D ( signal_5144 ), .Q ( signal_19802 ) ) ;
    buf_clk cell_5113 ( .C ( clk ), .D ( signal_5145 ), .Q ( signal_19806 ) ) ;
    buf_clk cell_5117 ( .C ( clk ), .D ( signal_5146 ), .Q ( signal_19810 ) ) ;
    buf_clk cell_5121 ( .C ( clk ), .D ( signal_5147 ), .Q ( signal_19814 ) ) ;
    buf_clk cell_5125 ( .C ( clk ), .D ( signal_1533 ), .Q ( signal_19818 ) ) ;
    buf_clk cell_5129 ( .C ( clk ), .D ( signal_4788 ), .Q ( signal_19822 ) ) ;
    buf_clk cell_5133 ( .C ( clk ), .D ( signal_4789 ), .Q ( signal_19826 ) ) ;
    buf_clk cell_5137 ( .C ( clk ), .D ( signal_4790 ), .Q ( signal_19830 ) ) ;
    buf_clk cell_5141 ( .C ( clk ), .D ( signal_4791 ), .Q ( signal_19834 ) ) ;
    buf_clk cell_5147 ( .C ( clk ), .D ( signal_19839 ), .Q ( signal_19840 ) ) ;
    buf_clk cell_5153 ( .C ( clk ), .D ( signal_19845 ), .Q ( signal_19846 ) ) ;
    buf_clk cell_5159 ( .C ( clk ), .D ( signal_19851 ), .Q ( signal_19852 ) ) ;
    buf_clk cell_5165 ( .C ( clk ), .D ( signal_19857 ), .Q ( signal_19858 ) ) ;
    buf_clk cell_5171 ( .C ( clk ), .D ( signal_19863 ), .Q ( signal_19864 ) ) ;
    buf_clk cell_5175 ( .C ( clk ), .D ( signal_17979 ), .Q ( signal_19868 ) ) ;
    buf_clk cell_5179 ( .C ( clk ), .D ( signal_17981 ), .Q ( signal_19872 ) ) ;
    buf_clk cell_5183 ( .C ( clk ), .D ( signal_17983 ), .Q ( signal_19876 ) ) ;
    buf_clk cell_5187 ( .C ( clk ), .D ( signal_17985 ), .Q ( signal_19880 ) ) ;
    buf_clk cell_5191 ( .C ( clk ), .D ( signal_17987 ), .Q ( signal_19884 ) ) ;
    buf_clk cell_5245 ( .C ( clk ), .D ( signal_1591 ), .Q ( signal_19938 ) ) ;
    buf_clk cell_5249 ( .C ( clk ), .D ( signal_5020 ), .Q ( signal_19942 ) ) ;
    buf_clk cell_5253 ( .C ( clk ), .D ( signal_5021 ), .Q ( signal_19946 ) ) ;
    buf_clk cell_5257 ( .C ( clk ), .D ( signal_5022 ), .Q ( signal_19950 ) ) ;
    buf_clk cell_5261 ( .C ( clk ), .D ( signal_5023 ), .Q ( signal_19954 ) ) ;
    buf_clk cell_5297 ( .C ( clk ), .D ( signal_19989 ), .Q ( signal_19990 ) ) ;
    buf_clk cell_5303 ( .C ( clk ), .D ( signal_19995 ), .Q ( signal_19996 ) ) ;
    buf_clk cell_5309 ( .C ( clk ), .D ( signal_20001 ), .Q ( signal_20002 ) ) ;
    buf_clk cell_5315 ( .C ( clk ), .D ( signal_20007 ), .Q ( signal_20008 ) ) ;
    buf_clk cell_5321 ( .C ( clk ), .D ( signal_20013 ), .Q ( signal_20014 ) ) ;
    buf_clk cell_5335 ( .C ( clk ), .D ( signal_1621 ), .Q ( signal_20028 ) ) ;
    buf_clk cell_5339 ( .C ( clk ), .D ( signal_5140 ), .Q ( signal_20032 ) ) ;
    buf_clk cell_5343 ( .C ( clk ), .D ( signal_5141 ), .Q ( signal_20036 ) ) ;
    buf_clk cell_5347 ( .C ( clk ), .D ( signal_5142 ), .Q ( signal_20040 ) ) ;
    buf_clk cell_5351 ( .C ( clk ), .D ( signal_5143 ), .Q ( signal_20044 ) ) ;
    buf_clk cell_5377 ( .C ( clk ), .D ( signal_20069 ), .Q ( signal_20070 ) ) ;
    buf_clk cell_5383 ( .C ( clk ), .D ( signal_20075 ), .Q ( signal_20076 ) ) ;
    buf_clk cell_5389 ( .C ( clk ), .D ( signal_20081 ), .Q ( signal_20082 ) ) ;
    buf_clk cell_5395 ( .C ( clk ), .D ( signal_20087 ), .Q ( signal_20088 ) ) ;
    buf_clk cell_5401 ( .C ( clk ), .D ( signal_20093 ), .Q ( signal_20094 ) ) ;
    buf_clk cell_5405 ( .C ( clk ), .D ( signal_18619 ), .Q ( signal_20098 ) ) ;
    buf_clk cell_5409 ( .C ( clk ), .D ( signal_18621 ), .Q ( signal_20102 ) ) ;
    buf_clk cell_5413 ( .C ( clk ), .D ( signal_18623 ), .Q ( signal_20106 ) ) ;
    buf_clk cell_5417 ( .C ( clk ), .D ( signal_18625 ), .Q ( signal_20110 ) ) ;
    buf_clk cell_5421 ( .C ( clk ), .D ( signal_18627 ), .Q ( signal_20114 ) ) ;
    buf_clk cell_5445 ( .C ( clk ), .D ( signal_1606 ), .Q ( signal_20138 ) ) ;
    buf_clk cell_5449 ( .C ( clk ), .D ( signal_5080 ), .Q ( signal_20142 ) ) ;
    buf_clk cell_5453 ( .C ( clk ), .D ( signal_5081 ), .Q ( signal_20146 ) ) ;
    buf_clk cell_5457 ( .C ( clk ), .D ( signal_5082 ), .Q ( signal_20150 ) ) ;
    buf_clk cell_5461 ( .C ( clk ), .D ( signal_5083 ), .Q ( signal_20154 ) ) ;
    buf_clk cell_5465 ( .C ( clk ), .D ( signal_1691 ), .Q ( signal_20158 ) ) ;
    buf_clk cell_5469 ( .C ( clk ), .D ( signal_5420 ), .Q ( signal_20162 ) ) ;
    buf_clk cell_5473 ( .C ( clk ), .D ( signal_5421 ), .Q ( signal_20166 ) ) ;
    buf_clk cell_5477 ( .C ( clk ), .D ( signal_5422 ), .Q ( signal_20170 ) ) ;
    buf_clk cell_5481 ( .C ( clk ), .D ( signal_5423 ), .Q ( signal_20174 ) ) ;
    buf_clk cell_5485 ( .C ( clk ), .D ( signal_1570 ), .Q ( signal_20178 ) ) ;
    buf_clk cell_5489 ( .C ( clk ), .D ( signal_4936 ), .Q ( signal_20182 ) ) ;
    buf_clk cell_5493 ( .C ( clk ), .D ( signal_4937 ), .Q ( signal_20186 ) ) ;
    buf_clk cell_5497 ( .C ( clk ), .D ( signal_4938 ), .Q ( signal_20190 ) ) ;
    buf_clk cell_5501 ( .C ( clk ), .D ( signal_4939 ), .Q ( signal_20194 ) ) ;
    buf_clk cell_5517 ( .C ( clk ), .D ( signal_20209 ), .Q ( signal_20210 ) ) ;
    buf_clk cell_5523 ( .C ( clk ), .D ( signal_20215 ), .Q ( signal_20216 ) ) ;
    buf_clk cell_5529 ( .C ( clk ), .D ( signal_20221 ), .Q ( signal_20222 ) ) ;
    buf_clk cell_5535 ( .C ( clk ), .D ( signal_20227 ), .Q ( signal_20228 ) ) ;
    buf_clk cell_5541 ( .C ( clk ), .D ( signal_20233 ), .Q ( signal_20234 ) ) ;
    buf_clk cell_5545 ( .C ( clk ), .D ( signal_1584 ), .Q ( signal_20238 ) ) ;
    buf_clk cell_5549 ( .C ( clk ), .D ( signal_4992 ), .Q ( signal_20242 ) ) ;
    buf_clk cell_5553 ( .C ( clk ), .D ( signal_4993 ), .Q ( signal_20246 ) ) ;
    buf_clk cell_5557 ( .C ( clk ), .D ( signal_4994 ), .Q ( signal_20250 ) ) ;
    buf_clk cell_5561 ( .C ( clk ), .D ( signal_4995 ), .Q ( signal_20254 ) ) ;
    buf_clk cell_5567 ( .C ( clk ), .D ( signal_20259 ), .Q ( signal_20260 ) ) ;
    buf_clk cell_5573 ( .C ( clk ), .D ( signal_20265 ), .Q ( signal_20266 ) ) ;
    buf_clk cell_5579 ( .C ( clk ), .D ( signal_20271 ), .Q ( signal_20272 ) ) ;
    buf_clk cell_5585 ( .C ( clk ), .D ( signal_20277 ), .Q ( signal_20278 ) ) ;
    buf_clk cell_5591 ( .C ( clk ), .D ( signal_20283 ), .Q ( signal_20284 ) ) ;
    buf_clk cell_5595 ( .C ( clk ), .D ( signal_1590 ), .Q ( signal_20288 ) ) ;
    buf_clk cell_5599 ( .C ( clk ), .D ( signal_5016 ), .Q ( signal_20292 ) ) ;
    buf_clk cell_5603 ( .C ( clk ), .D ( signal_5017 ), .Q ( signal_20296 ) ) ;
    buf_clk cell_5607 ( .C ( clk ), .D ( signal_5018 ), .Q ( signal_20300 ) ) ;
    buf_clk cell_5611 ( .C ( clk ), .D ( signal_5019 ), .Q ( signal_20304 ) ) ;
    buf_clk cell_5615 ( .C ( clk ), .D ( signal_1675 ), .Q ( signal_20308 ) ) ;
    buf_clk cell_5619 ( .C ( clk ), .D ( signal_5356 ), .Q ( signal_20312 ) ) ;
    buf_clk cell_5623 ( .C ( clk ), .D ( signal_5357 ), .Q ( signal_20316 ) ) ;
    buf_clk cell_5627 ( .C ( clk ), .D ( signal_5358 ), .Q ( signal_20320 ) ) ;
    buf_clk cell_5631 ( .C ( clk ), .D ( signal_5359 ), .Q ( signal_20324 ) ) ;
    buf_clk cell_5635 ( .C ( clk ), .D ( signal_1598 ), .Q ( signal_20328 ) ) ;
    buf_clk cell_5639 ( .C ( clk ), .D ( signal_5048 ), .Q ( signal_20332 ) ) ;
    buf_clk cell_5643 ( .C ( clk ), .D ( signal_5049 ), .Q ( signal_20336 ) ) ;
    buf_clk cell_5647 ( .C ( clk ), .D ( signal_5050 ), .Q ( signal_20340 ) ) ;
    buf_clk cell_5651 ( .C ( clk ), .D ( signal_5051 ), .Q ( signal_20344 ) ) ;
    buf_clk cell_5665 ( .C ( clk ), .D ( signal_1601 ), .Q ( signal_20358 ) ) ;
    buf_clk cell_5669 ( .C ( clk ), .D ( signal_5060 ), .Q ( signal_20362 ) ) ;
    buf_clk cell_5673 ( .C ( clk ), .D ( signal_5061 ), .Q ( signal_20366 ) ) ;
    buf_clk cell_5677 ( .C ( clk ), .D ( signal_5062 ), .Q ( signal_20370 ) ) ;
    buf_clk cell_5681 ( .C ( clk ), .D ( signal_5063 ), .Q ( signal_20374 ) ) ;
    buf_clk cell_5685 ( .C ( clk ), .D ( signal_1543 ), .Q ( signal_20378 ) ) ;
    buf_clk cell_5689 ( .C ( clk ), .D ( signal_4828 ), .Q ( signal_20382 ) ) ;
    buf_clk cell_5693 ( .C ( clk ), .D ( signal_4829 ), .Q ( signal_20386 ) ) ;
    buf_clk cell_5697 ( .C ( clk ), .D ( signal_4830 ), .Q ( signal_20390 ) ) ;
    buf_clk cell_5701 ( .C ( clk ), .D ( signal_4831 ), .Q ( signal_20394 ) ) ;
    buf_clk cell_5707 ( .C ( clk ), .D ( signal_20399 ), .Q ( signal_20400 ) ) ;
    buf_clk cell_5713 ( .C ( clk ), .D ( signal_20405 ), .Q ( signal_20406 ) ) ;
    buf_clk cell_5719 ( .C ( clk ), .D ( signal_20411 ), .Q ( signal_20412 ) ) ;
    buf_clk cell_5725 ( .C ( clk ), .D ( signal_20417 ), .Q ( signal_20418 ) ) ;
    buf_clk cell_5731 ( .C ( clk ), .D ( signal_20423 ), .Q ( signal_20424 ) ) ;
    buf_clk cell_5755 ( .C ( clk ), .D ( signal_1625 ), .Q ( signal_20448 ) ) ;
    buf_clk cell_5759 ( .C ( clk ), .D ( signal_5156 ), .Q ( signal_20452 ) ) ;
    buf_clk cell_5763 ( .C ( clk ), .D ( signal_5157 ), .Q ( signal_20456 ) ) ;
    buf_clk cell_5767 ( .C ( clk ), .D ( signal_5158 ), .Q ( signal_20460 ) ) ;
    buf_clk cell_5771 ( .C ( clk ), .D ( signal_5159 ), .Q ( signal_20464 ) ) ;
    buf_clk cell_5777 ( .C ( clk ), .D ( signal_20469 ), .Q ( signal_20470 ) ) ;
    buf_clk cell_5783 ( .C ( clk ), .D ( signal_20475 ), .Q ( signal_20476 ) ) ;
    buf_clk cell_5789 ( .C ( clk ), .D ( signal_20481 ), .Q ( signal_20482 ) ) ;
    buf_clk cell_5795 ( .C ( clk ), .D ( signal_20487 ), .Q ( signal_20488 ) ) ;
    buf_clk cell_5801 ( .C ( clk ), .D ( signal_20493 ), .Q ( signal_20494 ) ) ;
    buf_clk cell_5807 ( .C ( clk ), .D ( signal_20499 ), .Q ( signal_20500 ) ) ;
    buf_clk cell_5813 ( .C ( clk ), .D ( signal_20505 ), .Q ( signal_20506 ) ) ;
    buf_clk cell_5819 ( .C ( clk ), .D ( signal_20511 ), .Q ( signal_20512 ) ) ;
    buf_clk cell_5825 ( .C ( clk ), .D ( signal_20517 ), .Q ( signal_20518 ) ) ;
    buf_clk cell_5831 ( .C ( clk ), .D ( signal_20523 ), .Q ( signal_20524 ) ) ;
    buf_clk cell_5837 ( .C ( clk ), .D ( signal_20529 ), .Q ( signal_20530 ) ) ;
    buf_clk cell_5843 ( .C ( clk ), .D ( signal_20535 ), .Q ( signal_20536 ) ) ;
    buf_clk cell_5849 ( .C ( clk ), .D ( signal_20541 ), .Q ( signal_20542 ) ) ;
    buf_clk cell_5855 ( .C ( clk ), .D ( signal_20547 ), .Q ( signal_20548 ) ) ;
    buf_clk cell_5861 ( .C ( clk ), .D ( signal_20553 ), .Q ( signal_20554 ) ) ;
    buf_clk cell_5865 ( .C ( clk ), .D ( signal_18403 ), .Q ( signal_20558 ) ) ;
    buf_clk cell_5869 ( .C ( clk ), .D ( signal_18409 ), .Q ( signal_20562 ) ) ;
    buf_clk cell_5873 ( .C ( clk ), .D ( signal_18415 ), .Q ( signal_20566 ) ) ;
    buf_clk cell_5877 ( .C ( clk ), .D ( signal_18421 ), .Q ( signal_20570 ) ) ;
    buf_clk cell_5881 ( .C ( clk ), .D ( signal_18427 ), .Q ( signal_20574 ) ) ;
    buf_clk cell_5907 ( .C ( clk ), .D ( signal_20599 ), .Q ( signal_20600 ) ) ;
    buf_clk cell_5915 ( .C ( clk ), .D ( signal_20607 ), .Q ( signal_20608 ) ) ;
    buf_clk cell_5923 ( .C ( clk ), .D ( signal_20615 ), .Q ( signal_20616 ) ) ;
    buf_clk cell_5931 ( .C ( clk ), .D ( signal_20623 ), .Q ( signal_20624 ) ) ;
    buf_clk cell_5939 ( .C ( clk ), .D ( signal_20631 ), .Q ( signal_20632 ) ) ;
    buf_clk cell_5965 ( .C ( clk ), .D ( signal_1645 ), .Q ( signal_20658 ) ) ;
    buf_clk cell_5971 ( .C ( clk ), .D ( signal_5236 ), .Q ( signal_20664 ) ) ;
    buf_clk cell_5977 ( .C ( clk ), .D ( signal_5237 ), .Q ( signal_20670 ) ) ;
    buf_clk cell_5983 ( .C ( clk ), .D ( signal_5238 ), .Q ( signal_20676 ) ) ;
    buf_clk cell_5989 ( .C ( clk ), .D ( signal_5239 ), .Q ( signal_20682 ) ) ;
    buf_clk cell_5995 ( .C ( clk ), .D ( signal_1616 ), .Q ( signal_20688 ) ) ;
    buf_clk cell_6001 ( .C ( clk ), .D ( signal_5120 ), .Q ( signal_20694 ) ) ;
    buf_clk cell_6007 ( .C ( clk ), .D ( signal_5121 ), .Q ( signal_20700 ) ) ;
    buf_clk cell_6013 ( .C ( clk ), .D ( signal_5122 ), .Q ( signal_20706 ) ) ;
    buf_clk cell_6019 ( .C ( clk ), .D ( signal_5123 ), .Q ( signal_20712 ) ) ;
    buf_clk cell_6045 ( .C ( clk ), .D ( signal_1534 ), .Q ( signal_20738 ) ) ;
    buf_clk cell_6051 ( .C ( clk ), .D ( signal_4792 ), .Q ( signal_20744 ) ) ;
    buf_clk cell_6057 ( .C ( clk ), .D ( signal_4793 ), .Q ( signal_20750 ) ) ;
    buf_clk cell_6063 ( .C ( clk ), .D ( signal_4794 ), .Q ( signal_20756 ) ) ;
    buf_clk cell_6069 ( .C ( clk ), .D ( signal_4795 ), .Q ( signal_20762 ) ) ;
    buf_clk cell_6135 ( .C ( clk ), .D ( signal_1850 ), .Q ( signal_20828 ) ) ;
    buf_clk cell_6141 ( .C ( clk ), .D ( signal_6056 ), .Q ( signal_20834 ) ) ;
    buf_clk cell_6147 ( .C ( clk ), .D ( signal_6057 ), .Q ( signal_20840 ) ) ;
    buf_clk cell_6153 ( .C ( clk ), .D ( signal_6058 ), .Q ( signal_20846 ) ) ;
    buf_clk cell_6159 ( .C ( clk ), .D ( signal_6059 ), .Q ( signal_20852 ) ) ;
    buf_clk cell_6165 ( .C ( clk ), .D ( signal_1631 ), .Q ( signal_20858 ) ) ;
    buf_clk cell_6171 ( .C ( clk ), .D ( signal_5180 ), .Q ( signal_20864 ) ) ;
    buf_clk cell_6177 ( .C ( clk ), .D ( signal_5181 ), .Q ( signal_20870 ) ) ;
    buf_clk cell_6183 ( .C ( clk ), .D ( signal_5182 ), .Q ( signal_20876 ) ) ;
    buf_clk cell_6189 ( .C ( clk ), .D ( signal_5183 ), .Q ( signal_20882 ) ) ;
    buf_clk cell_6195 ( .C ( clk ), .D ( signal_1683 ), .Q ( signal_20888 ) ) ;
    buf_clk cell_6201 ( .C ( clk ), .D ( signal_5388 ), .Q ( signal_20894 ) ) ;
    buf_clk cell_6207 ( .C ( clk ), .D ( signal_5389 ), .Q ( signal_20900 ) ) ;
    buf_clk cell_6213 ( .C ( clk ), .D ( signal_5390 ), .Q ( signal_20906 ) ) ;
    buf_clk cell_6219 ( .C ( clk ), .D ( signal_5391 ), .Q ( signal_20912 ) ) ;
    buf_clk cell_6255 ( .C ( clk ), .D ( signal_1299 ), .Q ( signal_20948 ) ) ;
    buf_clk cell_6261 ( .C ( clk ), .D ( signal_3852 ), .Q ( signal_20954 ) ) ;
    buf_clk cell_6267 ( .C ( clk ), .D ( signal_3853 ), .Q ( signal_20960 ) ) ;
    buf_clk cell_6273 ( .C ( clk ), .D ( signal_3854 ), .Q ( signal_20966 ) ) ;
    buf_clk cell_6279 ( .C ( clk ), .D ( signal_3855 ), .Q ( signal_20972 ) ) ;
    buf_clk cell_6295 ( .C ( clk ), .D ( signal_1557 ), .Q ( signal_20988 ) ) ;
    buf_clk cell_6301 ( .C ( clk ), .D ( signal_4884 ), .Q ( signal_20994 ) ) ;
    buf_clk cell_6307 ( .C ( clk ), .D ( signal_4885 ), .Q ( signal_21000 ) ) ;
    buf_clk cell_6313 ( .C ( clk ), .D ( signal_4886 ), .Q ( signal_21006 ) ) ;
    buf_clk cell_6319 ( .C ( clk ), .D ( signal_4887 ), .Q ( signal_21012 ) ) ;
    buf_clk cell_6337 ( .C ( clk ), .D ( signal_21029 ), .Q ( signal_21030 ) ) ;
    buf_clk cell_6345 ( .C ( clk ), .D ( signal_21037 ), .Q ( signal_21038 ) ) ;
    buf_clk cell_6353 ( .C ( clk ), .D ( signal_21045 ), .Q ( signal_21046 ) ) ;
    buf_clk cell_6361 ( .C ( clk ), .D ( signal_21053 ), .Q ( signal_21054 ) ) ;
    buf_clk cell_6369 ( .C ( clk ), .D ( signal_21061 ), .Q ( signal_21062 ) ) ;
    buf_clk cell_6415 ( .C ( clk ), .D ( signal_1506 ), .Q ( signal_21108 ) ) ;
    buf_clk cell_6421 ( .C ( clk ), .D ( signal_4680 ), .Q ( signal_21114 ) ) ;
    buf_clk cell_6427 ( .C ( clk ), .D ( signal_4681 ), .Q ( signal_21120 ) ) ;
    buf_clk cell_6433 ( .C ( clk ), .D ( signal_4682 ), .Q ( signal_21126 ) ) ;
    buf_clk cell_6439 ( .C ( clk ), .D ( signal_4683 ), .Q ( signal_21132 ) ) ;
    buf_clk cell_6445 ( .C ( clk ), .D ( signal_1593 ), .Q ( signal_21138 ) ) ;
    buf_clk cell_6451 ( .C ( clk ), .D ( signal_5028 ), .Q ( signal_21144 ) ) ;
    buf_clk cell_6457 ( .C ( clk ), .D ( signal_5029 ), .Q ( signal_21150 ) ) ;
    buf_clk cell_6463 ( .C ( clk ), .D ( signal_5030 ), .Q ( signal_21156 ) ) ;
    buf_clk cell_6469 ( .C ( clk ), .D ( signal_5031 ), .Q ( signal_21162 ) ) ;
    buf_clk cell_6497 ( .C ( clk ), .D ( signal_21189 ), .Q ( signal_21190 ) ) ;
    buf_clk cell_6505 ( .C ( clk ), .D ( signal_21197 ), .Q ( signal_21198 ) ) ;
    buf_clk cell_6513 ( .C ( clk ), .D ( signal_21205 ), .Q ( signal_21206 ) ) ;
    buf_clk cell_6521 ( .C ( clk ), .D ( signal_21213 ), .Q ( signal_21214 ) ) ;
    buf_clk cell_6529 ( .C ( clk ), .D ( signal_21221 ), .Q ( signal_21222 ) ) ;
    buf_clk cell_6535 ( .C ( clk ), .D ( signal_1338 ), .Q ( signal_21228 ) ) ;
    buf_clk cell_6541 ( .C ( clk ), .D ( signal_4008 ), .Q ( signal_21234 ) ) ;
    buf_clk cell_6547 ( .C ( clk ), .D ( signal_4009 ), .Q ( signal_21240 ) ) ;
    buf_clk cell_6553 ( .C ( clk ), .D ( signal_4010 ), .Q ( signal_21246 ) ) ;
    buf_clk cell_6559 ( .C ( clk ), .D ( signal_4011 ), .Q ( signal_21252 ) ) ;
    buf_clk cell_6565 ( .C ( clk ), .D ( signal_17889 ), .Q ( signal_21258 ) ) ;
    buf_clk cell_6571 ( .C ( clk ), .D ( signal_17891 ), .Q ( signal_21264 ) ) ;
    buf_clk cell_6577 ( .C ( clk ), .D ( signal_17893 ), .Q ( signal_21270 ) ) ;
    buf_clk cell_6583 ( .C ( clk ), .D ( signal_17895 ), .Q ( signal_21276 ) ) ;
    buf_clk cell_6589 ( .C ( clk ), .D ( signal_17897 ), .Q ( signal_21282 ) ) ;
    buf_clk cell_6615 ( .C ( clk ), .D ( signal_18339 ), .Q ( signal_21308 ) ) ;
    buf_clk cell_6621 ( .C ( clk ), .D ( signal_18341 ), .Q ( signal_21314 ) ) ;
    buf_clk cell_6627 ( .C ( clk ), .D ( signal_18343 ), .Q ( signal_21320 ) ) ;
    buf_clk cell_6633 ( .C ( clk ), .D ( signal_18345 ), .Q ( signal_21326 ) ) ;
    buf_clk cell_6639 ( .C ( clk ), .D ( signal_18347 ), .Q ( signal_21332 ) ) ;
    buf_clk cell_6665 ( .C ( clk ), .D ( signal_1637 ), .Q ( signal_21358 ) ) ;
    buf_clk cell_6671 ( .C ( clk ), .D ( signal_5204 ), .Q ( signal_21364 ) ) ;
    buf_clk cell_6677 ( .C ( clk ), .D ( signal_5205 ), .Q ( signal_21370 ) ) ;
    buf_clk cell_6683 ( .C ( clk ), .D ( signal_5206 ), .Q ( signal_21376 ) ) ;
    buf_clk cell_6689 ( .C ( clk ), .D ( signal_5207 ), .Q ( signal_21382 ) ) ;
    buf_clk cell_6695 ( .C ( clk ), .D ( signal_1518 ), .Q ( signal_21388 ) ) ;
    buf_clk cell_6701 ( .C ( clk ), .D ( signal_4728 ), .Q ( signal_21394 ) ) ;
    buf_clk cell_6707 ( .C ( clk ), .D ( signal_4729 ), .Q ( signal_21400 ) ) ;
    buf_clk cell_6713 ( .C ( clk ), .D ( signal_4730 ), .Q ( signal_21406 ) ) ;
    buf_clk cell_6719 ( .C ( clk ), .D ( signal_4731 ), .Q ( signal_21412 ) ) ;
    buf_clk cell_6747 ( .C ( clk ), .D ( signal_21439 ), .Q ( signal_21440 ) ) ;
    buf_clk cell_6757 ( .C ( clk ), .D ( signal_21449 ), .Q ( signal_21450 ) ) ;
    buf_clk cell_6767 ( .C ( clk ), .D ( signal_21459 ), .Q ( signal_21460 ) ) ;
    buf_clk cell_6777 ( .C ( clk ), .D ( signal_21469 ), .Q ( signal_21470 ) ) ;
    buf_clk cell_6787 ( .C ( clk ), .D ( signal_21479 ), .Q ( signal_21480 ) ) ;
    buf_clk cell_6825 ( .C ( clk ), .D ( signal_1619 ), .Q ( signal_21518 ) ) ;
    buf_clk cell_6833 ( .C ( clk ), .D ( signal_5132 ), .Q ( signal_21526 ) ) ;
    buf_clk cell_6841 ( .C ( clk ), .D ( signal_5133 ), .Q ( signal_21534 ) ) ;
    buf_clk cell_6849 ( .C ( clk ), .D ( signal_5134 ), .Q ( signal_21542 ) ) ;
    buf_clk cell_6857 ( .C ( clk ), .D ( signal_5135 ), .Q ( signal_21550 ) ) ;
    buf_clk cell_6865 ( .C ( clk ), .D ( signal_1350 ), .Q ( signal_21558 ) ) ;
    buf_clk cell_6873 ( .C ( clk ), .D ( signal_4056 ), .Q ( signal_21566 ) ) ;
    buf_clk cell_6881 ( .C ( clk ), .D ( signal_4057 ), .Q ( signal_21574 ) ) ;
    buf_clk cell_6889 ( .C ( clk ), .D ( signal_4058 ), .Q ( signal_21582 ) ) ;
    buf_clk cell_6897 ( .C ( clk ), .D ( signal_4059 ), .Q ( signal_21590 ) ) ;
    buf_clk cell_6987 ( .C ( clk ), .D ( signal_21679 ), .Q ( signal_21680 ) ) ;
    buf_clk cell_6997 ( .C ( clk ), .D ( signal_21689 ), .Q ( signal_21690 ) ) ;
    buf_clk cell_7007 ( .C ( clk ), .D ( signal_21699 ), .Q ( signal_21700 ) ) ;
    buf_clk cell_7017 ( .C ( clk ), .D ( signal_21709 ), .Q ( signal_21710 ) ) ;
    buf_clk cell_7027 ( .C ( clk ), .D ( signal_21719 ), .Q ( signal_21720 ) ) ;
    buf_clk cell_7075 ( .C ( clk ), .D ( signal_1575 ), .Q ( signal_21768 ) ) ;
    buf_clk cell_7083 ( .C ( clk ), .D ( signal_4956 ), .Q ( signal_21776 ) ) ;
    buf_clk cell_7091 ( .C ( clk ), .D ( signal_4957 ), .Q ( signal_21784 ) ) ;
    buf_clk cell_7099 ( .C ( clk ), .D ( signal_4958 ), .Q ( signal_21792 ) ) ;
    buf_clk cell_7107 ( .C ( clk ), .D ( signal_4959 ), .Q ( signal_21800 ) ) ;
    buf_clk cell_7145 ( .C ( clk ), .D ( signal_1587 ), .Q ( signal_21838 ) ) ;
    buf_clk cell_7153 ( .C ( clk ), .D ( signal_5004 ), .Q ( signal_21846 ) ) ;
    buf_clk cell_7161 ( .C ( clk ), .D ( signal_5005 ), .Q ( signal_21854 ) ) ;
    buf_clk cell_7169 ( .C ( clk ), .D ( signal_5006 ), .Q ( signal_21862 ) ) ;
    buf_clk cell_7177 ( .C ( clk ), .D ( signal_5007 ), .Q ( signal_21870 ) ) ;
    buf_clk cell_7185 ( .C ( clk ), .D ( signal_1861 ), .Q ( signal_21878 ) ) ;
    buf_clk cell_7193 ( .C ( clk ), .D ( signal_6100 ), .Q ( signal_21886 ) ) ;
    buf_clk cell_7201 ( .C ( clk ), .D ( signal_6101 ), .Q ( signal_21894 ) ) ;
    buf_clk cell_7209 ( .C ( clk ), .D ( signal_6102 ), .Q ( signal_21902 ) ) ;
    buf_clk cell_7217 ( .C ( clk ), .D ( signal_6103 ), .Q ( signal_21910 ) ) ;
    buf_clk cell_7225 ( .C ( clk ), .D ( signal_1258 ), .Q ( signal_21918 ) ) ;
    buf_clk cell_7233 ( .C ( clk ), .D ( signal_3688 ), .Q ( signal_21926 ) ) ;
    buf_clk cell_7241 ( .C ( clk ), .D ( signal_3689 ), .Q ( signal_21934 ) ) ;
    buf_clk cell_7249 ( .C ( clk ), .D ( signal_3690 ), .Q ( signal_21942 ) ) ;
    buf_clk cell_7257 ( .C ( clk ), .D ( signal_3691 ), .Q ( signal_21950 ) ) ;
    buf_clk cell_7267 ( .C ( clk ), .D ( signal_21959 ), .Q ( signal_21960 ) ) ;
    buf_clk cell_7277 ( .C ( clk ), .D ( signal_21969 ), .Q ( signal_21970 ) ) ;
    buf_clk cell_7287 ( .C ( clk ), .D ( signal_21979 ), .Q ( signal_21980 ) ) ;
    buf_clk cell_7297 ( .C ( clk ), .D ( signal_21989 ), .Q ( signal_21990 ) ) ;
    buf_clk cell_7307 ( .C ( clk ), .D ( signal_21999 ), .Q ( signal_22000 ) ) ;
    buf_clk cell_7315 ( .C ( clk ), .D ( signal_17969 ), .Q ( signal_22008 ) ) ;
    buf_clk cell_7323 ( .C ( clk ), .D ( signal_17971 ), .Q ( signal_22016 ) ) ;
    buf_clk cell_7331 ( .C ( clk ), .D ( signal_17973 ), .Q ( signal_22024 ) ) ;
    buf_clk cell_7339 ( .C ( clk ), .D ( signal_17975 ), .Q ( signal_22032 ) ) ;
    buf_clk cell_7347 ( .C ( clk ), .D ( signal_17977 ), .Q ( signal_22040 ) ) ;
    buf_clk cell_7355 ( .C ( clk ), .D ( signal_1614 ), .Q ( signal_22048 ) ) ;
    buf_clk cell_7363 ( .C ( clk ), .D ( signal_5112 ), .Q ( signal_22056 ) ) ;
    buf_clk cell_7371 ( .C ( clk ), .D ( signal_5113 ), .Q ( signal_22064 ) ) ;
    buf_clk cell_7379 ( .C ( clk ), .D ( signal_5114 ), .Q ( signal_22072 ) ) ;
    buf_clk cell_7387 ( .C ( clk ), .D ( signal_5115 ), .Q ( signal_22080 ) ) ;
    buf_clk cell_7405 ( .C ( clk ), .D ( signal_1549 ), .Q ( signal_22098 ) ) ;
    buf_clk cell_7413 ( .C ( clk ), .D ( signal_4852 ), .Q ( signal_22106 ) ) ;
    buf_clk cell_7421 ( .C ( clk ), .D ( signal_4853 ), .Q ( signal_22114 ) ) ;
    buf_clk cell_7429 ( .C ( clk ), .D ( signal_4854 ), .Q ( signal_22122 ) ) ;
    buf_clk cell_7437 ( .C ( clk ), .D ( signal_4855 ), .Q ( signal_22130 ) ) ;
    buf_clk cell_7445 ( .C ( clk ), .D ( signal_1578 ), .Q ( signal_22138 ) ) ;
    buf_clk cell_7453 ( .C ( clk ), .D ( signal_4968 ), .Q ( signal_22146 ) ) ;
    buf_clk cell_7461 ( .C ( clk ), .D ( signal_4969 ), .Q ( signal_22154 ) ) ;
    buf_clk cell_7469 ( .C ( clk ), .D ( signal_4970 ), .Q ( signal_22162 ) ) ;
    buf_clk cell_7477 ( .C ( clk ), .D ( signal_4971 ), .Q ( signal_22170 ) ) ;
    buf_clk cell_7485 ( .C ( clk ), .D ( signal_1581 ), .Q ( signal_22178 ) ) ;
    buf_clk cell_7493 ( .C ( clk ), .D ( signal_4980 ), .Q ( signal_22186 ) ) ;
    buf_clk cell_7501 ( .C ( clk ), .D ( signal_4981 ), .Q ( signal_22194 ) ) ;
    buf_clk cell_7509 ( .C ( clk ), .D ( signal_4982 ), .Q ( signal_22202 ) ) ;
    buf_clk cell_7517 ( .C ( clk ), .D ( signal_4983 ), .Q ( signal_22210 ) ) ;
    buf_clk cell_7695 ( .C ( clk ), .D ( signal_1505 ), .Q ( signal_22388 ) ) ;
    buf_clk cell_7705 ( .C ( clk ), .D ( signal_4676 ), .Q ( signal_22398 ) ) ;
    buf_clk cell_7715 ( .C ( clk ), .D ( signal_4677 ), .Q ( signal_22408 ) ) ;
    buf_clk cell_7725 ( .C ( clk ), .D ( signal_4678 ), .Q ( signal_22418 ) ) ;
    buf_clk cell_7735 ( .C ( clk ), .D ( signal_4679 ), .Q ( signal_22428 ) ) ;
    buf_clk cell_7825 ( .C ( clk ), .D ( signal_1589 ), .Q ( signal_22518 ) ) ;
    buf_clk cell_7835 ( .C ( clk ), .D ( signal_5012 ), .Q ( signal_22528 ) ) ;
    buf_clk cell_7845 ( .C ( clk ), .D ( signal_5013 ), .Q ( signal_22538 ) ) ;
    buf_clk cell_7855 ( .C ( clk ), .D ( signal_5014 ), .Q ( signal_22548 ) ) ;
    buf_clk cell_7865 ( .C ( clk ), .D ( signal_5015 ), .Q ( signal_22558 ) ) ;
    buf_clk cell_8835 ( .C ( clk ), .D ( signal_1527 ), .Q ( signal_23528 ) ) ;
    buf_clk cell_8849 ( .C ( clk ), .D ( signal_4764 ), .Q ( signal_23542 ) ) ;
    buf_clk cell_8863 ( .C ( clk ), .D ( signal_4765 ), .Q ( signal_23556 ) ) ;
    buf_clk cell_8877 ( .C ( clk ), .D ( signal_4766 ), .Q ( signal_23570 ) ) ;
    buf_clk cell_8891 ( .C ( clk ), .D ( signal_4767 ), .Q ( signal_23584 ) ) ;
    buf_clk cell_8945 ( .C ( clk ), .D ( signal_1633 ), .Q ( signal_23638 ) ) ;
    buf_clk cell_8959 ( .C ( clk ), .D ( signal_5188 ), .Q ( signal_23652 ) ) ;
    buf_clk cell_8973 ( .C ( clk ), .D ( signal_5189 ), .Q ( signal_23666 ) ) ;
    buf_clk cell_8987 ( .C ( clk ), .D ( signal_5190 ), .Q ( signal_23680 ) ) ;
    buf_clk cell_9001 ( .C ( clk ), .D ( signal_5191 ), .Q ( signal_23694 ) ) ;
    buf_clk cell_9145 ( .C ( clk ), .D ( signal_1588 ), .Q ( signal_23838 ) ) ;
    buf_clk cell_9161 ( .C ( clk ), .D ( signal_5008 ), .Q ( signal_23854 ) ) ;
    buf_clk cell_9177 ( .C ( clk ), .D ( signal_5009 ), .Q ( signal_23870 ) ) ;
    buf_clk cell_9193 ( .C ( clk ), .D ( signal_5010 ), .Q ( signal_23886 ) ) ;
    buf_clk cell_9209 ( .C ( clk ), .D ( signal_5011 ), .Q ( signal_23902 ) ) ;
    buf_clk cell_9245 ( .C ( clk ), .D ( signal_1602 ), .Q ( signal_23938 ) ) ;
    buf_clk cell_9261 ( .C ( clk ), .D ( signal_5064 ), .Q ( signal_23954 ) ) ;
    buf_clk cell_9277 ( .C ( clk ), .D ( signal_5065 ), .Q ( signal_23970 ) ) ;
    buf_clk cell_9293 ( .C ( clk ), .D ( signal_5066 ), .Q ( signal_23986 ) ) ;
    buf_clk cell_9309 ( .C ( clk ), .D ( signal_5067 ), .Q ( signal_24002 ) ) ;
    buf_clk cell_9635 ( .C ( clk ), .D ( signal_1539 ), .Q ( signal_24328 ) ) ;
    buf_clk cell_9653 ( .C ( clk ), .D ( signal_4812 ), .Q ( signal_24346 ) ) ;
    buf_clk cell_9671 ( .C ( clk ), .D ( signal_4813 ), .Q ( signal_24364 ) ) ;
    buf_clk cell_9689 ( .C ( clk ), .D ( signal_4814 ), .Q ( signal_24382 ) ) ;
    buf_clk cell_9707 ( .C ( clk ), .D ( signal_4815 ), .Q ( signal_24400 ) ) ;
    buf_clk cell_9885 ( .C ( clk ), .D ( signal_1603 ), .Q ( signal_24578 ) ) ;
    buf_clk cell_9905 ( .C ( clk ), .D ( signal_5068 ), .Q ( signal_24598 ) ) ;
    buf_clk cell_9925 ( .C ( clk ), .D ( signal_5069 ), .Q ( signal_24618 ) ) ;
    buf_clk cell_9945 ( .C ( clk ), .D ( signal_5070 ), .Q ( signal_24638 ) ) ;
    buf_clk cell_9965 ( .C ( clk ), .D ( signal_5071 ), .Q ( signal_24658 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1644 ( .a ({signal_3827, signal_3826, signal_3825, signal_3824, signal_1292}), .b ({signal_17817, signal_17815, signal_17813, signal_17811, signal_17809}), .clk ( clk ), .r ({Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540]}), .c ({signal_5295, signal_5294, signal_5293, signal_5292, signal_1659}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1652 ( .a ({signal_17827, signal_17825, signal_17823, signal_17821, signal_17819}), .b ({signal_4199, signal_4198, signal_4197, signal_4196, signal_1385}), .clk ( clk ), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550]}), .c ({signal_5327, signal_5326, signal_5325, signal_5324, signal_1667}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1662 ( .a ({signal_17837, signal_17835, signal_17833, signal_17831, signal_17829}), .b ({signal_3975, signal_3974, signal_3973, signal_3972, signal_1329}), .clk ( clk ), .r ({Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({signal_5367, signal_5366, signal_5365, signal_5364, signal_1677}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1672 ( .a ({signal_17847, signal_17845, signal_17843, signal_17841, signal_17839}), .b ({signal_4031, signal_4030, signal_4029, signal_4028, signal_1343}), .clk ( clk ), .r ({Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570]}), .c ({signal_5407, signal_5406, signal_5405, signal_5404, signal_1687}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1683 ( .a ({signal_17857, signal_17855, signal_17853, signal_17851, signal_17849}), .b ({signal_4091, signal_4090, signal_4089, signal_4088, signal_1358}), .clk ( clk ), .r ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580]}), .c ({signal_5451, signal_5450, signal_5449, signal_5448, signal_1698}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1685 ( .a ({signal_17867, signal_17865, signal_17863, signal_17861, signal_17859}), .b ({signal_4099, signal_4098, signal_4097, signal_4096, signal_1360}), .clk ( clk ), .r ({Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .c ({signal_5459, signal_5458, signal_5457, signal_5456, signal_1700}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1686 ( .a ({signal_17877, signal_17875, signal_17873, signal_17871, signal_17869}), .b ({signal_4443, signal_4442, signal_4441, signal_4440, signal_1446}), .clk ( clk ), .r ({Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600]}), .c ({signal_5463, signal_5462, signal_5461, signal_5460, signal_1701}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1688 ( .a ({signal_17887, signal_17885, signal_17883, signal_17881, signal_17879}), .b ({signal_4443, signal_4442, signal_4441, signal_4440, signal_1446}), .clk ( clk ), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610]}), .c ({signal_5471, signal_5470, signal_5469, signal_5468, signal_1703}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1689 ( .a ({signal_17887, signal_17885, signal_17883, signal_17881, signal_17879}), .b ({signal_4499, signal_4498, signal_4497, signal_4496, signal_1460}), .clk ( clk ), .r ({Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({signal_5475, signal_5474, signal_5473, signal_5472, signal_1704}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1690 ( .a ({signal_17897, signal_17895, signal_17893, signal_17891, signal_17889}), .b ({signal_4503, signal_4502, signal_4501, signal_4500, signal_1461}), .clk ( clk ), .r ({Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630]}), .c ({signal_5479, signal_5478, signal_5477, signal_5476, signal_1705}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1691 ( .a ({signal_17907, signal_17905, signal_17903, signal_17901, signal_17899}), .b ({signal_4507, signal_4506, signal_4505, signal_4504, signal_1462}), .clk ( clk ), .r ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640]}), .c ({signal_5483, signal_5482, signal_5481, signal_5480, signal_1706}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1692 ( .a ({signal_17917, signal_17915, signal_17913, signal_17911, signal_17909}), .b ({signal_4459, signal_4458, signal_4457, signal_4456, signal_1450}), .clk ( clk ), .r ({Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .c ({signal_5487, signal_5486, signal_5485, signal_5484, signal_1707}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1694 ( .a ({signal_17947, signal_17941, signal_17935, signal_17929, signal_17923}), .b ({signal_4571, signal_4570, signal_4569, signal_4568, signal_1478}), .clk ( clk ), .r ({Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660]}), .c ({signal_5495, signal_5494, signal_5493, signal_5492, signal_1709}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1695 ( .a ({signal_17957, signal_17955, signal_17953, signal_17951, signal_17949}), .b ({signal_4111, signal_4110, signal_4109, signal_4108, signal_1363}), .clk ( clk ), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670]}), .c ({signal_5499, signal_5498, signal_5497, signal_5496, signal_1710}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1696 ( .a ({signal_17967, signal_17965, signal_17963, signal_17961, signal_17959}), .b ({signal_4399, signal_4398, signal_4397, signal_4396, signal_1435}), .clk ( clk ), .r ({Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({signal_5503, signal_5502, signal_5501, signal_5500, signal_1711}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1697 ( .a ({signal_17977, signal_17975, signal_17973, signal_17971, signal_17969}), .b ({signal_4555, signal_4554, signal_4553, signal_4552, signal_1474}), .clk ( clk ), .r ({Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690]}), .c ({signal_5507, signal_5506, signal_5505, signal_5504, signal_1712}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1699 ( .a ({signal_17987, signal_17985, signal_17983, signal_17981, signal_17979}), .b ({signal_4647, signal_4646, signal_4645, signal_4644, signal_1497}), .clk ( clk ), .r ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700]}), .c ({signal_5515, signal_5514, signal_5513, signal_5512, signal_1714}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1715 ( .a ({signal_5295, signal_5294, signal_5293, signal_5292, signal_1659}), .b ({signal_5579, signal_5578, signal_5577, signal_5576, signal_1730}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1721 ( .a ({signal_5327, signal_5326, signal_5325, signal_5324, signal_1667}), .b ({signal_5603, signal_5602, signal_5601, signal_5600, signal_1736}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1725 ( .a ({signal_5367, signal_5366, signal_5365, signal_5364, signal_1677}), .b ({signal_5619, signal_5618, signal_5617, signal_5616, signal_1740}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1737 ( .a ({signal_5459, signal_5458, signal_5457, signal_5456, signal_1700}), .b ({signal_5667, signal_5666, signal_5665, signal_5664, signal_1752}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1738 ( .a ({signal_5463, signal_5462, signal_5461, signal_5460, signal_1701}), .b ({signal_5671, signal_5670, signal_5669, signal_5668, signal_1753}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1740 ( .a ({signal_5471, signal_5470, signal_5469, signal_5468, signal_1703}), .b ({signal_5679, signal_5678, signal_5677, signal_5676, signal_1755}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1741 ( .a ({signal_5475, signal_5474, signal_5473, signal_5472, signal_1704}), .b ({signal_5683, signal_5682, signal_5681, signal_5680, signal_1756}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1742 ( .a ({signal_5479, signal_5478, signal_5477, signal_5476, signal_1705}), .b ({signal_5687, signal_5686, signal_5685, signal_5684, signal_1757}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1743 ( .a ({signal_5483, signal_5482, signal_5481, signal_5480, signal_1706}), .b ({signal_5691, signal_5690, signal_5689, signal_5688, signal_1758}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1744 ( .a ({signal_5487, signal_5486, signal_5485, signal_5484, signal_1707}), .b ({signal_5695, signal_5694, signal_5693, signal_5692, signal_1759}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1746 ( .a ({signal_5495, signal_5494, signal_5493, signal_5492, signal_1709}), .b ({signal_5703, signal_5702, signal_5701, signal_5700, signal_1761}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1747 ( .a ({signal_5503, signal_5502, signal_5501, signal_5500, signal_1711}), .b ({signal_5707, signal_5706, signal_5705, signal_5704, signal_1762}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1748 ( .a ({signal_5507, signal_5506, signal_5505, signal_5504, signal_1712}), .b ({signal_5711, signal_5710, signal_5709, signal_5708, signal_1763}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1750 ( .a ({signal_5515, signal_5514, signal_5513, signal_5512, signal_1714}), .b ({signal_5719, signal_5718, signal_5717, signal_5716, signal_1765}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1752 ( .a ({signal_4783, signal_4782, signal_4781, signal_4780, signal_1531}), .b ({signal_4787, signal_4786, signal_4785, signal_4784, signal_1532}), .clk ( clk ), .r ({Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .c ({signal_5727, signal_5726, signal_5725, signal_5724, signal_1767}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1759 ( .a ({signal_17997, signal_17995, signal_17993, signal_17991, signal_17989}), .b ({signal_4707, signal_4706, signal_4705, signal_4704, signal_1512}), .clk ( clk ), .r ({Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720]}), .c ({signal_5755, signal_5754, signal_5753, signal_5752, signal_1774}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1763 ( .a ({signal_18007, signal_18005, signal_18003, signal_18001, signal_17999}), .b ({signal_4727, signal_4726, signal_4725, signal_4724, signal_1517}), .clk ( clk ), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730]}), .c ({signal_5771, signal_5770, signal_5769, signal_5768, signal_1778}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1768 ( .a ({signal_4759, signal_4758, signal_4757, signal_4756, signal_1525}), .b ({signal_4763, signal_4762, signal_4761, signal_4760, signal_1526}), .clk ( clk ), .r ({Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({signal_5791, signal_5790, signal_5789, signal_5788, signal_1783}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1771 ( .a ({signal_4751, signal_4750, signal_4749, signal_4748, signal_1523}), .b ({signal_4779, signal_4778, signal_4777, signal_4776, signal_1530}), .clk ( clk ), .r ({Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750]}), .c ({signal_5803, signal_5802, signal_5801, signal_5800, signal_1786}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1774 ( .a ({signal_18017, signal_18015, signal_18013, signal_18011, signal_18009}), .b ({signal_4803, signal_4802, signal_4801, signal_4800, signal_1536}), .clk ( clk ), .r ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760]}), .c ({signal_5815, signal_5814, signal_5813, signal_5812, signal_1789}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1775 ( .a ({signal_4823, signal_4822, signal_4821, signal_4820, signal_1541}), .b ({signal_4827, signal_4826, signal_4825, signal_4824, signal_1542}), .clk ( clk ), .r ({Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .c ({signal_5819, signal_5818, signal_5817, signal_5816, signal_1790}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1777 ( .a ({signal_18027, signal_18025, signal_18023, signal_18021, signal_18019}), .b ({signal_4843, signal_4842, signal_4841, signal_4840, signal_1546}), .clk ( clk ), .r ({Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780]}), .c ({signal_5827, signal_5826, signal_5825, signal_5824, signal_1792}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1780 ( .a ({signal_18037, signal_18035, signal_18033, signal_18031, signal_18029}), .b ({signal_5255, signal_5254, signal_5253, signal_5252, signal_1649}), .clk ( clk ), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790]}), .c ({signal_5839, signal_5838, signal_5837, signal_5836, signal_1795}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1781 ( .a ({signal_5035, signal_5034, signal_5033, signal_5032, signal_1594}), .b ({signal_5103, signal_5102, signal_5101, signal_5100, signal_1611}), .clk ( clk ), .r ({Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({signal_5843, signal_5842, signal_5841, signal_5840, signal_1796}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1787 ( .a ({signal_18047, signal_18045, signal_18043, signal_18041, signal_18039}), .b ({signal_4903, signal_4902, signal_4901, signal_4900, signal_1561}), .clk ( clk ), .r ({Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810]}), .c ({signal_5867, signal_5866, signal_5865, signal_5864, signal_1802}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1788 ( .a ({signal_4911, signal_4910, signal_4909, signal_4908, signal_1563}), .b ({signal_18057, signal_18055, signal_18053, signal_18051, signal_18049}), .clk ( clk ), .r ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820]}), .c ({signal_5871, signal_5870, signal_5869, signal_5868, signal_1803}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1789 ( .a ({signal_18067, signal_18065, signal_18063, signal_18061, signal_18059}), .b ({signal_5271, signal_5270, signal_5269, signal_5268, signal_1653}), .clk ( clk ), .r ({Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .c ({signal_5875, signal_5874, signal_5873, signal_5872, signal_1804}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1790 ( .a ({signal_18077, signal_18075, signal_18073, signal_18071, signal_18069}), .b ({signal_5275, signal_5274, signal_5273, signal_5272, signal_1654}), .clk ( clk ), .r ({Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840]}), .c ({signal_5879, signal_5878, signal_5877, signal_5876, signal_1805}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1791 ( .a ({signal_18087, signal_18085, signal_18083, signal_18081, signal_18079}), .b ({signal_5279, signal_5278, signal_5277, signal_5276, signal_1655}), .clk ( clk ), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850]}), .c ({signal_5883, signal_5882, signal_5881, signal_5880, signal_1806}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1792 ( .a ({signal_4923, signal_4922, signal_4921, signal_4920, signal_1566}), .b ({signal_4927, signal_4926, signal_4925, signal_4924, signal_1567}), .clk ( clk ), .r ({Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({signal_5887, signal_5886, signal_5885, signal_5884, signal_1807}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1793 ( .a ({signal_3807, signal_3806, signal_3805, signal_3804, signal_1287}), .b ({signal_4931, signal_4930, signal_4929, signal_4928, signal_1568}), .clk ( clk ), .r ({Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870]}), .c ({signal_5891, signal_5890, signal_5889, signal_5888, signal_1808}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1794 ( .a ({signal_5219, signal_5218, signal_5217, signal_5216, signal_1640}), .b ({signal_4935, signal_4934, signal_4933, signal_4932, signal_1569}), .clk ( clk ), .r ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880]}), .c ({signal_5895, signal_5894, signal_5893, signal_5892, signal_1809}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1795 ( .a ({signal_17897, signal_17895, signal_17893, signal_17891, signal_17889}), .b ({signal_4943, signal_4942, signal_4941, signal_4940, signal_1571}), .clk ( clk ), .r ({Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .c ({signal_5899, signal_5898, signal_5897, signal_5896, signal_1810}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1796 ( .a ({signal_4711, signal_4710, signal_4709, signal_4708, signal_1513}), .b ({signal_4947, signal_4946, signal_4945, signal_4944, signal_1572}), .clk ( clk ), .r ({Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900]}), .c ({signal_5903, signal_5902, signal_5901, signal_5900, signal_1811}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1797 ( .a ({signal_18097, signal_18095, signal_18093, signal_18091, signal_18089}), .b ({signal_4951, signal_4950, signal_4949, signal_4948, signal_1573}), .clk ( clk ), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910]}), .c ({signal_5907, signal_5906, signal_5905, signal_5904, signal_1812}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1798 ( .a ({signal_18107, signal_18105, signal_18103, signal_18101, signal_18099}), .b ({signal_5299, signal_5298, signal_5297, signal_5296, signal_1660}), .clk ( clk ), .r ({Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({signal_5911, signal_5910, signal_5909, signal_5908, signal_1813}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1799 ( .a ({signal_18117, signal_18115, signal_18113, signal_18111, signal_18109}), .b ({signal_4955, signal_4954, signal_4953, signal_4952, signal_1574}), .clk ( clk ), .r ({Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930]}), .c ({signal_5915, signal_5914, signal_5913, signal_5912, signal_1814}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1800 ( .a ({signal_18127, signal_18125, signal_18123, signal_18121, signal_18119}), .b ({signal_4967, signal_4966, signal_4965, signal_4964, signal_1577}), .clk ( clk ), .r ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940]}), .c ({signal_5919, signal_5918, signal_5917, signal_5916, signal_1815}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1801 ( .a ({signal_18137, signal_18135, signal_18133, signal_18131, signal_18129}), .b ({signal_5303, signal_5302, signal_5301, signal_5300, signal_1661}), .clk ( clk ), .r ({Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .c ({signal_5923, signal_5922, signal_5921, signal_5920, signal_1816}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1802 ( .a ({signal_18147, signal_18145, signal_18143, signal_18141, signal_18139}), .b ({signal_4923, signal_4922, signal_4921, signal_4920, signal_1566}), .clk ( clk ), .r ({Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960]}), .c ({signal_5927, signal_5926, signal_5925, signal_5924, signal_1817}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1803 ( .a ({signal_4975, signal_4974, signal_4973, signal_4972, signal_1579}), .b ({signal_4979, signal_4978, signal_4977, signal_4976, signal_1580}), .clk ( clk ), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970]}), .c ({signal_5931, signal_5930, signal_5929, signal_5928, signal_1818}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1804 ( .a ({signal_4755, signal_4754, signal_4753, signal_4752, signal_1524}), .b ({signal_4999, signal_4998, signal_4997, signal_4996, signal_1585}), .clk ( clk ), .r ({Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({signal_5935, signal_5934, signal_5933, signal_5932, signal_1819}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1805 ( .a ({signal_4955, signal_4954, signal_4953, signal_4952, signal_1574}), .b ({signal_5003, signal_5002, signal_5001, signal_5000, signal_1586}), .clk ( clk ), .r ({Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990]}), .c ({signal_5939, signal_5938, signal_5937, signal_5936, signal_1820}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1806 ( .a ({signal_18167, signal_18163, signal_18159, signal_18155, signal_18151}), .b ({signal_5331, signal_5330, signal_5329, signal_5328, signal_1668}), .clk ( clk ), .r ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000]}), .c ({signal_5943, signal_5942, signal_5941, signal_5940, signal_1821}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1807 ( .a ({signal_18177, signal_18175, signal_18173, signal_18171, signal_18169}), .b ({signal_5323, signal_5322, signal_5321, signal_5320, signal_1666}), .clk ( clk ), .r ({Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .c ({signal_5947, signal_5946, signal_5945, signal_5944, signal_1822}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1808 ( .a ({signal_18187, signal_18185, signal_18183, signal_18181, signal_18179}), .b ({signal_5339, signal_5338, signal_5337, signal_5336, signal_1670}), .clk ( clk ), .r ({Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020]}), .c ({signal_5951, signal_5950, signal_5949, signal_5948, signal_1823}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1809 ( .a ({signal_18207, signal_18203, signal_18199, signal_18195, signal_18191}), .b ({signal_5343, signal_5342, signal_5341, signal_5340, signal_1671}), .clk ( clk ), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030]}), .c ({signal_5955, signal_5954, signal_5953, signal_5952, signal_1824}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1810 ( .a ({signal_5175, signal_5174, signal_5173, signal_5172, signal_1629}), .b ({signal_5179, signal_5178, signal_5177, signal_5176, signal_1630}), .clk ( clk ), .r ({Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({signal_5959, signal_5958, signal_5957, signal_5956, signal_1825}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1811 ( .a ({signal_4775, signal_4774, signal_4773, signal_4772, signal_1529}), .b ({signal_5347, signal_5346, signal_5345, signal_5344, signal_1672}), .clk ( clk ), .r ({Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050]}), .c ({signal_5963, signal_5962, signal_5961, signal_5960, signal_1826}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1812 ( .a ({signal_4811, signal_4810, signal_4809, signal_4808, signal_1538}), .b ({signal_5055, signal_5054, signal_5053, signal_5052, signal_1599}), .clk ( clk ), .r ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060]}), .c ({signal_5967, signal_5966, signal_5965, signal_5964, signal_1827}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1813 ( .a ({signal_4835, signal_4834, signal_4833, signal_4832, signal_1544}), .b ({signal_5079, signal_5078, signal_5077, signal_5076, signal_1605}), .clk ( clk ), .r ({Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .c ({signal_5971, signal_5970, signal_5969, signal_5968, signal_1828}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1814 ( .a ({signal_4839, signal_4838, signal_4837, signal_4836, signal_1545}), .b ({signal_5087, signal_5086, signal_5085, signal_5084, signal_1607}), .clk ( clk ), .r ({Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080]}), .c ({signal_5975, signal_5974, signal_5973, signal_5972, signal_1829}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1815 ( .a ({signal_18217, signal_18215, signal_18213, signal_18211, signal_18209}), .b ({signal_5091, signal_5090, signal_5089, signal_5088, signal_1608}), .clk ( clk ), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090]}), .c ({signal_5979, signal_5978, signal_5977, signal_5976, signal_1830}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1816 ( .a ({signal_18227, signal_18225, signal_18223, signal_18221, signal_18219}), .b ({signal_5395, signal_5394, signal_5393, signal_5392, signal_1684}), .clk ( clk ), .r ({Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({signal_5983, signal_5982, signal_5981, signal_5980, signal_1831}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1817 ( .a ({signal_18237, signal_18235, signal_18233, signal_18231, signal_18229}), .b ({signal_5399, signal_5398, signal_5397, signal_5396, signal_1685}), .clk ( clk ), .r ({Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110]}), .c ({signal_5987, signal_5986, signal_5985, signal_5984, signal_1832}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1818 ( .a ({signal_4943, signal_4942, signal_4941, signal_4940, signal_1571}), .b ({signal_5043, signal_5042, signal_5041, signal_5040, signal_1596}), .clk ( clk ), .r ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120]}), .c ({signal_5991, signal_5990, signal_5989, signal_5988, signal_1833}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1820 ( .a ({signal_4035, signal_4034, signal_4033, signal_4032, signal_1344}), .b ({signal_5099, signal_5098, signal_5097, signal_5096, signal_1610}), .clk ( clk ), .r ({Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .c ({signal_5999, signal_5998, signal_5997, signal_5996, signal_1835}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1821 ( .a ({signal_18247, signal_18245, signal_18243, signal_18241, signal_18239}), .b ({signal_5107, signal_5106, signal_5105, signal_5104, signal_1612}), .clk ( clk ), .r ({Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140]}), .c ({signal_6003, signal_6002, signal_6001, signal_6000, signal_1836}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1822 ( .a ({signal_18257, signal_18255, signal_18253, signal_18251, signal_18249}), .b ({signal_5119, signal_5118, signal_5117, signal_5116, signal_1615}), .clk ( clk ), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150]}), .c ({signal_6007, signal_6006, signal_6005, signal_6004, signal_1837}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1823 ( .a ({signal_4883, signal_4882, signal_4881, signal_4880, signal_1556}), .b ({signal_5127, signal_5126, signal_5125, signal_5124, signal_1617}), .clk ( clk ), .r ({Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({signal_6011, signal_6010, signal_6009, signal_6008, signal_1838}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1824 ( .a ({signal_18267, signal_18265, signal_18263, signal_18261, signal_18259}), .b ({signal_5427, signal_5426, signal_5425, signal_5424, signal_1692}), .clk ( clk ), .r ({Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170]}), .c ({signal_6015, signal_6014, signal_6013, signal_6012, signal_1839}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1825 ( .a ({signal_18277, signal_18275, signal_18273, signal_18271, signal_18269}), .b ({signal_5139, signal_5138, signal_5137, signal_5136, signal_1620}), .clk ( clk ), .r ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180]}), .c ({signal_6019, signal_6018, signal_6017, signal_6016, signal_1840}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1826 ( .a ({signal_18287, signal_18285, signal_18283, signal_18281, signal_18279}), .b ({signal_5119, signal_5118, signal_5117, signal_5116, signal_1615}), .clk ( clk ), .r ({Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .c ({signal_6023, signal_6022, signal_6021, signal_6020, signal_1841}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1827 ( .a ({signal_18297, signal_18295, signal_18293, signal_18291, signal_18289}), .b ({signal_5439, signal_5438, signal_5437, signal_5436, signal_1695}), .clk ( clk ), .r ({Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200]}), .c ({signal_6027, signal_6026, signal_6025, signal_6024, signal_1842}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1828 ( .a ({signal_4915, signal_4914, signal_4913, signal_4912, signal_1564}), .b ({signal_5151, signal_5150, signal_5149, signal_5148, signal_1623}), .clk ( clk ), .r ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210]}), .c ({signal_6031, signal_6030, signal_6029, signal_6028, signal_1843}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1829 ( .a ({signal_18307, signal_18305, signal_18303, signal_18301, signal_18299}), .b ({signal_5155, signal_5154, signal_5153, signal_5152, signal_1624}), .clk ( clk ), .r ({Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .c ({signal_6035, signal_6034, signal_6033, signal_6032, signal_1844}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1830 ( .a ({signal_5163, signal_5162, signal_5161, signal_5160, signal_1626}), .b ({signal_5167, signal_5166, signal_5165, signal_5164, signal_1627}), .clk ( clk ), .r ({Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230]}), .c ({signal_6039, signal_6038, signal_6037, signal_6036, signal_1845}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1831 ( .a ({signal_5027, signal_5026, signal_5025, signal_5024, signal_1592}), .b ({signal_5171, signal_5170, signal_5169, signal_5168, signal_1628}), .clk ( clk ), .r ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240]}), .c ({signal_6043, signal_6042, signal_6041, signal_6040, signal_1846}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1832 ( .a ({signal_4751, signal_4750, signal_4749, signal_4748, signal_1523}), .b ({signal_5195, signal_5194, signal_5193, signal_5192, signal_1634}), .clk ( clk ), .r ({Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .c ({signal_6047, signal_6046, signal_6045, signal_6044, signal_1847}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1833 ( .a ({signal_4107, signal_4106, signal_4105, signal_4104, signal_1362}), .b ({signal_5199, signal_5198, signal_5197, signal_5196, signal_1635}), .clk ( clk ), .r ({Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260]}), .c ({signal_6051, signal_6050, signal_6049, signal_6048, signal_1848}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1842 ( .a ({signal_5771, signal_5770, signal_5769, signal_5768, signal_1778}), .b ({signal_6087, signal_6086, signal_6085, signal_6084, signal_1857}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1853 ( .a ({signal_5839, signal_5838, signal_5837, signal_5836, signal_1795}), .b ({signal_6131, signal_6130, signal_6129, signal_6128, signal_1868}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1859 ( .a ({signal_5879, signal_5878, signal_5877, signal_5876, signal_1805}), .b ({signal_6155, signal_6154, signal_6153, signal_6152, signal_1874}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1860 ( .a ({signal_5887, signal_5886, signal_5885, signal_5884, signal_1807}), .b ({signal_6159, signal_6158, signal_6157, signal_6156, signal_1875}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1861 ( .a ({signal_5907, signal_5906, signal_5905, signal_5904, signal_1812}), .b ({signal_6163, signal_6162, signal_6161, signal_6160, signal_1876}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1862 ( .a ({signal_5923, signal_5922, signal_5921, signal_5920, signal_1816}), .b ({signal_6167, signal_6166, signal_6165, signal_6164, signal_1877}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1863 ( .a ({signal_5927, signal_5926, signal_5925, signal_5924, signal_1817}), .b ({signal_6171, signal_6170, signal_6169, signal_6168, signal_1878}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1864 ( .a ({signal_5943, signal_5942, signal_5941, signal_5940, signal_1821}), .b ({signal_6175, signal_6174, signal_6173, signal_6172, signal_1879}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1865 ( .a ({signal_5947, signal_5946, signal_5945, signal_5944, signal_1822}), .b ({signal_6179, signal_6178, signal_6177, signal_6176, signal_1880}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1866 ( .a ({signal_5951, signal_5950, signal_5949, signal_5948, signal_1823}), .b ({signal_6183, signal_6182, signal_6181, signal_6180, signal_1881}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1867 ( .a ({signal_5955, signal_5954, signal_5953, signal_5952, signal_1824}), .b ({signal_6187, signal_6186, signal_6185, signal_6184, signal_1882}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1868 ( .a ({signal_5971, signal_5970, signal_5969, signal_5968, signal_1828}), .b ({signal_6191, signal_6190, signal_6189, signal_6188, signal_1883}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1869 ( .a ({signal_5975, signal_5974, signal_5973, signal_5972, signal_1829}), .b ({signal_6195, signal_6194, signal_6193, signal_6192, signal_1884}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1870 ( .a ({signal_5983, signal_5982, signal_5981, signal_5980, signal_1831}), .b ({signal_6199, signal_6198, signal_6197, signal_6196, signal_1885}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1871 ( .a ({signal_5987, signal_5986, signal_5985, signal_5984, signal_1832}), .b ({signal_6203, signal_6202, signal_6201, signal_6200, signal_1886}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1873 ( .a ({signal_6027, signal_6026, signal_6025, signal_6024, signal_1842}), .b ({signal_6211, signal_6210, signal_6209, signal_6208, signal_1888}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1874 ( .a ({signal_6035, signal_6034, signal_6033, signal_6032, signal_1844}), .b ({signal_6215, signal_6214, signal_6213, signal_6212, signal_1889}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1876 ( .a ({signal_5519, signal_5518, signal_5517, signal_5516, signal_1715}), .b ({signal_18317, signal_18315, signal_18313, signal_18311, signal_18309}), .clk ( clk ), .r ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270]}), .c ({signal_6223, signal_6222, signal_6221, signal_6220, signal_1891}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1877 ( .a ({signal_18337, signal_18333, signal_18329, signal_18325, signal_18321}), .b ({signal_5523, signal_5522, signal_5521, signal_5520, signal_1716}), .clk ( clk ), .r ({Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .c ({signal_6227, signal_6226, signal_6225, signal_6224, signal_1892}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1878 ( .a ({signal_18347, signal_18345, signal_18343, signal_18341, signal_18339}), .b ({signal_5527, signal_5526, signal_5525, signal_5524, signal_1717}), .clk ( clk ), .r ({Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290]}), .c ({signal_6231, signal_6230, signal_6229, signal_6228, signal_1893}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1879 ( .a ({signal_17887, signal_17885, signal_17883, signal_17881, signal_17879}), .b ({signal_5531, signal_5530, signal_5529, signal_5528, signal_1718}), .clk ( clk ), .r ({Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300]}), .c ({signal_6235, signal_6234, signal_6233, signal_6232, signal_1894}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1880 ( .a ({signal_17987, signal_17985, signal_17983, signal_17981, signal_17979}), .b ({signal_5731, signal_5730, signal_5729, signal_5728, signal_1768}), .clk ( clk ), .r ({Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310]}), .c ({signal_6239, signal_6238, signal_6237, signal_6236, signal_1895}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1881 ( .a ({signal_18367, signal_18363, signal_18359, signal_18355, signal_18351}), .b ({signal_5535, signal_5534, signal_5533, signal_5532, signal_1719}), .clk ( clk ), .r ({Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320]}), .c ({signal_6243, signal_6242, signal_6241, signal_6240, signal_1896}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1882 ( .a ({signal_5539, signal_5538, signal_5537, signal_5536, signal_1720}), .b ({signal_18377, signal_18375, signal_18373, signal_18371, signal_18369}), .clk ( clk ), .r ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330]}), .c ({signal_6247, signal_6246, signal_6245, signal_6244, signal_1897}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1883 ( .a ({signal_18387, signal_18385, signal_18383, signal_18381, signal_18379}), .b ({signal_5543, signal_5542, signal_5541, signal_5540, signal_1721}), .clk ( clk ), .r ({Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .c ({signal_6251, signal_6250, signal_6249, signal_6248, signal_1898}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1884 ( .a ({signal_18397, signal_18395, signal_18393, signal_18391, signal_18389}), .b ({signal_5547, signal_5546, signal_5545, signal_5544, signal_1722}), .clk ( clk ), .r ({Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350]}), .c ({signal_6255, signal_6254, signal_6253, signal_6252, signal_1899}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1885 ( .a ({signal_18427, signal_18421, signal_18415, signal_18409, signal_18403}), .b ({signal_5551, signal_5550, signal_5549, signal_5548, signal_1723}), .clk ( clk ), .r ({Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360]}), .c ({signal_6259, signal_6258, signal_6257, signal_6256, signal_1900}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1886 ( .a ({signal_17917, signal_17915, signal_17913, signal_17911, signal_17909}), .b ({signal_5735, signal_5734, signal_5733, signal_5732, signal_1769}), .clk ( clk ), .r ({Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370]}), .c ({signal_6263, signal_6262, signal_6261, signal_6260, signal_1901}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1887 ( .a ({signal_18437, signal_18435, signal_18433, signal_18431, signal_18429}), .b ({signal_5555, signal_5554, signal_5553, signal_5552, signal_1724}), .clk ( clk ), .r ({Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380]}), .c ({signal_6267, signal_6266, signal_6265, signal_6264, signal_1902}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1888 ( .a ({signal_18447, signal_18445, signal_18443, signal_18441, signal_18439}), .b ({signal_5563, signal_5562, signal_5561, signal_5560, signal_1726}), .clk ( clk ), .r ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390]}), .c ({signal_6271, signal_6270, signal_6269, signal_6268, signal_1903}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1889 ( .a ({signal_18457, signal_18455, signal_18453, signal_18451, signal_18449}), .b ({signal_5743, signal_5742, signal_5741, signal_5740, signal_1771}), .clk ( clk ), .r ({Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .c ({signal_6275, signal_6274, signal_6273, signal_6272, signal_1904}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1890 ( .a ({signal_17887, signal_17885, signal_17883, signal_17881, signal_17879}), .b ({signal_5567, signal_5566, signal_5565, signal_5564, signal_1727}), .clk ( clk ), .r ({Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410]}), .c ({signal_6279, signal_6278, signal_6277, signal_6276, signal_1905}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1891 ( .a ({signal_17987, signal_17985, signal_17983, signal_17981, signal_17979}), .b ({signal_5571, signal_5570, signal_5569, signal_5568, signal_1728}), .clk ( clk ), .r ({Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420]}), .c ({signal_6283, signal_6282, signal_6281, signal_6280, signal_1906}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1892 ( .a ({signal_18467, signal_18465, signal_18463, signal_18461, signal_18459}), .b ({signal_5575, signal_5574, signal_5573, signal_5572, signal_1729}), .clk ( clk ), .r ({Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430]}), .c ({signal_6287, signal_6286, signal_6285, signal_6284, signal_1907}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1894 ( .a ({signal_18007, signal_18005, signal_18003, signal_18001, signal_17999}), .b ({signal_5583, signal_5582, signal_5581, signal_5580, signal_1731}), .clk ( clk ), .r ({Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440]}), .c ({signal_6295, signal_6294, signal_6293, signal_6292, signal_1909}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1895 ( .a ({signal_18487, signal_18483, signal_18479, signal_18475, signal_18471}), .b ({signal_5587, signal_5586, signal_5585, signal_5584, signal_1732}), .clk ( clk ), .r ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450]}), .c ({signal_6299, signal_6298, signal_6297, signal_6296, signal_1910}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1896 ( .a ({signal_18497, signal_18495, signal_18493, signal_18491, signal_18489}), .b ({signal_5591, signal_5590, signal_5589, signal_5588, signal_1733}), .clk ( clk ), .r ({Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .c ({signal_6303, signal_6302, signal_6301, signal_6300, signal_1911}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1897 ( .a ({signal_18507, signal_18505, signal_18503, signal_18501, signal_18499}), .b ({signal_5595, signal_5594, signal_5593, signal_5592, signal_1734}), .clk ( clk ), .r ({Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470]}), .c ({signal_6307, signal_6306, signal_6305, signal_6304, signal_1912}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1898 ( .a ({signal_18517, signal_18515, signal_18513, signal_18511, signal_18509}), .b ({signal_5787, signal_5786, signal_5785, signal_5784, signal_1782}), .clk ( clk ), .r ({Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480]}), .c ({signal_6311, signal_6310, signal_6309, signal_6308, signal_1913}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1899 ( .a ({signal_18527, signal_18525, signal_18523, signal_18521, signal_18519}), .b ({signal_5599, signal_5598, signal_5597, signal_5596, signal_1735}), .clk ( clk ), .r ({Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490]}), .c ({signal_6315, signal_6314, signal_6313, signal_6312, signal_1914}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1900 ( .a ({signal_18447, signal_18445, signal_18443, signal_18441, signal_18439}), .b ({signal_5607, signal_5606, signal_5605, signal_5604, signal_1737}), .clk ( clk ), .r ({Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500]}), .c ({signal_6319, signal_6318, signal_6317, signal_6316, signal_1915}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1901 ( .a ({signal_5611, signal_5610, signal_5609, signal_5608, signal_1738}), .b ({signal_5355, signal_5354, signal_5353, signal_5352, signal_1674}), .clk ( clk ), .r ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510]}), .c ({signal_6323, signal_6322, signal_6321, signal_6320, signal_1916}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1903 ( .a ({signal_17897, signal_17895, signal_17893, signal_17891, signal_17889}), .b ({signal_5615, signal_5614, signal_5613, signal_5612, signal_1739}), .clk ( clk ), .r ({Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .c ({signal_6331, signal_6330, signal_6329, signal_6328, signal_1918}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1905 ( .a ({signal_18497, signal_18495, signal_18493, signal_18491, signal_18489}), .b ({signal_5623, signal_5622, signal_5621, signal_5620, signal_1741}), .clk ( clk ), .r ({Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530]}), .c ({signal_6339, signal_6338, signal_6337, signal_6336, signal_1920}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1906 ( .a ({signal_17977, signal_17975, signal_17973, signal_17971, signal_17969}), .b ({signal_5627, signal_5626, signal_5625, signal_5624, signal_1742}), .clk ( clk ), .r ({Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540]}), .c ({signal_6343, signal_6342, signal_6341, signal_6340, signal_1921}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1907 ( .a ({signal_18227, signal_18225, signal_18223, signal_18221, signal_18219}), .b ({signal_5631, signal_5630, signal_5629, signal_5628, signal_1743}), .clk ( clk ), .r ({Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550]}), .c ({signal_6347, signal_6346, signal_6345, signal_6344, signal_1922}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1908 ( .a ({signal_18367, signal_18363, signal_18359, signal_18355, signal_18351}), .b ({signal_5635, signal_5634, signal_5633, signal_5632, signal_1744}), .clk ( clk ), .r ({Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560]}), .c ({signal_6351, signal_6350, signal_6349, signal_6348, signal_1923}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1909 ( .a ({signal_18537, signal_18535, signal_18533, signal_18531, signal_18529}), .b ({signal_5787, signal_5786, signal_5785, signal_5784, signal_1782}), .clk ( clk ), .r ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570]}), .c ({signal_6355, signal_6354, signal_6353, signal_6352, signal_1924}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1910 ( .a ({signal_18547, signal_18545, signal_18543, signal_18541, signal_18539}), .b ({signal_5639, signal_5638, signal_5637, signal_5636, signal_1745}), .clk ( clk ), .r ({Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .c ({signal_6359, signal_6358, signal_6357, signal_6356, signal_1925}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1913 ( .a ({signal_18557, signal_18555, signal_18553, signal_18551, signal_18549}), .b ({signal_5643, signal_5642, signal_5641, signal_5640, signal_1746}), .clk ( clk ), .r ({Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590]}), .c ({signal_6371, signal_6370, signal_6369, signal_6368, signal_1928}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1914 ( .a ({signal_17977, signal_17975, signal_17973, signal_17971, signal_17969}), .b ({signal_5647, signal_5646, signal_5645, signal_5644, signal_1747}), .clk ( clk ), .r ({Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600]}), .c ({signal_6375, signal_6374, signal_6373, signal_6372, signal_1929}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1915 ( .a ({signal_17887, signal_17885, signal_17883, signal_17881, signal_17879}), .b ({signal_5651, signal_5650, signal_5649, signal_5648, signal_1748}), .clk ( clk ), .r ({Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610]}), .c ({signal_6379, signal_6378, signal_6377, signal_6376, signal_1930}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1916 ( .a ({signal_18567, signal_18565, signal_18563, signal_18561, signal_18559}), .b ({signal_5559, signal_5558, signal_5557, signal_5556, signal_1725}), .clk ( clk ), .r ({Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620]}), .c ({signal_6383, signal_6382, signal_6381, signal_6380, signal_1931}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1917 ( .a ({signal_18577, signal_18575, signal_18573, signal_18571, signal_18569}), .b ({signal_5575, signal_5574, signal_5573, signal_5572, signal_1729}), .clk ( clk ), .r ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630]}), .c ({signal_6387, signal_6386, signal_6385, signal_6384, signal_1932}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1919 ( .a ({signal_18597, signal_18593, signal_18589, signal_18585, signal_18581}), .b ({signal_5655, signal_5654, signal_5653, signal_5652, signal_1749}), .clk ( clk ), .r ({Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .c ({signal_6395, signal_6394, signal_6393, signal_6392, signal_1934}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1920 ( .a ({signal_18227, signal_18225, signal_18223, signal_18221, signal_18219}), .b ({signal_5659, signal_5658, signal_5657, signal_5656, signal_1750}), .clk ( clk ), .r ({Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650]}), .c ({signal_6399, signal_6398, signal_6397, signal_6396, signal_1935}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1923 ( .a ({signal_18607, signal_18605, signal_18603, signal_18601, signal_18599}), .b ({signal_5663, signal_5662, signal_5661, signal_5660, signal_1751}), .clk ( clk ), .r ({Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660]}), .c ({signal_6411, signal_6410, signal_6409, signal_6408, signal_1938}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1927 ( .a ({signal_18617, signal_18615, signal_18613, signal_18611, signal_18609}), .b ({signal_5675, signal_5674, signal_5673, signal_5672, signal_1754}), .clk ( clk ), .r ({Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670]}), .c ({signal_6427, signal_6426, signal_6425, signal_6424, signal_1942}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1932 ( .a ({signal_17877, signal_17875, signal_17873, signal_17871, signal_17869}), .b ({signal_5699, signal_5698, signal_5697, signal_5696, signal_1760}), .clk ( clk ), .r ({Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680]}), .c ({signal_6447, signal_6446, signal_6445, signal_6444, signal_1947}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1944 ( .a ({signal_18627, signal_18625, signal_18623, signal_18621, signal_18619}), .b ({signal_5715, signal_5714, signal_5713, signal_5712, signal_1764}), .clk ( clk ), .r ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690]}), .c ({signal_6495, signal_6494, signal_6493, signal_6492, signal_1959}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1948 ( .a ({signal_6227, signal_6226, signal_6225, signal_6224, signal_1892}), .b ({signal_6511, signal_6510, signal_6509, signal_6508, signal_1963}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1949 ( .a ({signal_6231, signal_6230, signal_6229, signal_6228, signal_1893}), .b ({signal_6515, signal_6514, signal_6513, signal_6512, signal_1964}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1950 ( .a ({signal_6239, signal_6238, signal_6237, signal_6236, signal_1895}), .b ({signal_6519, signal_6518, signal_6517, signal_6516, signal_1965}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1951 ( .a ({signal_6247, signal_6246, signal_6245, signal_6244, signal_1897}), .b ({signal_6523, signal_6522, signal_6521, signal_6520, signal_1966}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1952 ( .a ({signal_6251, signal_6250, signal_6249, signal_6248, signal_1898}), .b ({signal_6527, signal_6526, signal_6525, signal_6524, signal_1967}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1953 ( .a ({signal_6259, signal_6258, signal_6257, signal_6256, signal_1900}), .b ({signal_6531, signal_6530, signal_6529, signal_6528, signal_1968}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1954 ( .a ({signal_6263, signal_6262, signal_6261, signal_6260, signal_1901}), .b ({signal_6535, signal_6534, signal_6533, signal_6532, signal_1969}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1955 ( .a ({signal_6267, signal_6266, signal_6265, signal_6264, signal_1902}), .b ({signal_6539, signal_6538, signal_6537, signal_6536, signal_1970}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1956 ( .a ({signal_6271, signal_6270, signal_6269, signal_6268, signal_1903}), .b ({signal_6543, signal_6542, signal_6541, signal_6540, signal_1971}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1957 ( .a ({signal_6275, signal_6274, signal_6273, signal_6272, signal_1904}), .b ({signal_6547, signal_6546, signal_6545, signal_6544, signal_1972}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1958 ( .a ({signal_6279, signal_6278, signal_6277, signal_6276, signal_1905}), .b ({signal_6551, signal_6550, signal_6549, signal_6548, signal_1973}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1959 ( .a ({signal_6283, signal_6282, signal_6281, signal_6280, signal_1906}), .b ({signal_6555, signal_6554, signal_6553, signal_6552, signal_1974}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1960 ( .a ({signal_6287, signal_6286, signal_6285, signal_6284, signal_1907}), .b ({signal_6559, signal_6558, signal_6557, signal_6556, signal_1975}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1962 ( .a ({signal_6295, signal_6294, signal_6293, signal_6292, signal_1909}), .b ({signal_6567, signal_6566, signal_6565, signal_6564, signal_1977}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1963 ( .a ({signal_6299, signal_6298, signal_6297, signal_6296, signal_1910}), .b ({signal_6571, signal_6570, signal_6569, signal_6568, signal_1978}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1964 ( .a ({signal_6303, signal_6302, signal_6301, signal_6300, signal_1911}), .b ({signal_6575, signal_6574, signal_6573, signal_6572, signal_1979}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1965 ( .a ({signal_6307, signal_6306, signal_6305, signal_6304, signal_1912}), .b ({signal_6579, signal_6578, signal_6577, signal_6576, signal_1980}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1966 ( .a ({signal_6311, signal_6310, signal_6309, signal_6308, signal_1913}), .b ({signal_6583, signal_6582, signal_6581, signal_6580, signal_1981}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1967 ( .a ({signal_6315, signal_6314, signal_6313, signal_6312, signal_1914}), .b ({signal_6587, signal_6586, signal_6585, signal_6584, signal_1982}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1968 ( .a ({signal_6319, signal_6318, signal_6317, signal_6316, signal_1915}), .b ({signal_6591, signal_6590, signal_6589, signal_6588, signal_1983}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1970 ( .a ({signal_6331, signal_6330, signal_6329, signal_6328, signal_1918}), .b ({signal_6599, signal_6598, signal_6597, signal_6596, signal_1985}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1972 ( .a ({signal_6339, signal_6338, signal_6337, signal_6336, signal_1920}), .b ({signal_6607, signal_6606, signal_6605, signal_6604, signal_1987}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1973 ( .a ({signal_6343, signal_6342, signal_6341, signal_6340, signal_1921}), .b ({signal_6611, signal_6610, signal_6609, signal_6608, signal_1988}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1974 ( .a ({signal_6347, signal_6346, signal_6345, signal_6344, signal_1922}), .b ({signal_6615, signal_6614, signal_6613, signal_6612, signal_1989}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1975 ( .a ({signal_6351, signal_6350, signal_6349, signal_6348, signal_1923}), .b ({signal_6619, signal_6618, signal_6617, signal_6616, signal_1990}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1976 ( .a ({signal_6355, signal_6354, signal_6353, signal_6352, signal_1924}), .b ({signal_6623, signal_6622, signal_6621, signal_6620, signal_1991}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1977 ( .a ({signal_6359, signal_6358, signal_6357, signal_6356, signal_1925}), .b ({signal_6627, signal_6626, signal_6625, signal_6624, signal_1992}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1979 ( .a ({signal_6371, signal_6370, signal_6369, signal_6368, signal_1928}), .b ({signal_6635, signal_6634, signal_6633, signal_6632, signal_1994}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1980 ( .a ({signal_6375, signal_6374, signal_6373, signal_6372, signal_1929}), .b ({signal_6639, signal_6638, signal_6637, signal_6636, signal_1995}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1981 ( .a ({signal_6379, signal_6378, signal_6377, signal_6376, signal_1930}), .b ({signal_6643, signal_6642, signal_6641, signal_6640, signal_1996}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1982 ( .a ({signal_6383, signal_6382, signal_6381, signal_6380, signal_1931}), .b ({signal_6647, signal_6646, signal_6645, signal_6644, signal_1997}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1983 ( .a ({signal_6387, signal_6386, signal_6385, signal_6384, signal_1932}), .b ({signal_6651, signal_6650, signal_6649, signal_6648, signal_1998}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1984 ( .a ({signal_6395, signal_6394, signal_6393, signal_6392, signal_1934}), .b ({signal_6655, signal_6654, signal_6653, signal_6652, signal_1999}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1985 ( .a ({signal_6399, signal_6398, signal_6397, signal_6396, signal_1935}), .b ({signal_6659, signal_6658, signal_6657, signal_6656, signal_2000}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1988 ( .a ({signal_6411, signal_6410, signal_6409, signal_6408, signal_1938}), .b ({signal_6671, signal_6670, signal_6669, signal_6668, signal_2003}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1990 ( .a ({signal_6427, signal_6426, signal_6425, signal_6424, signal_1942}), .b ({signal_6679, signal_6678, signal_6677, signal_6676, signal_2005}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1991 ( .a ({signal_6447, signal_6446, signal_6445, signal_6444, signal_1947}), .b ({signal_6683, signal_6682, signal_6681, signal_6680, signal_2006}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1996 ( .a ({signal_6495, signal_6494, signal_6493, signal_6492, signal_1959}), .b ({signal_6703, signal_6702, signal_6701, signal_6700, signal_2011}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2000 ( .a ({signal_6111, signal_6110, signal_6109, signal_6108, signal_1863}), .b ({signal_5035, signal_5034, signal_5033, signal_5032, signal_1594}), .clk ( clk ), .r ({Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .c ({signal_6719, signal_6718, signal_6717, signal_6716, signal_2015}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2001 ( .a ({signal_6067, signal_6066, signal_6065, signal_6064, signal_1852}), .b ({signal_4919, signal_4918, signal_4917, signal_4916, signal_1565}), .clk ( clk ), .r ({Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710]}), .c ({signal_6723, signal_6722, signal_6721, signal_6720, signal_2016}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2003 ( .a ({signal_6079, signal_6078, signal_6077, signal_6076, signal_1855}), .b ({signal_6083, signal_6082, signal_6081, signal_6080, signal_1856}), .clk ( clk ), .r ({Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720]}), .c ({signal_6731, signal_6730, signal_6729, signal_6728, signal_2018}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2004 ( .a ({signal_18637, signal_18635, signal_18633, signal_18631, signal_18629}), .b ({signal_6091, signal_6090, signal_6089, signal_6088, signal_1858}), .clk ( clk ), .r ({Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730]}), .c ({signal_6735, signal_6734, signal_6733, signal_6732, signal_2019}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2005 ( .a ({signal_18247, signal_18245, signal_18243, signal_18241, signal_18239}), .b ({signal_6095, signal_6094, signal_6093, signal_6092, signal_1859}), .clk ( clk ), .r ({Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740]}), .c ({signal_6739, signal_6738, signal_6737, signal_6736, signal_2020}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2006 ( .a ({signal_18647, signal_18645, signal_18643, signal_18641, signal_18639}), .b ({signal_6099, signal_6098, signal_6097, signal_6096, signal_1860}), .clk ( clk ), .r ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750]}), .c ({signal_6743, signal_6742, signal_6741, signal_6740, signal_2021}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2008 ( .a ({signal_18657, signal_18655, signal_18653, signal_18651, signal_18649}), .b ({signal_6115, signal_6114, signal_6113, signal_6112, signal_1864}), .clk ( clk ), .r ({Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .c ({signal_6751, signal_6750, signal_6749, signal_6748, signal_2023}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2011 ( .a ({signal_18247, signal_18245, signal_18243, signal_18241, signal_18239}), .b ({signal_6119, signal_6118, signal_6117, signal_6116, signal_1865}), .clk ( clk ), .r ({Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770]}), .c ({signal_6763, signal_6762, signal_6761, signal_6760, signal_2026}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2012 ( .a ({signal_5095, signal_5094, signal_5093, signal_5092, signal_1609}), .b ({signal_6127, signal_6126, signal_6125, signal_6124, signal_1867}), .clk ( clk ), .r ({Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780]}), .c ({signal_6767, signal_6766, signal_6765, signal_6764, signal_2027}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2014 ( .a ({signal_6135, signal_6134, signal_6133, signal_6132, signal_1869}), .b ({signal_5411, signal_5410, signal_5409, signal_5408, signal_1688}), .clk ( clk ), .r ({Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790]}), .c ({signal_6775, signal_6774, signal_6773, signal_6772, signal_2029}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2015 ( .a ({signal_5087, signal_5086, signal_5085, signal_5084, signal_1607}), .b ({signal_6143, signal_6142, signal_6141, signal_6140, signal_1871}), .clk ( clk ), .r ({Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800]}), .c ({signal_6779, signal_6778, signal_6777, signal_6776, signal_2030}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2048 ( .a ({signal_6735, signal_6734, signal_6733, signal_6732, signal_2019}), .b ({signal_6911, signal_6910, signal_6909, signal_6908, signal_2063}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2052 ( .a ({signal_6763, signal_6762, signal_6761, signal_6760, signal_2026}), .b ({signal_6927, signal_6926, signal_6925, signal_6924, signal_2067}) ) ;
    buf_clk cell_3966 ( .C ( clk ), .D ( signal_18658 ), .Q ( signal_18659 ) ) ;
    buf_clk cell_3968 ( .C ( clk ), .D ( signal_18660 ), .Q ( signal_18661 ) ) ;
    buf_clk cell_3970 ( .C ( clk ), .D ( signal_18662 ), .Q ( signal_18663 ) ) ;
    buf_clk cell_3972 ( .C ( clk ), .D ( signal_18664 ), .Q ( signal_18665 ) ) ;
    buf_clk cell_3974 ( .C ( clk ), .D ( signal_18666 ), .Q ( signal_18667 ) ) ;
    buf_clk cell_3976 ( .C ( clk ), .D ( signal_18668 ), .Q ( signal_18669 ) ) ;
    buf_clk cell_3978 ( .C ( clk ), .D ( signal_18670 ), .Q ( signal_18671 ) ) ;
    buf_clk cell_3980 ( .C ( clk ), .D ( signal_18672 ), .Q ( signal_18673 ) ) ;
    buf_clk cell_3982 ( .C ( clk ), .D ( signal_18674 ), .Q ( signal_18675 ) ) ;
    buf_clk cell_3984 ( .C ( clk ), .D ( signal_18676 ), .Q ( signal_18677 ) ) ;
    buf_clk cell_3988 ( .C ( clk ), .D ( signal_18680 ), .Q ( signal_18681 ) ) ;
    buf_clk cell_3992 ( .C ( clk ), .D ( signal_18684 ), .Q ( signal_18685 ) ) ;
    buf_clk cell_3996 ( .C ( clk ), .D ( signal_18688 ), .Q ( signal_18689 ) ) ;
    buf_clk cell_4000 ( .C ( clk ), .D ( signal_18692 ), .Q ( signal_18693 ) ) ;
    buf_clk cell_4004 ( .C ( clk ), .D ( signal_18696 ), .Q ( signal_18697 ) ) ;
    buf_clk cell_4006 ( .C ( clk ), .D ( signal_18698 ), .Q ( signal_18699 ) ) ;
    buf_clk cell_4008 ( .C ( clk ), .D ( signal_18700 ), .Q ( signal_18701 ) ) ;
    buf_clk cell_4010 ( .C ( clk ), .D ( signal_18702 ), .Q ( signal_18703 ) ) ;
    buf_clk cell_4012 ( .C ( clk ), .D ( signal_18704 ), .Q ( signal_18705 ) ) ;
    buf_clk cell_4014 ( .C ( clk ), .D ( signal_18706 ), .Q ( signal_18707 ) ) ;
    buf_clk cell_4018 ( .C ( clk ), .D ( signal_18710 ), .Q ( signal_18711 ) ) ;
    buf_clk cell_4022 ( .C ( clk ), .D ( signal_18714 ), .Q ( signal_18715 ) ) ;
    buf_clk cell_4026 ( .C ( clk ), .D ( signal_18718 ), .Q ( signal_18719 ) ) ;
    buf_clk cell_4030 ( .C ( clk ), .D ( signal_18722 ), .Q ( signal_18723 ) ) ;
    buf_clk cell_4034 ( .C ( clk ), .D ( signal_18726 ), .Q ( signal_18727 ) ) ;
    buf_clk cell_4038 ( .C ( clk ), .D ( signal_18730 ), .Q ( signal_18731 ) ) ;
    buf_clk cell_4042 ( .C ( clk ), .D ( signal_18734 ), .Q ( signal_18735 ) ) ;
    buf_clk cell_4046 ( .C ( clk ), .D ( signal_18738 ), .Q ( signal_18739 ) ) ;
    buf_clk cell_4050 ( .C ( clk ), .D ( signal_18742 ), .Q ( signal_18743 ) ) ;
    buf_clk cell_4054 ( .C ( clk ), .D ( signal_18746 ), .Q ( signal_18747 ) ) ;
    buf_clk cell_4058 ( .C ( clk ), .D ( signal_18750 ), .Q ( signal_18751 ) ) ;
    buf_clk cell_4062 ( .C ( clk ), .D ( signal_18754 ), .Q ( signal_18755 ) ) ;
    buf_clk cell_4066 ( .C ( clk ), .D ( signal_18758 ), .Q ( signal_18759 ) ) ;
    buf_clk cell_4070 ( .C ( clk ), .D ( signal_18762 ), .Q ( signal_18763 ) ) ;
    buf_clk cell_4074 ( .C ( clk ), .D ( signal_18766 ), .Q ( signal_18767 ) ) ;
    buf_clk cell_4082 ( .C ( clk ), .D ( signal_18774 ), .Q ( signal_18775 ) ) ;
    buf_clk cell_4090 ( .C ( clk ), .D ( signal_18782 ), .Q ( signal_18783 ) ) ;
    buf_clk cell_4098 ( .C ( clk ), .D ( signal_18790 ), .Q ( signal_18791 ) ) ;
    buf_clk cell_4106 ( .C ( clk ), .D ( signal_18798 ), .Q ( signal_18799 ) ) ;
    buf_clk cell_4114 ( .C ( clk ), .D ( signal_18806 ), .Q ( signal_18807 ) ) ;
    buf_clk cell_4116 ( .C ( clk ), .D ( signal_18808 ), .Q ( signal_18809 ) ) ;
    buf_clk cell_4118 ( .C ( clk ), .D ( signal_18810 ), .Q ( signal_18811 ) ) ;
    buf_clk cell_4120 ( .C ( clk ), .D ( signal_18812 ), .Q ( signal_18813 ) ) ;
    buf_clk cell_4122 ( .C ( clk ), .D ( signal_18814 ), .Q ( signal_18815 ) ) ;
    buf_clk cell_4124 ( .C ( clk ), .D ( signal_18816 ), .Q ( signal_18817 ) ) ;
    buf_clk cell_4126 ( .C ( clk ), .D ( signal_18818 ), .Q ( signal_18819 ) ) ;
    buf_clk cell_4128 ( .C ( clk ), .D ( signal_18820 ), .Q ( signal_18821 ) ) ;
    buf_clk cell_4130 ( .C ( clk ), .D ( signal_18822 ), .Q ( signal_18823 ) ) ;
    buf_clk cell_4132 ( .C ( clk ), .D ( signal_18824 ), .Q ( signal_18825 ) ) ;
    buf_clk cell_4134 ( .C ( clk ), .D ( signal_18826 ), .Q ( signal_18827 ) ) ;
    buf_clk cell_4138 ( .C ( clk ), .D ( signal_18830 ), .Q ( signal_18831 ) ) ;
    buf_clk cell_4142 ( .C ( clk ), .D ( signal_18834 ), .Q ( signal_18835 ) ) ;
    buf_clk cell_4146 ( .C ( clk ), .D ( signal_18838 ), .Q ( signal_18839 ) ) ;
    buf_clk cell_4150 ( .C ( clk ), .D ( signal_18842 ), .Q ( signal_18843 ) ) ;
    buf_clk cell_4154 ( .C ( clk ), .D ( signal_18846 ), .Q ( signal_18847 ) ) ;
    buf_clk cell_4156 ( .C ( clk ), .D ( signal_18848 ), .Q ( signal_18849 ) ) ;
    buf_clk cell_4158 ( .C ( clk ), .D ( signal_18850 ), .Q ( signal_18851 ) ) ;
    buf_clk cell_4160 ( .C ( clk ), .D ( signal_18852 ), .Q ( signal_18853 ) ) ;
    buf_clk cell_4162 ( .C ( clk ), .D ( signal_18854 ), .Q ( signal_18855 ) ) ;
    buf_clk cell_4164 ( .C ( clk ), .D ( signal_18856 ), .Q ( signal_18857 ) ) ;
    buf_clk cell_4166 ( .C ( clk ), .D ( signal_18858 ), .Q ( signal_18859 ) ) ;
    buf_clk cell_4168 ( .C ( clk ), .D ( signal_18860 ), .Q ( signal_18861 ) ) ;
    buf_clk cell_4170 ( .C ( clk ), .D ( signal_18862 ), .Q ( signal_18863 ) ) ;
    buf_clk cell_4172 ( .C ( clk ), .D ( signal_18864 ), .Q ( signal_18865 ) ) ;
    buf_clk cell_4174 ( .C ( clk ), .D ( signal_18866 ), .Q ( signal_18867 ) ) ;
    buf_clk cell_4178 ( .C ( clk ), .D ( signal_18870 ), .Q ( signal_18871 ) ) ;
    buf_clk cell_4182 ( .C ( clk ), .D ( signal_18874 ), .Q ( signal_18875 ) ) ;
    buf_clk cell_4186 ( .C ( clk ), .D ( signal_18878 ), .Q ( signal_18879 ) ) ;
    buf_clk cell_4190 ( .C ( clk ), .D ( signal_18882 ), .Q ( signal_18883 ) ) ;
    buf_clk cell_4194 ( .C ( clk ), .D ( signal_18886 ), .Q ( signal_18887 ) ) ;
    buf_clk cell_4196 ( .C ( clk ), .D ( signal_18888 ), .Q ( signal_18889 ) ) ;
    buf_clk cell_4198 ( .C ( clk ), .D ( signal_18890 ), .Q ( signal_18891 ) ) ;
    buf_clk cell_4200 ( .C ( clk ), .D ( signal_18892 ), .Q ( signal_18893 ) ) ;
    buf_clk cell_4202 ( .C ( clk ), .D ( signal_18894 ), .Q ( signal_18895 ) ) ;
    buf_clk cell_4204 ( .C ( clk ), .D ( signal_18896 ), .Q ( signal_18897 ) ) ;
    buf_clk cell_4206 ( .C ( clk ), .D ( signal_18898 ), .Q ( signal_18899 ) ) ;
    buf_clk cell_4208 ( .C ( clk ), .D ( signal_18900 ), .Q ( signal_18901 ) ) ;
    buf_clk cell_4210 ( .C ( clk ), .D ( signal_18902 ), .Q ( signal_18903 ) ) ;
    buf_clk cell_4212 ( .C ( clk ), .D ( signal_18904 ), .Q ( signal_18905 ) ) ;
    buf_clk cell_4214 ( .C ( clk ), .D ( signal_18906 ), .Q ( signal_18907 ) ) ;
    buf_clk cell_4216 ( .C ( clk ), .D ( signal_18908 ), .Q ( signal_18909 ) ) ;
    buf_clk cell_4218 ( .C ( clk ), .D ( signal_18910 ), .Q ( signal_18911 ) ) ;
    buf_clk cell_4220 ( .C ( clk ), .D ( signal_18912 ), .Q ( signal_18913 ) ) ;
    buf_clk cell_4222 ( .C ( clk ), .D ( signal_18914 ), .Q ( signal_18915 ) ) ;
    buf_clk cell_4224 ( .C ( clk ), .D ( signal_18916 ), .Q ( signal_18917 ) ) ;
    buf_clk cell_4226 ( .C ( clk ), .D ( signal_18918 ), .Q ( signal_18919 ) ) ;
    buf_clk cell_4228 ( .C ( clk ), .D ( signal_18920 ), .Q ( signal_18921 ) ) ;
    buf_clk cell_4230 ( .C ( clk ), .D ( signal_18922 ), .Q ( signal_18923 ) ) ;
    buf_clk cell_4232 ( .C ( clk ), .D ( signal_18924 ), .Q ( signal_18925 ) ) ;
    buf_clk cell_4234 ( .C ( clk ), .D ( signal_18926 ), .Q ( signal_18927 ) ) ;
    buf_clk cell_4236 ( .C ( clk ), .D ( signal_18928 ), .Q ( signal_18929 ) ) ;
    buf_clk cell_4238 ( .C ( clk ), .D ( signal_18930 ), .Q ( signal_18931 ) ) ;
    buf_clk cell_4240 ( .C ( clk ), .D ( signal_18932 ), .Q ( signal_18933 ) ) ;
    buf_clk cell_4242 ( .C ( clk ), .D ( signal_18934 ), .Q ( signal_18935 ) ) ;
    buf_clk cell_4244 ( .C ( clk ), .D ( signal_18936 ), .Q ( signal_18937 ) ) ;
    buf_clk cell_4248 ( .C ( clk ), .D ( signal_18940 ), .Q ( signal_18941 ) ) ;
    buf_clk cell_4252 ( .C ( clk ), .D ( signal_18944 ), .Q ( signal_18945 ) ) ;
    buf_clk cell_4256 ( .C ( clk ), .D ( signal_18948 ), .Q ( signal_18949 ) ) ;
    buf_clk cell_4260 ( .C ( clk ), .D ( signal_18952 ), .Q ( signal_18953 ) ) ;
    buf_clk cell_4264 ( .C ( clk ), .D ( signal_18956 ), .Q ( signal_18957 ) ) ;
    buf_clk cell_4266 ( .C ( clk ), .D ( signal_18958 ), .Q ( signal_18959 ) ) ;
    buf_clk cell_4268 ( .C ( clk ), .D ( signal_18960 ), .Q ( signal_18961 ) ) ;
    buf_clk cell_4270 ( .C ( clk ), .D ( signal_18962 ), .Q ( signal_18963 ) ) ;
    buf_clk cell_4272 ( .C ( clk ), .D ( signal_18964 ), .Q ( signal_18965 ) ) ;
    buf_clk cell_4274 ( .C ( clk ), .D ( signal_18966 ), .Q ( signal_18967 ) ) ;
    buf_clk cell_4276 ( .C ( clk ), .D ( signal_18968 ), .Q ( signal_18969 ) ) ;
    buf_clk cell_4278 ( .C ( clk ), .D ( signal_18970 ), .Q ( signal_18971 ) ) ;
    buf_clk cell_4280 ( .C ( clk ), .D ( signal_18972 ), .Q ( signal_18973 ) ) ;
    buf_clk cell_4282 ( .C ( clk ), .D ( signal_18974 ), .Q ( signal_18975 ) ) ;
    buf_clk cell_4284 ( .C ( clk ), .D ( signal_18976 ), .Q ( signal_18977 ) ) ;
    buf_clk cell_4286 ( .C ( clk ), .D ( signal_18978 ), .Q ( signal_18979 ) ) ;
    buf_clk cell_4288 ( .C ( clk ), .D ( signal_18980 ), .Q ( signal_18981 ) ) ;
    buf_clk cell_4290 ( .C ( clk ), .D ( signal_18982 ), .Q ( signal_18983 ) ) ;
    buf_clk cell_4292 ( .C ( clk ), .D ( signal_18984 ), .Q ( signal_18985 ) ) ;
    buf_clk cell_4294 ( .C ( clk ), .D ( signal_18986 ), .Q ( signal_18987 ) ) ;
    buf_clk cell_4296 ( .C ( clk ), .D ( signal_18988 ), .Q ( signal_18989 ) ) ;
    buf_clk cell_4298 ( .C ( clk ), .D ( signal_18990 ), .Q ( signal_18991 ) ) ;
    buf_clk cell_4300 ( .C ( clk ), .D ( signal_18992 ), .Q ( signal_18993 ) ) ;
    buf_clk cell_4302 ( .C ( clk ), .D ( signal_18994 ), .Q ( signal_18995 ) ) ;
    buf_clk cell_4304 ( .C ( clk ), .D ( signal_18996 ), .Q ( signal_18997 ) ) ;
    buf_clk cell_4308 ( .C ( clk ), .D ( signal_19000 ), .Q ( signal_19001 ) ) ;
    buf_clk cell_4312 ( .C ( clk ), .D ( signal_19004 ), .Q ( signal_19005 ) ) ;
    buf_clk cell_4316 ( .C ( clk ), .D ( signal_19008 ), .Q ( signal_19009 ) ) ;
    buf_clk cell_4320 ( .C ( clk ), .D ( signal_19012 ), .Q ( signal_19013 ) ) ;
    buf_clk cell_4324 ( .C ( clk ), .D ( signal_19016 ), .Q ( signal_19017 ) ) ;
    buf_clk cell_4326 ( .C ( clk ), .D ( signal_19018 ), .Q ( signal_19019 ) ) ;
    buf_clk cell_4328 ( .C ( clk ), .D ( signal_19020 ), .Q ( signal_19021 ) ) ;
    buf_clk cell_4330 ( .C ( clk ), .D ( signal_19022 ), .Q ( signal_19023 ) ) ;
    buf_clk cell_4332 ( .C ( clk ), .D ( signal_19024 ), .Q ( signal_19025 ) ) ;
    buf_clk cell_4334 ( .C ( clk ), .D ( signal_19026 ), .Q ( signal_19027 ) ) ;
    buf_clk cell_4336 ( .C ( clk ), .D ( signal_19028 ), .Q ( signal_19029 ) ) ;
    buf_clk cell_4338 ( .C ( clk ), .D ( signal_19030 ), .Q ( signal_19031 ) ) ;
    buf_clk cell_4340 ( .C ( clk ), .D ( signal_19032 ), .Q ( signal_19033 ) ) ;
    buf_clk cell_4342 ( .C ( clk ), .D ( signal_19034 ), .Q ( signal_19035 ) ) ;
    buf_clk cell_4344 ( .C ( clk ), .D ( signal_19036 ), .Q ( signal_19037 ) ) ;
    buf_clk cell_4348 ( .C ( clk ), .D ( signal_19040 ), .Q ( signal_19041 ) ) ;
    buf_clk cell_4352 ( .C ( clk ), .D ( signal_19044 ), .Q ( signal_19045 ) ) ;
    buf_clk cell_4356 ( .C ( clk ), .D ( signal_19048 ), .Q ( signal_19049 ) ) ;
    buf_clk cell_4360 ( .C ( clk ), .D ( signal_19052 ), .Q ( signal_19053 ) ) ;
    buf_clk cell_4364 ( .C ( clk ), .D ( signal_19056 ), .Q ( signal_19057 ) ) ;
    buf_clk cell_4368 ( .C ( clk ), .D ( signal_19060 ), .Q ( signal_19061 ) ) ;
    buf_clk cell_4372 ( .C ( clk ), .D ( signal_19064 ), .Q ( signal_19065 ) ) ;
    buf_clk cell_4376 ( .C ( clk ), .D ( signal_19068 ), .Q ( signal_19069 ) ) ;
    buf_clk cell_4380 ( .C ( clk ), .D ( signal_19072 ), .Q ( signal_19073 ) ) ;
    buf_clk cell_4384 ( .C ( clk ), .D ( signal_19076 ), .Q ( signal_19077 ) ) ;
    buf_clk cell_4388 ( .C ( clk ), .D ( signal_19080 ), .Q ( signal_19081 ) ) ;
    buf_clk cell_4392 ( .C ( clk ), .D ( signal_19084 ), .Q ( signal_19085 ) ) ;
    buf_clk cell_4396 ( .C ( clk ), .D ( signal_19088 ), .Q ( signal_19089 ) ) ;
    buf_clk cell_4400 ( .C ( clk ), .D ( signal_19092 ), .Q ( signal_19093 ) ) ;
    buf_clk cell_4404 ( .C ( clk ), .D ( signal_19096 ), .Q ( signal_19097 ) ) ;
    buf_clk cell_4408 ( .C ( clk ), .D ( signal_19100 ), .Q ( signal_19101 ) ) ;
    buf_clk cell_4412 ( .C ( clk ), .D ( signal_19104 ), .Q ( signal_19105 ) ) ;
    buf_clk cell_4416 ( .C ( clk ), .D ( signal_19108 ), .Q ( signal_19109 ) ) ;
    buf_clk cell_4420 ( .C ( clk ), .D ( signal_19112 ), .Q ( signal_19113 ) ) ;
    buf_clk cell_4424 ( .C ( clk ), .D ( signal_19116 ), .Q ( signal_19117 ) ) ;
    buf_clk cell_4426 ( .C ( clk ), .D ( signal_19118 ), .Q ( signal_19119 ) ) ;
    buf_clk cell_4428 ( .C ( clk ), .D ( signal_19120 ), .Q ( signal_19121 ) ) ;
    buf_clk cell_4430 ( .C ( clk ), .D ( signal_19122 ), .Q ( signal_19123 ) ) ;
    buf_clk cell_4432 ( .C ( clk ), .D ( signal_19124 ), .Q ( signal_19125 ) ) ;
    buf_clk cell_4434 ( .C ( clk ), .D ( signal_19126 ), .Q ( signal_19127 ) ) ;
    buf_clk cell_4436 ( .C ( clk ), .D ( signal_19128 ), .Q ( signal_19129 ) ) ;
    buf_clk cell_4438 ( .C ( clk ), .D ( signal_19130 ), .Q ( signal_19131 ) ) ;
    buf_clk cell_4440 ( .C ( clk ), .D ( signal_19132 ), .Q ( signal_19133 ) ) ;
    buf_clk cell_4442 ( .C ( clk ), .D ( signal_19134 ), .Q ( signal_19135 ) ) ;
    buf_clk cell_4444 ( .C ( clk ), .D ( signal_19136 ), .Q ( signal_19137 ) ) ;
    buf_clk cell_4446 ( .C ( clk ), .D ( signal_19138 ), .Q ( signal_19139 ) ) ;
    buf_clk cell_4448 ( .C ( clk ), .D ( signal_19140 ), .Q ( signal_19141 ) ) ;
    buf_clk cell_4450 ( .C ( clk ), .D ( signal_19142 ), .Q ( signal_19143 ) ) ;
    buf_clk cell_4452 ( .C ( clk ), .D ( signal_19144 ), .Q ( signal_19145 ) ) ;
    buf_clk cell_4454 ( .C ( clk ), .D ( signal_19146 ), .Q ( signal_19147 ) ) ;
    buf_clk cell_4456 ( .C ( clk ), .D ( signal_19148 ), .Q ( signal_19149 ) ) ;
    buf_clk cell_4458 ( .C ( clk ), .D ( signal_19150 ), .Q ( signal_19151 ) ) ;
    buf_clk cell_4460 ( .C ( clk ), .D ( signal_19152 ), .Q ( signal_19153 ) ) ;
    buf_clk cell_4462 ( .C ( clk ), .D ( signal_19154 ), .Q ( signal_19155 ) ) ;
    buf_clk cell_4464 ( .C ( clk ), .D ( signal_19156 ), .Q ( signal_19157 ) ) ;
    buf_clk cell_4466 ( .C ( clk ), .D ( signal_19158 ), .Q ( signal_19159 ) ) ;
    buf_clk cell_4468 ( .C ( clk ), .D ( signal_19160 ), .Q ( signal_19161 ) ) ;
    buf_clk cell_4470 ( .C ( clk ), .D ( signal_19162 ), .Q ( signal_19163 ) ) ;
    buf_clk cell_4472 ( .C ( clk ), .D ( signal_19164 ), .Q ( signal_19165 ) ) ;
    buf_clk cell_4474 ( .C ( clk ), .D ( signal_19166 ), .Q ( signal_19167 ) ) ;
    buf_clk cell_4478 ( .C ( clk ), .D ( signal_19170 ), .Q ( signal_19171 ) ) ;
    buf_clk cell_4482 ( .C ( clk ), .D ( signal_19174 ), .Q ( signal_19175 ) ) ;
    buf_clk cell_4486 ( .C ( clk ), .D ( signal_19178 ), .Q ( signal_19179 ) ) ;
    buf_clk cell_4490 ( .C ( clk ), .D ( signal_19182 ), .Q ( signal_19183 ) ) ;
    buf_clk cell_4494 ( .C ( clk ), .D ( signal_19186 ), .Q ( signal_19187 ) ) ;
    buf_clk cell_4498 ( .C ( clk ), .D ( signal_19190 ), .Q ( signal_19191 ) ) ;
    buf_clk cell_4502 ( .C ( clk ), .D ( signal_19194 ), .Q ( signal_19195 ) ) ;
    buf_clk cell_4506 ( .C ( clk ), .D ( signal_19198 ), .Q ( signal_19199 ) ) ;
    buf_clk cell_4510 ( .C ( clk ), .D ( signal_19202 ), .Q ( signal_19203 ) ) ;
    buf_clk cell_4514 ( .C ( clk ), .D ( signal_19206 ), .Q ( signal_19207 ) ) ;
    buf_clk cell_4518 ( .C ( clk ), .D ( signal_19210 ), .Q ( signal_19211 ) ) ;
    buf_clk cell_4522 ( .C ( clk ), .D ( signal_19214 ), .Q ( signal_19215 ) ) ;
    buf_clk cell_4526 ( .C ( clk ), .D ( signal_19218 ), .Q ( signal_19219 ) ) ;
    buf_clk cell_4530 ( .C ( clk ), .D ( signal_19222 ), .Q ( signal_19223 ) ) ;
    buf_clk cell_4534 ( .C ( clk ), .D ( signal_19226 ), .Q ( signal_19227 ) ) ;
    buf_clk cell_4536 ( .C ( clk ), .D ( signal_19228 ), .Q ( signal_19229 ) ) ;
    buf_clk cell_4538 ( .C ( clk ), .D ( signal_19230 ), .Q ( signal_19231 ) ) ;
    buf_clk cell_4540 ( .C ( clk ), .D ( signal_19232 ), .Q ( signal_19233 ) ) ;
    buf_clk cell_4542 ( .C ( clk ), .D ( signal_19234 ), .Q ( signal_19235 ) ) ;
    buf_clk cell_4544 ( .C ( clk ), .D ( signal_19236 ), .Q ( signal_19237 ) ) ;
    buf_clk cell_4548 ( .C ( clk ), .D ( signal_19240 ), .Q ( signal_19241 ) ) ;
    buf_clk cell_4552 ( .C ( clk ), .D ( signal_19244 ), .Q ( signal_19245 ) ) ;
    buf_clk cell_4556 ( .C ( clk ), .D ( signal_19248 ), .Q ( signal_19249 ) ) ;
    buf_clk cell_4560 ( .C ( clk ), .D ( signal_19252 ), .Q ( signal_19253 ) ) ;
    buf_clk cell_4564 ( .C ( clk ), .D ( signal_19256 ), .Q ( signal_19257 ) ) ;
    buf_clk cell_4566 ( .C ( clk ), .D ( signal_19258 ), .Q ( signal_19259 ) ) ;
    buf_clk cell_4568 ( .C ( clk ), .D ( signal_19260 ), .Q ( signal_19261 ) ) ;
    buf_clk cell_4570 ( .C ( clk ), .D ( signal_19262 ), .Q ( signal_19263 ) ) ;
    buf_clk cell_4572 ( .C ( clk ), .D ( signal_19264 ), .Q ( signal_19265 ) ) ;
    buf_clk cell_4574 ( .C ( clk ), .D ( signal_19266 ), .Q ( signal_19267 ) ) ;
    buf_clk cell_4576 ( .C ( clk ), .D ( signal_19268 ), .Q ( signal_19269 ) ) ;
    buf_clk cell_4578 ( .C ( clk ), .D ( signal_19270 ), .Q ( signal_19271 ) ) ;
    buf_clk cell_4580 ( .C ( clk ), .D ( signal_19272 ), .Q ( signal_19273 ) ) ;
    buf_clk cell_4582 ( .C ( clk ), .D ( signal_19274 ), .Q ( signal_19275 ) ) ;
    buf_clk cell_4584 ( .C ( clk ), .D ( signal_19276 ), .Q ( signal_19277 ) ) ;
    buf_clk cell_4586 ( .C ( clk ), .D ( signal_19278 ), .Q ( signal_19279 ) ) ;
    buf_clk cell_4588 ( .C ( clk ), .D ( signal_19280 ), .Q ( signal_19281 ) ) ;
    buf_clk cell_4590 ( .C ( clk ), .D ( signal_19282 ), .Q ( signal_19283 ) ) ;
    buf_clk cell_4592 ( .C ( clk ), .D ( signal_19284 ), .Q ( signal_19285 ) ) ;
    buf_clk cell_4594 ( .C ( clk ), .D ( signal_19286 ), .Q ( signal_19287 ) ) ;
    buf_clk cell_4596 ( .C ( clk ), .D ( signal_19288 ), .Q ( signal_19289 ) ) ;
    buf_clk cell_4598 ( .C ( clk ), .D ( signal_19290 ), .Q ( signal_19291 ) ) ;
    buf_clk cell_4600 ( .C ( clk ), .D ( signal_19292 ), .Q ( signal_19293 ) ) ;
    buf_clk cell_4602 ( .C ( clk ), .D ( signal_19294 ), .Q ( signal_19295 ) ) ;
    buf_clk cell_4604 ( .C ( clk ), .D ( signal_19296 ), .Q ( signal_19297 ) ) ;
    buf_clk cell_4606 ( .C ( clk ), .D ( signal_19298 ), .Q ( signal_19299 ) ) ;
    buf_clk cell_4608 ( .C ( clk ), .D ( signal_19300 ), .Q ( signal_19301 ) ) ;
    buf_clk cell_4610 ( .C ( clk ), .D ( signal_19302 ), .Q ( signal_19303 ) ) ;
    buf_clk cell_4612 ( .C ( clk ), .D ( signal_19304 ), .Q ( signal_19305 ) ) ;
    buf_clk cell_4614 ( .C ( clk ), .D ( signal_19306 ), .Q ( signal_19307 ) ) ;
    buf_clk cell_4618 ( .C ( clk ), .D ( signal_19310 ), .Q ( signal_19311 ) ) ;
    buf_clk cell_4622 ( .C ( clk ), .D ( signal_19314 ), .Q ( signal_19315 ) ) ;
    buf_clk cell_4626 ( .C ( clk ), .D ( signal_19318 ), .Q ( signal_19319 ) ) ;
    buf_clk cell_4630 ( .C ( clk ), .D ( signal_19322 ), .Q ( signal_19323 ) ) ;
    buf_clk cell_4634 ( .C ( clk ), .D ( signal_19326 ), .Q ( signal_19327 ) ) ;
    buf_clk cell_4638 ( .C ( clk ), .D ( signal_19330 ), .Q ( signal_19331 ) ) ;
    buf_clk cell_4642 ( .C ( clk ), .D ( signal_19334 ), .Q ( signal_19335 ) ) ;
    buf_clk cell_4646 ( .C ( clk ), .D ( signal_19338 ), .Q ( signal_19339 ) ) ;
    buf_clk cell_4650 ( .C ( clk ), .D ( signal_19342 ), .Q ( signal_19343 ) ) ;
    buf_clk cell_4654 ( .C ( clk ), .D ( signal_19346 ), .Q ( signal_19347 ) ) ;
    buf_clk cell_4656 ( .C ( clk ), .D ( signal_19348 ), .Q ( signal_19349 ) ) ;
    buf_clk cell_4658 ( .C ( clk ), .D ( signal_19350 ), .Q ( signal_19351 ) ) ;
    buf_clk cell_4660 ( .C ( clk ), .D ( signal_19352 ), .Q ( signal_19353 ) ) ;
    buf_clk cell_4662 ( .C ( clk ), .D ( signal_19354 ), .Q ( signal_19355 ) ) ;
    buf_clk cell_4664 ( .C ( clk ), .D ( signal_19356 ), .Q ( signal_19357 ) ) ;
    buf_clk cell_4668 ( .C ( clk ), .D ( signal_19360 ), .Q ( signal_19361 ) ) ;
    buf_clk cell_4672 ( .C ( clk ), .D ( signal_19364 ), .Q ( signal_19365 ) ) ;
    buf_clk cell_4676 ( .C ( clk ), .D ( signal_19368 ), .Q ( signal_19369 ) ) ;
    buf_clk cell_4680 ( .C ( clk ), .D ( signal_19372 ), .Q ( signal_19373 ) ) ;
    buf_clk cell_4684 ( .C ( clk ), .D ( signal_19376 ), .Q ( signal_19377 ) ) ;
    buf_clk cell_4686 ( .C ( clk ), .D ( signal_19378 ), .Q ( signal_19379 ) ) ;
    buf_clk cell_4688 ( .C ( clk ), .D ( signal_19380 ), .Q ( signal_19381 ) ) ;
    buf_clk cell_4690 ( .C ( clk ), .D ( signal_19382 ), .Q ( signal_19383 ) ) ;
    buf_clk cell_4692 ( .C ( clk ), .D ( signal_19384 ), .Q ( signal_19385 ) ) ;
    buf_clk cell_4694 ( .C ( clk ), .D ( signal_19386 ), .Q ( signal_19387 ) ) ;
    buf_clk cell_4696 ( .C ( clk ), .D ( signal_19388 ), .Q ( signal_19389 ) ) ;
    buf_clk cell_4698 ( .C ( clk ), .D ( signal_19390 ), .Q ( signal_19391 ) ) ;
    buf_clk cell_4700 ( .C ( clk ), .D ( signal_19392 ), .Q ( signal_19393 ) ) ;
    buf_clk cell_4702 ( .C ( clk ), .D ( signal_19394 ), .Q ( signal_19395 ) ) ;
    buf_clk cell_4704 ( .C ( clk ), .D ( signal_19396 ), .Q ( signal_19397 ) ) ;
    buf_clk cell_4708 ( .C ( clk ), .D ( signal_19400 ), .Q ( signal_19401 ) ) ;
    buf_clk cell_4712 ( .C ( clk ), .D ( signal_19404 ), .Q ( signal_19405 ) ) ;
    buf_clk cell_4716 ( .C ( clk ), .D ( signal_19408 ), .Q ( signal_19409 ) ) ;
    buf_clk cell_4720 ( .C ( clk ), .D ( signal_19412 ), .Q ( signal_19413 ) ) ;
    buf_clk cell_4724 ( .C ( clk ), .D ( signal_19416 ), .Q ( signal_19417 ) ) ;
    buf_clk cell_4728 ( .C ( clk ), .D ( signal_19420 ), .Q ( signal_19421 ) ) ;
    buf_clk cell_4732 ( .C ( clk ), .D ( signal_19424 ), .Q ( signal_19425 ) ) ;
    buf_clk cell_4736 ( .C ( clk ), .D ( signal_19428 ), .Q ( signal_19429 ) ) ;
    buf_clk cell_4740 ( .C ( clk ), .D ( signal_19432 ), .Q ( signal_19433 ) ) ;
    buf_clk cell_4744 ( .C ( clk ), .D ( signal_19436 ), .Q ( signal_19437 ) ) ;
    buf_clk cell_4748 ( .C ( clk ), .D ( signal_19440 ), .Q ( signal_19441 ) ) ;
    buf_clk cell_4752 ( .C ( clk ), .D ( signal_19444 ), .Q ( signal_19445 ) ) ;
    buf_clk cell_4756 ( .C ( clk ), .D ( signal_19448 ), .Q ( signal_19449 ) ) ;
    buf_clk cell_4760 ( .C ( clk ), .D ( signal_19452 ), .Q ( signal_19453 ) ) ;
    buf_clk cell_4764 ( .C ( clk ), .D ( signal_19456 ), .Q ( signal_19457 ) ) ;
    buf_clk cell_4766 ( .C ( clk ), .D ( signal_19458 ), .Q ( signal_19459 ) ) ;
    buf_clk cell_4768 ( .C ( clk ), .D ( signal_19460 ), .Q ( signal_19461 ) ) ;
    buf_clk cell_4770 ( .C ( clk ), .D ( signal_19462 ), .Q ( signal_19463 ) ) ;
    buf_clk cell_4772 ( .C ( clk ), .D ( signal_19464 ), .Q ( signal_19465 ) ) ;
    buf_clk cell_4774 ( .C ( clk ), .D ( signal_19466 ), .Q ( signal_19467 ) ) ;
    buf_clk cell_4778 ( .C ( clk ), .D ( signal_19470 ), .Q ( signal_19471 ) ) ;
    buf_clk cell_4782 ( .C ( clk ), .D ( signal_19474 ), .Q ( signal_19475 ) ) ;
    buf_clk cell_4786 ( .C ( clk ), .D ( signal_19478 ), .Q ( signal_19479 ) ) ;
    buf_clk cell_4790 ( .C ( clk ), .D ( signal_19482 ), .Q ( signal_19483 ) ) ;
    buf_clk cell_4794 ( .C ( clk ), .D ( signal_19486 ), .Q ( signal_19487 ) ) ;
    buf_clk cell_4798 ( .C ( clk ), .D ( signal_19490 ), .Q ( signal_19491 ) ) ;
    buf_clk cell_4802 ( .C ( clk ), .D ( signal_19494 ), .Q ( signal_19495 ) ) ;
    buf_clk cell_4806 ( .C ( clk ), .D ( signal_19498 ), .Q ( signal_19499 ) ) ;
    buf_clk cell_4810 ( .C ( clk ), .D ( signal_19502 ), .Q ( signal_19503 ) ) ;
    buf_clk cell_4814 ( .C ( clk ), .D ( signal_19506 ), .Q ( signal_19507 ) ) ;
    buf_clk cell_4816 ( .C ( clk ), .D ( signal_19508 ), .Q ( signal_19509 ) ) ;
    buf_clk cell_4818 ( .C ( clk ), .D ( signal_19510 ), .Q ( signal_19511 ) ) ;
    buf_clk cell_4820 ( .C ( clk ), .D ( signal_19512 ), .Q ( signal_19513 ) ) ;
    buf_clk cell_4822 ( .C ( clk ), .D ( signal_19514 ), .Q ( signal_19515 ) ) ;
    buf_clk cell_4824 ( .C ( clk ), .D ( signal_19516 ), .Q ( signal_19517 ) ) ;
    buf_clk cell_4828 ( .C ( clk ), .D ( signal_19520 ), .Q ( signal_19521 ) ) ;
    buf_clk cell_4832 ( .C ( clk ), .D ( signal_19524 ), .Q ( signal_19525 ) ) ;
    buf_clk cell_4836 ( .C ( clk ), .D ( signal_19528 ), .Q ( signal_19529 ) ) ;
    buf_clk cell_4840 ( .C ( clk ), .D ( signal_19532 ), .Q ( signal_19533 ) ) ;
    buf_clk cell_4844 ( .C ( clk ), .D ( signal_19536 ), .Q ( signal_19537 ) ) ;
    buf_clk cell_4846 ( .C ( clk ), .D ( signal_19538 ), .Q ( signal_19539 ) ) ;
    buf_clk cell_4848 ( .C ( clk ), .D ( signal_19540 ), .Q ( signal_19541 ) ) ;
    buf_clk cell_4850 ( .C ( clk ), .D ( signal_19542 ), .Q ( signal_19543 ) ) ;
    buf_clk cell_4852 ( .C ( clk ), .D ( signal_19544 ), .Q ( signal_19545 ) ) ;
    buf_clk cell_4854 ( .C ( clk ), .D ( signal_19546 ), .Q ( signal_19547 ) ) ;
    buf_clk cell_4856 ( .C ( clk ), .D ( signal_19548 ), .Q ( signal_19549 ) ) ;
    buf_clk cell_4858 ( .C ( clk ), .D ( signal_19550 ), .Q ( signal_19551 ) ) ;
    buf_clk cell_4860 ( .C ( clk ), .D ( signal_19552 ), .Q ( signal_19553 ) ) ;
    buf_clk cell_4862 ( .C ( clk ), .D ( signal_19554 ), .Q ( signal_19555 ) ) ;
    buf_clk cell_4864 ( .C ( clk ), .D ( signal_19556 ), .Q ( signal_19557 ) ) ;
    buf_clk cell_4866 ( .C ( clk ), .D ( signal_19558 ), .Q ( signal_19559 ) ) ;
    buf_clk cell_4868 ( .C ( clk ), .D ( signal_19560 ), .Q ( signal_19561 ) ) ;
    buf_clk cell_4870 ( .C ( clk ), .D ( signal_19562 ), .Q ( signal_19563 ) ) ;
    buf_clk cell_4872 ( .C ( clk ), .D ( signal_19564 ), .Q ( signal_19565 ) ) ;
    buf_clk cell_4874 ( .C ( clk ), .D ( signal_19566 ), .Q ( signal_19567 ) ) ;
    buf_clk cell_4878 ( .C ( clk ), .D ( signal_19570 ), .Q ( signal_19571 ) ) ;
    buf_clk cell_4882 ( .C ( clk ), .D ( signal_19574 ), .Q ( signal_19575 ) ) ;
    buf_clk cell_4886 ( .C ( clk ), .D ( signal_19578 ), .Q ( signal_19579 ) ) ;
    buf_clk cell_4890 ( .C ( clk ), .D ( signal_19582 ), .Q ( signal_19583 ) ) ;
    buf_clk cell_4894 ( .C ( clk ), .D ( signal_19586 ), .Q ( signal_19587 ) ) ;
    buf_clk cell_4908 ( .C ( clk ), .D ( signal_19600 ), .Q ( signal_19601 ) ) ;
    buf_clk cell_4914 ( .C ( clk ), .D ( signal_19606 ), .Q ( signal_19607 ) ) ;
    buf_clk cell_4920 ( .C ( clk ), .D ( signal_19612 ), .Q ( signal_19613 ) ) ;
    buf_clk cell_4926 ( .C ( clk ), .D ( signal_19618 ), .Q ( signal_19619 ) ) ;
    buf_clk cell_4932 ( .C ( clk ), .D ( signal_19624 ), .Q ( signal_19625 ) ) ;
    buf_clk cell_4938 ( .C ( clk ), .D ( signal_19630 ), .Q ( signal_19631 ) ) ;
    buf_clk cell_4944 ( .C ( clk ), .D ( signal_19636 ), .Q ( signal_19637 ) ) ;
    buf_clk cell_4950 ( .C ( clk ), .D ( signal_19642 ), .Q ( signal_19643 ) ) ;
    buf_clk cell_4956 ( .C ( clk ), .D ( signal_19648 ), .Q ( signal_19649 ) ) ;
    buf_clk cell_4962 ( .C ( clk ), .D ( signal_19654 ), .Q ( signal_19655 ) ) ;
    buf_clk cell_4968 ( .C ( clk ), .D ( signal_19660 ), .Q ( signal_19661 ) ) ;
    buf_clk cell_4974 ( .C ( clk ), .D ( signal_19666 ), .Q ( signal_19667 ) ) ;
    buf_clk cell_4980 ( .C ( clk ), .D ( signal_19672 ), .Q ( signal_19673 ) ) ;
    buf_clk cell_4986 ( .C ( clk ), .D ( signal_19678 ), .Q ( signal_19679 ) ) ;
    buf_clk cell_4992 ( .C ( clk ), .D ( signal_19684 ), .Q ( signal_19685 ) ) ;
    buf_clk cell_4996 ( .C ( clk ), .D ( signal_19688 ), .Q ( signal_19689 ) ) ;
    buf_clk cell_5000 ( .C ( clk ), .D ( signal_19692 ), .Q ( signal_19693 ) ) ;
    buf_clk cell_5004 ( .C ( clk ), .D ( signal_19696 ), .Q ( signal_19697 ) ) ;
    buf_clk cell_5008 ( .C ( clk ), .D ( signal_19700 ), .Q ( signal_19701 ) ) ;
    buf_clk cell_5012 ( .C ( clk ), .D ( signal_19704 ), .Q ( signal_19705 ) ) ;
    buf_clk cell_5018 ( .C ( clk ), .D ( signal_19710 ), .Q ( signal_19711 ) ) ;
    buf_clk cell_5024 ( .C ( clk ), .D ( signal_19716 ), .Q ( signal_19717 ) ) ;
    buf_clk cell_5030 ( .C ( clk ), .D ( signal_19722 ), .Q ( signal_19723 ) ) ;
    buf_clk cell_5036 ( .C ( clk ), .D ( signal_19728 ), .Q ( signal_19729 ) ) ;
    buf_clk cell_5042 ( .C ( clk ), .D ( signal_19734 ), .Q ( signal_19735 ) ) ;
    buf_clk cell_5046 ( .C ( clk ), .D ( signal_19738 ), .Q ( signal_19739 ) ) ;
    buf_clk cell_5050 ( .C ( clk ), .D ( signal_19742 ), .Q ( signal_19743 ) ) ;
    buf_clk cell_5054 ( .C ( clk ), .D ( signal_19746 ), .Q ( signal_19747 ) ) ;
    buf_clk cell_5058 ( .C ( clk ), .D ( signal_19750 ), .Q ( signal_19751 ) ) ;
    buf_clk cell_5062 ( .C ( clk ), .D ( signal_19754 ), .Q ( signal_19755 ) ) ;
    buf_clk cell_5066 ( .C ( clk ), .D ( signal_19758 ), .Q ( signal_19759 ) ) ;
    buf_clk cell_5070 ( .C ( clk ), .D ( signal_19762 ), .Q ( signal_19763 ) ) ;
    buf_clk cell_5074 ( .C ( clk ), .D ( signal_19766 ), .Q ( signal_19767 ) ) ;
    buf_clk cell_5078 ( .C ( clk ), .D ( signal_19770 ), .Q ( signal_19771 ) ) ;
    buf_clk cell_5082 ( .C ( clk ), .D ( signal_19774 ), .Q ( signal_19775 ) ) ;
    buf_clk cell_5086 ( .C ( clk ), .D ( signal_19778 ), .Q ( signal_19779 ) ) ;
    buf_clk cell_5090 ( .C ( clk ), .D ( signal_19782 ), .Q ( signal_19783 ) ) ;
    buf_clk cell_5094 ( .C ( clk ), .D ( signal_19786 ), .Q ( signal_19787 ) ) ;
    buf_clk cell_5098 ( .C ( clk ), .D ( signal_19790 ), .Q ( signal_19791 ) ) ;
    buf_clk cell_5102 ( .C ( clk ), .D ( signal_19794 ), .Q ( signal_19795 ) ) ;
    buf_clk cell_5106 ( .C ( clk ), .D ( signal_19798 ), .Q ( signal_19799 ) ) ;
    buf_clk cell_5110 ( .C ( clk ), .D ( signal_19802 ), .Q ( signal_19803 ) ) ;
    buf_clk cell_5114 ( .C ( clk ), .D ( signal_19806 ), .Q ( signal_19807 ) ) ;
    buf_clk cell_5118 ( .C ( clk ), .D ( signal_19810 ), .Q ( signal_19811 ) ) ;
    buf_clk cell_5122 ( .C ( clk ), .D ( signal_19814 ), .Q ( signal_19815 ) ) ;
    buf_clk cell_5126 ( .C ( clk ), .D ( signal_19818 ), .Q ( signal_19819 ) ) ;
    buf_clk cell_5130 ( .C ( clk ), .D ( signal_19822 ), .Q ( signal_19823 ) ) ;
    buf_clk cell_5134 ( .C ( clk ), .D ( signal_19826 ), .Q ( signal_19827 ) ) ;
    buf_clk cell_5138 ( .C ( clk ), .D ( signal_19830 ), .Q ( signal_19831 ) ) ;
    buf_clk cell_5142 ( .C ( clk ), .D ( signal_19834 ), .Q ( signal_19835 ) ) ;
    buf_clk cell_5148 ( .C ( clk ), .D ( signal_19840 ), .Q ( signal_19841 ) ) ;
    buf_clk cell_5154 ( .C ( clk ), .D ( signal_19846 ), .Q ( signal_19847 ) ) ;
    buf_clk cell_5160 ( .C ( clk ), .D ( signal_19852 ), .Q ( signal_19853 ) ) ;
    buf_clk cell_5166 ( .C ( clk ), .D ( signal_19858 ), .Q ( signal_19859 ) ) ;
    buf_clk cell_5172 ( .C ( clk ), .D ( signal_19864 ), .Q ( signal_19865 ) ) ;
    buf_clk cell_5176 ( .C ( clk ), .D ( signal_19868 ), .Q ( signal_19869 ) ) ;
    buf_clk cell_5180 ( .C ( clk ), .D ( signal_19872 ), .Q ( signal_19873 ) ) ;
    buf_clk cell_5184 ( .C ( clk ), .D ( signal_19876 ), .Q ( signal_19877 ) ) ;
    buf_clk cell_5188 ( .C ( clk ), .D ( signal_19880 ), .Q ( signal_19881 ) ) ;
    buf_clk cell_5192 ( .C ( clk ), .D ( signal_19884 ), .Q ( signal_19885 ) ) ;
    buf_clk cell_5246 ( .C ( clk ), .D ( signal_19938 ), .Q ( signal_19939 ) ) ;
    buf_clk cell_5250 ( .C ( clk ), .D ( signal_19942 ), .Q ( signal_19943 ) ) ;
    buf_clk cell_5254 ( .C ( clk ), .D ( signal_19946 ), .Q ( signal_19947 ) ) ;
    buf_clk cell_5258 ( .C ( clk ), .D ( signal_19950 ), .Q ( signal_19951 ) ) ;
    buf_clk cell_5262 ( .C ( clk ), .D ( signal_19954 ), .Q ( signal_19955 ) ) ;
    buf_clk cell_5298 ( .C ( clk ), .D ( signal_19990 ), .Q ( signal_19991 ) ) ;
    buf_clk cell_5304 ( .C ( clk ), .D ( signal_19996 ), .Q ( signal_19997 ) ) ;
    buf_clk cell_5310 ( .C ( clk ), .D ( signal_20002 ), .Q ( signal_20003 ) ) ;
    buf_clk cell_5316 ( .C ( clk ), .D ( signal_20008 ), .Q ( signal_20009 ) ) ;
    buf_clk cell_5322 ( .C ( clk ), .D ( signal_20014 ), .Q ( signal_20015 ) ) ;
    buf_clk cell_5336 ( .C ( clk ), .D ( signal_20028 ), .Q ( signal_20029 ) ) ;
    buf_clk cell_5340 ( .C ( clk ), .D ( signal_20032 ), .Q ( signal_20033 ) ) ;
    buf_clk cell_5344 ( .C ( clk ), .D ( signal_20036 ), .Q ( signal_20037 ) ) ;
    buf_clk cell_5348 ( .C ( clk ), .D ( signal_20040 ), .Q ( signal_20041 ) ) ;
    buf_clk cell_5352 ( .C ( clk ), .D ( signal_20044 ), .Q ( signal_20045 ) ) ;
    buf_clk cell_5378 ( .C ( clk ), .D ( signal_20070 ), .Q ( signal_20071 ) ) ;
    buf_clk cell_5384 ( .C ( clk ), .D ( signal_20076 ), .Q ( signal_20077 ) ) ;
    buf_clk cell_5390 ( .C ( clk ), .D ( signal_20082 ), .Q ( signal_20083 ) ) ;
    buf_clk cell_5396 ( .C ( clk ), .D ( signal_20088 ), .Q ( signal_20089 ) ) ;
    buf_clk cell_5402 ( .C ( clk ), .D ( signal_20094 ), .Q ( signal_20095 ) ) ;
    buf_clk cell_5406 ( .C ( clk ), .D ( signal_20098 ), .Q ( signal_20099 ) ) ;
    buf_clk cell_5410 ( .C ( clk ), .D ( signal_20102 ), .Q ( signal_20103 ) ) ;
    buf_clk cell_5414 ( .C ( clk ), .D ( signal_20106 ), .Q ( signal_20107 ) ) ;
    buf_clk cell_5418 ( .C ( clk ), .D ( signal_20110 ), .Q ( signal_20111 ) ) ;
    buf_clk cell_5422 ( .C ( clk ), .D ( signal_20114 ), .Q ( signal_20115 ) ) ;
    buf_clk cell_5446 ( .C ( clk ), .D ( signal_20138 ), .Q ( signal_20139 ) ) ;
    buf_clk cell_5450 ( .C ( clk ), .D ( signal_20142 ), .Q ( signal_20143 ) ) ;
    buf_clk cell_5454 ( .C ( clk ), .D ( signal_20146 ), .Q ( signal_20147 ) ) ;
    buf_clk cell_5458 ( .C ( clk ), .D ( signal_20150 ), .Q ( signal_20151 ) ) ;
    buf_clk cell_5462 ( .C ( clk ), .D ( signal_20154 ), .Q ( signal_20155 ) ) ;
    buf_clk cell_5466 ( .C ( clk ), .D ( signal_20158 ), .Q ( signal_20159 ) ) ;
    buf_clk cell_5470 ( .C ( clk ), .D ( signal_20162 ), .Q ( signal_20163 ) ) ;
    buf_clk cell_5474 ( .C ( clk ), .D ( signal_20166 ), .Q ( signal_20167 ) ) ;
    buf_clk cell_5478 ( .C ( clk ), .D ( signal_20170 ), .Q ( signal_20171 ) ) ;
    buf_clk cell_5482 ( .C ( clk ), .D ( signal_20174 ), .Q ( signal_20175 ) ) ;
    buf_clk cell_5486 ( .C ( clk ), .D ( signal_20178 ), .Q ( signal_20179 ) ) ;
    buf_clk cell_5490 ( .C ( clk ), .D ( signal_20182 ), .Q ( signal_20183 ) ) ;
    buf_clk cell_5494 ( .C ( clk ), .D ( signal_20186 ), .Q ( signal_20187 ) ) ;
    buf_clk cell_5498 ( .C ( clk ), .D ( signal_20190 ), .Q ( signal_20191 ) ) ;
    buf_clk cell_5502 ( .C ( clk ), .D ( signal_20194 ), .Q ( signal_20195 ) ) ;
    buf_clk cell_5518 ( .C ( clk ), .D ( signal_20210 ), .Q ( signal_20211 ) ) ;
    buf_clk cell_5524 ( .C ( clk ), .D ( signal_20216 ), .Q ( signal_20217 ) ) ;
    buf_clk cell_5530 ( .C ( clk ), .D ( signal_20222 ), .Q ( signal_20223 ) ) ;
    buf_clk cell_5536 ( .C ( clk ), .D ( signal_20228 ), .Q ( signal_20229 ) ) ;
    buf_clk cell_5542 ( .C ( clk ), .D ( signal_20234 ), .Q ( signal_20235 ) ) ;
    buf_clk cell_5546 ( .C ( clk ), .D ( signal_20238 ), .Q ( signal_20239 ) ) ;
    buf_clk cell_5550 ( .C ( clk ), .D ( signal_20242 ), .Q ( signal_20243 ) ) ;
    buf_clk cell_5554 ( .C ( clk ), .D ( signal_20246 ), .Q ( signal_20247 ) ) ;
    buf_clk cell_5558 ( .C ( clk ), .D ( signal_20250 ), .Q ( signal_20251 ) ) ;
    buf_clk cell_5562 ( .C ( clk ), .D ( signal_20254 ), .Q ( signal_20255 ) ) ;
    buf_clk cell_5568 ( .C ( clk ), .D ( signal_20260 ), .Q ( signal_20261 ) ) ;
    buf_clk cell_5574 ( .C ( clk ), .D ( signal_20266 ), .Q ( signal_20267 ) ) ;
    buf_clk cell_5580 ( .C ( clk ), .D ( signal_20272 ), .Q ( signal_20273 ) ) ;
    buf_clk cell_5586 ( .C ( clk ), .D ( signal_20278 ), .Q ( signal_20279 ) ) ;
    buf_clk cell_5592 ( .C ( clk ), .D ( signal_20284 ), .Q ( signal_20285 ) ) ;
    buf_clk cell_5596 ( .C ( clk ), .D ( signal_20288 ), .Q ( signal_20289 ) ) ;
    buf_clk cell_5600 ( .C ( clk ), .D ( signal_20292 ), .Q ( signal_20293 ) ) ;
    buf_clk cell_5604 ( .C ( clk ), .D ( signal_20296 ), .Q ( signal_20297 ) ) ;
    buf_clk cell_5608 ( .C ( clk ), .D ( signal_20300 ), .Q ( signal_20301 ) ) ;
    buf_clk cell_5612 ( .C ( clk ), .D ( signal_20304 ), .Q ( signal_20305 ) ) ;
    buf_clk cell_5616 ( .C ( clk ), .D ( signal_20308 ), .Q ( signal_20309 ) ) ;
    buf_clk cell_5620 ( .C ( clk ), .D ( signal_20312 ), .Q ( signal_20313 ) ) ;
    buf_clk cell_5624 ( .C ( clk ), .D ( signal_20316 ), .Q ( signal_20317 ) ) ;
    buf_clk cell_5628 ( .C ( clk ), .D ( signal_20320 ), .Q ( signal_20321 ) ) ;
    buf_clk cell_5632 ( .C ( clk ), .D ( signal_20324 ), .Q ( signal_20325 ) ) ;
    buf_clk cell_5636 ( .C ( clk ), .D ( signal_20328 ), .Q ( signal_20329 ) ) ;
    buf_clk cell_5640 ( .C ( clk ), .D ( signal_20332 ), .Q ( signal_20333 ) ) ;
    buf_clk cell_5644 ( .C ( clk ), .D ( signal_20336 ), .Q ( signal_20337 ) ) ;
    buf_clk cell_5648 ( .C ( clk ), .D ( signal_20340 ), .Q ( signal_20341 ) ) ;
    buf_clk cell_5652 ( .C ( clk ), .D ( signal_20344 ), .Q ( signal_20345 ) ) ;
    buf_clk cell_5666 ( .C ( clk ), .D ( signal_20358 ), .Q ( signal_20359 ) ) ;
    buf_clk cell_5670 ( .C ( clk ), .D ( signal_20362 ), .Q ( signal_20363 ) ) ;
    buf_clk cell_5674 ( .C ( clk ), .D ( signal_20366 ), .Q ( signal_20367 ) ) ;
    buf_clk cell_5678 ( .C ( clk ), .D ( signal_20370 ), .Q ( signal_20371 ) ) ;
    buf_clk cell_5682 ( .C ( clk ), .D ( signal_20374 ), .Q ( signal_20375 ) ) ;
    buf_clk cell_5686 ( .C ( clk ), .D ( signal_20378 ), .Q ( signal_20379 ) ) ;
    buf_clk cell_5690 ( .C ( clk ), .D ( signal_20382 ), .Q ( signal_20383 ) ) ;
    buf_clk cell_5694 ( .C ( clk ), .D ( signal_20386 ), .Q ( signal_20387 ) ) ;
    buf_clk cell_5698 ( .C ( clk ), .D ( signal_20390 ), .Q ( signal_20391 ) ) ;
    buf_clk cell_5702 ( .C ( clk ), .D ( signal_20394 ), .Q ( signal_20395 ) ) ;
    buf_clk cell_5708 ( .C ( clk ), .D ( signal_20400 ), .Q ( signal_20401 ) ) ;
    buf_clk cell_5714 ( .C ( clk ), .D ( signal_20406 ), .Q ( signal_20407 ) ) ;
    buf_clk cell_5720 ( .C ( clk ), .D ( signal_20412 ), .Q ( signal_20413 ) ) ;
    buf_clk cell_5726 ( .C ( clk ), .D ( signal_20418 ), .Q ( signal_20419 ) ) ;
    buf_clk cell_5732 ( .C ( clk ), .D ( signal_20424 ), .Q ( signal_20425 ) ) ;
    buf_clk cell_5756 ( .C ( clk ), .D ( signal_20448 ), .Q ( signal_20449 ) ) ;
    buf_clk cell_5760 ( .C ( clk ), .D ( signal_20452 ), .Q ( signal_20453 ) ) ;
    buf_clk cell_5764 ( .C ( clk ), .D ( signal_20456 ), .Q ( signal_20457 ) ) ;
    buf_clk cell_5768 ( .C ( clk ), .D ( signal_20460 ), .Q ( signal_20461 ) ) ;
    buf_clk cell_5772 ( .C ( clk ), .D ( signal_20464 ), .Q ( signal_20465 ) ) ;
    buf_clk cell_5778 ( .C ( clk ), .D ( signal_20470 ), .Q ( signal_20471 ) ) ;
    buf_clk cell_5784 ( .C ( clk ), .D ( signal_20476 ), .Q ( signal_20477 ) ) ;
    buf_clk cell_5790 ( .C ( clk ), .D ( signal_20482 ), .Q ( signal_20483 ) ) ;
    buf_clk cell_5796 ( .C ( clk ), .D ( signal_20488 ), .Q ( signal_20489 ) ) ;
    buf_clk cell_5802 ( .C ( clk ), .D ( signal_20494 ), .Q ( signal_20495 ) ) ;
    buf_clk cell_5808 ( .C ( clk ), .D ( signal_20500 ), .Q ( signal_20501 ) ) ;
    buf_clk cell_5814 ( .C ( clk ), .D ( signal_20506 ), .Q ( signal_20507 ) ) ;
    buf_clk cell_5820 ( .C ( clk ), .D ( signal_20512 ), .Q ( signal_20513 ) ) ;
    buf_clk cell_5826 ( .C ( clk ), .D ( signal_20518 ), .Q ( signal_20519 ) ) ;
    buf_clk cell_5832 ( .C ( clk ), .D ( signal_20524 ), .Q ( signal_20525 ) ) ;
    buf_clk cell_5838 ( .C ( clk ), .D ( signal_20530 ), .Q ( signal_20531 ) ) ;
    buf_clk cell_5844 ( .C ( clk ), .D ( signal_20536 ), .Q ( signal_20537 ) ) ;
    buf_clk cell_5850 ( .C ( clk ), .D ( signal_20542 ), .Q ( signal_20543 ) ) ;
    buf_clk cell_5856 ( .C ( clk ), .D ( signal_20548 ), .Q ( signal_20549 ) ) ;
    buf_clk cell_5862 ( .C ( clk ), .D ( signal_20554 ), .Q ( signal_20555 ) ) ;
    buf_clk cell_5866 ( .C ( clk ), .D ( signal_20558 ), .Q ( signal_20559 ) ) ;
    buf_clk cell_5870 ( .C ( clk ), .D ( signal_20562 ), .Q ( signal_20563 ) ) ;
    buf_clk cell_5874 ( .C ( clk ), .D ( signal_20566 ), .Q ( signal_20567 ) ) ;
    buf_clk cell_5878 ( .C ( clk ), .D ( signal_20570 ), .Q ( signal_20571 ) ) ;
    buf_clk cell_5882 ( .C ( clk ), .D ( signal_20574 ), .Q ( signal_20575 ) ) ;
    buf_clk cell_5908 ( .C ( clk ), .D ( signal_20600 ), .Q ( signal_20601 ) ) ;
    buf_clk cell_5916 ( .C ( clk ), .D ( signal_20608 ), .Q ( signal_20609 ) ) ;
    buf_clk cell_5924 ( .C ( clk ), .D ( signal_20616 ), .Q ( signal_20617 ) ) ;
    buf_clk cell_5932 ( .C ( clk ), .D ( signal_20624 ), .Q ( signal_20625 ) ) ;
    buf_clk cell_5940 ( .C ( clk ), .D ( signal_20632 ), .Q ( signal_20633 ) ) ;
    buf_clk cell_5966 ( .C ( clk ), .D ( signal_20658 ), .Q ( signal_20659 ) ) ;
    buf_clk cell_5972 ( .C ( clk ), .D ( signal_20664 ), .Q ( signal_20665 ) ) ;
    buf_clk cell_5978 ( .C ( clk ), .D ( signal_20670 ), .Q ( signal_20671 ) ) ;
    buf_clk cell_5984 ( .C ( clk ), .D ( signal_20676 ), .Q ( signal_20677 ) ) ;
    buf_clk cell_5990 ( .C ( clk ), .D ( signal_20682 ), .Q ( signal_20683 ) ) ;
    buf_clk cell_5996 ( .C ( clk ), .D ( signal_20688 ), .Q ( signal_20689 ) ) ;
    buf_clk cell_6002 ( .C ( clk ), .D ( signal_20694 ), .Q ( signal_20695 ) ) ;
    buf_clk cell_6008 ( .C ( clk ), .D ( signal_20700 ), .Q ( signal_20701 ) ) ;
    buf_clk cell_6014 ( .C ( clk ), .D ( signal_20706 ), .Q ( signal_20707 ) ) ;
    buf_clk cell_6020 ( .C ( clk ), .D ( signal_20712 ), .Q ( signal_20713 ) ) ;
    buf_clk cell_6046 ( .C ( clk ), .D ( signal_20738 ), .Q ( signal_20739 ) ) ;
    buf_clk cell_6052 ( .C ( clk ), .D ( signal_20744 ), .Q ( signal_20745 ) ) ;
    buf_clk cell_6058 ( .C ( clk ), .D ( signal_20750 ), .Q ( signal_20751 ) ) ;
    buf_clk cell_6064 ( .C ( clk ), .D ( signal_20756 ), .Q ( signal_20757 ) ) ;
    buf_clk cell_6070 ( .C ( clk ), .D ( signal_20762 ), .Q ( signal_20763 ) ) ;
    buf_clk cell_6136 ( .C ( clk ), .D ( signal_20828 ), .Q ( signal_20829 ) ) ;
    buf_clk cell_6142 ( .C ( clk ), .D ( signal_20834 ), .Q ( signal_20835 ) ) ;
    buf_clk cell_6148 ( .C ( clk ), .D ( signal_20840 ), .Q ( signal_20841 ) ) ;
    buf_clk cell_6154 ( .C ( clk ), .D ( signal_20846 ), .Q ( signal_20847 ) ) ;
    buf_clk cell_6160 ( .C ( clk ), .D ( signal_20852 ), .Q ( signal_20853 ) ) ;
    buf_clk cell_6166 ( .C ( clk ), .D ( signal_20858 ), .Q ( signal_20859 ) ) ;
    buf_clk cell_6172 ( .C ( clk ), .D ( signal_20864 ), .Q ( signal_20865 ) ) ;
    buf_clk cell_6178 ( .C ( clk ), .D ( signal_20870 ), .Q ( signal_20871 ) ) ;
    buf_clk cell_6184 ( .C ( clk ), .D ( signal_20876 ), .Q ( signal_20877 ) ) ;
    buf_clk cell_6190 ( .C ( clk ), .D ( signal_20882 ), .Q ( signal_20883 ) ) ;
    buf_clk cell_6196 ( .C ( clk ), .D ( signal_20888 ), .Q ( signal_20889 ) ) ;
    buf_clk cell_6202 ( .C ( clk ), .D ( signal_20894 ), .Q ( signal_20895 ) ) ;
    buf_clk cell_6208 ( .C ( clk ), .D ( signal_20900 ), .Q ( signal_20901 ) ) ;
    buf_clk cell_6214 ( .C ( clk ), .D ( signal_20906 ), .Q ( signal_20907 ) ) ;
    buf_clk cell_6220 ( .C ( clk ), .D ( signal_20912 ), .Q ( signal_20913 ) ) ;
    buf_clk cell_6256 ( .C ( clk ), .D ( signal_20948 ), .Q ( signal_20949 ) ) ;
    buf_clk cell_6262 ( .C ( clk ), .D ( signal_20954 ), .Q ( signal_20955 ) ) ;
    buf_clk cell_6268 ( .C ( clk ), .D ( signal_20960 ), .Q ( signal_20961 ) ) ;
    buf_clk cell_6274 ( .C ( clk ), .D ( signal_20966 ), .Q ( signal_20967 ) ) ;
    buf_clk cell_6280 ( .C ( clk ), .D ( signal_20972 ), .Q ( signal_20973 ) ) ;
    buf_clk cell_6296 ( .C ( clk ), .D ( signal_20988 ), .Q ( signal_20989 ) ) ;
    buf_clk cell_6302 ( .C ( clk ), .D ( signal_20994 ), .Q ( signal_20995 ) ) ;
    buf_clk cell_6308 ( .C ( clk ), .D ( signal_21000 ), .Q ( signal_21001 ) ) ;
    buf_clk cell_6314 ( .C ( clk ), .D ( signal_21006 ), .Q ( signal_21007 ) ) ;
    buf_clk cell_6320 ( .C ( clk ), .D ( signal_21012 ), .Q ( signal_21013 ) ) ;
    buf_clk cell_6338 ( .C ( clk ), .D ( signal_21030 ), .Q ( signal_21031 ) ) ;
    buf_clk cell_6346 ( .C ( clk ), .D ( signal_21038 ), .Q ( signal_21039 ) ) ;
    buf_clk cell_6354 ( .C ( clk ), .D ( signal_21046 ), .Q ( signal_21047 ) ) ;
    buf_clk cell_6362 ( .C ( clk ), .D ( signal_21054 ), .Q ( signal_21055 ) ) ;
    buf_clk cell_6370 ( .C ( clk ), .D ( signal_21062 ), .Q ( signal_21063 ) ) ;
    buf_clk cell_6416 ( .C ( clk ), .D ( signal_21108 ), .Q ( signal_21109 ) ) ;
    buf_clk cell_6422 ( .C ( clk ), .D ( signal_21114 ), .Q ( signal_21115 ) ) ;
    buf_clk cell_6428 ( .C ( clk ), .D ( signal_21120 ), .Q ( signal_21121 ) ) ;
    buf_clk cell_6434 ( .C ( clk ), .D ( signal_21126 ), .Q ( signal_21127 ) ) ;
    buf_clk cell_6440 ( .C ( clk ), .D ( signal_21132 ), .Q ( signal_21133 ) ) ;
    buf_clk cell_6446 ( .C ( clk ), .D ( signal_21138 ), .Q ( signal_21139 ) ) ;
    buf_clk cell_6452 ( .C ( clk ), .D ( signal_21144 ), .Q ( signal_21145 ) ) ;
    buf_clk cell_6458 ( .C ( clk ), .D ( signal_21150 ), .Q ( signal_21151 ) ) ;
    buf_clk cell_6464 ( .C ( clk ), .D ( signal_21156 ), .Q ( signal_21157 ) ) ;
    buf_clk cell_6470 ( .C ( clk ), .D ( signal_21162 ), .Q ( signal_21163 ) ) ;
    buf_clk cell_6498 ( .C ( clk ), .D ( signal_21190 ), .Q ( signal_21191 ) ) ;
    buf_clk cell_6506 ( .C ( clk ), .D ( signal_21198 ), .Q ( signal_21199 ) ) ;
    buf_clk cell_6514 ( .C ( clk ), .D ( signal_21206 ), .Q ( signal_21207 ) ) ;
    buf_clk cell_6522 ( .C ( clk ), .D ( signal_21214 ), .Q ( signal_21215 ) ) ;
    buf_clk cell_6530 ( .C ( clk ), .D ( signal_21222 ), .Q ( signal_21223 ) ) ;
    buf_clk cell_6536 ( .C ( clk ), .D ( signal_21228 ), .Q ( signal_21229 ) ) ;
    buf_clk cell_6542 ( .C ( clk ), .D ( signal_21234 ), .Q ( signal_21235 ) ) ;
    buf_clk cell_6548 ( .C ( clk ), .D ( signal_21240 ), .Q ( signal_21241 ) ) ;
    buf_clk cell_6554 ( .C ( clk ), .D ( signal_21246 ), .Q ( signal_21247 ) ) ;
    buf_clk cell_6560 ( .C ( clk ), .D ( signal_21252 ), .Q ( signal_21253 ) ) ;
    buf_clk cell_6566 ( .C ( clk ), .D ( signal_21258 ), .Q ( signal_21259 ) ) ;
    buf_clk cell_6572 ( .C ( clk ), .D ( signal_21264 ), .Q ( signal_21265 ) ) ;
    buf_clk cell_6578 ( .C ( clk ), .D ( signal_21270 ), .Q ( signal_21271 ) ) ;
    buf_clk cell_6584 ( .C ( clk ), .D ( signal_21276 ), .Q ( signal_21277 ) ) ;
    buf_clk cell_6590 ( .C ( clk ), .D ( signal_21282 ), .Q ( signal_21283 ) ) ;
    buf_clk cell_6616 ( .C ( clk ), .D ( signal_21308 ), .Q ( signal_21309 ) ) ;
    buf_clk cell_6622 ( .C ( clk ), .D ( signal_21314 ), .Q ( signal_21315 ) ) ;
    buf_clk cell_6628 ( .C ( clk ), .D ( signal_21320 ), .Q ( signal_21321 ) ) ;
    buf_clk cell_6634 ( .C ( clk ), .D ( signal_21326 ), .Q ( signal_21327 ) ) ;
    buf_clk cell_6640 ( .C ( clk ), .D ( signal_21332 ), .Q ( signal_21333 ) ) ;
    buf_clk cell_6666 ( .C ( clk ), .D ( signal_21358 ), .Q ( signal_21359 ) ) ;
    buf_clk cell_6672 ( .C ( clk ), .D ( signal_21364 ), .Q ( signal_21365 ) ) ;
    buf_clk cell_6678 ( .C ( clk ), .D ( signal_21370 ), .Q ( signal_21371 ) ) ;
    buf_clk cell_6684 ( .C ( clk ), .D ( signal_21376 ), .Q ( signal_21377 ) ) ;
    buf_clk cell_6690 ( .C ( clk ), .D ( signal_21382 ), .Q ( signal_21383 ) ) ;
    buf_clk cell_6696 ( .C ( clk ), .D ( signal_21388 ), .Q ( signal_21389 ) ) ;
    buf_clk cell_6702 ( .C ( clk ), .D ( signal_21394 ), .Q ( signal_21395 ) ) ;
    buf_clk cell_6708 ( .C ( clk ), .D ( signal_21400 ), .Q ( signal_21401 ) ) ;
    buf_clk cell_6714 ( .C ( clk ), .D ( signal_21406 ), .Q ( signal_21407 ) ) ;
    buf_clk cell_6720 ( .C ( clk ), .D ( signal_21412 ), .Q ( signal_21413 ) ) ;
    buf_clk cell_6748 ( .C ( clk ), .D ( signal_21440 ), .Q ( signal_21441 ) ) ;
    buf_clk cell_6758 ( .C ( clk ), .D ( signal_21450 ), .Q ( signal_21451 ) ) ;
    buf_clk cell_6768 ( .C ( clk ), .D ( signal_21460 ), .Q ( signal_21461 ) ) ;
    buf_clk cell_6778 ( .C ( clk ), .D ( signal_21470 ), .Q ( signal_21471 ) ) ;
    buf_clk cell_6788 ( .C ( clk ), .D ( signal_21480 ), .Q ( signal_21481 ) ) ;
    buf_clk cell_6826 ( .C ( clk ), .D ( signal_21518 ), .Q ( signal_21519 ) ) ;
    buf_clk cell_6834 ( .C ( clk ), .D ( signal_21526 ), .Q ( signal_21527 ) ) ;
    buf_clk cell_6842 ( .C ( clk ), .D ( signal_21534 ), .Q ( signal_21535 ) ) ;
    buf_clk cell_6850 ( .C ( clk ), .D ( signal_21542 ), .Q ( signal_21543 ) ) ;
    buf_clk cell_6858 ( .C ( clk ), .D ( signal_21550 ), .Q ( signal_21551 ) ) ;
    buf_clk cell_6866 ( .C ( clk ), .D ( signal_21558 ), .Q ( signal_21559 ) ) ;
    buf_clk cell_6874 ( .C ( clk ), .D ( signal_21566 ), .Q ( signal_21567 ) ) ;
    buf_clk cell_6882 ( .C ( clk ), .D ( signal_21574 ), .Q ( signal_21575 ) ) ;
    buf_clk cell_6890 ( .C ( clk ), .D ( signal_21582 ), .Q ( signal_21583 ) ) ;
    buf_clk cell_6898 ( .C ( clk ), .D ( signal_21590 ), .Q ( signal_21591 ) ) ;
    buf_clk cell_6988 ( .C ( clk ), .D ( signal_21680 ), .Q ( signal_21681 ) ) ;
    buf_clk cell_6998 ( .C ( clk ), .D ( signal_21690 ), .Q ( signal_21691 ) ) ;
    buf_clk cell_7008 ( .C ( clk ), .D ( signal_21700 ), .Q ( signal_21701 ) ) ;
    buf_clk cell_7018 ( .C ( clk ), .D ( signal_21710 ), .Q ( signal_21711 ) ) ;
    buf_clk cell_7028 ( .C ( clk ), .D ( signal_21720 ), .Q ( signal_21721 ) ) ;
    buf_clk cell_7076 ( .C ( clk ), .D ( signal_21768 ), .Q ( signal_21769 ) ) ;
    buf_clk cell_7084 ( .C ( clk ), .D ( signal_21776 ), .Q ( signal_21777 ) ) ;
    buf_clk cell_7092 ( .C ( clk ), .D ( signal_21784 ), .Q ( signal_21785 ) ) ;
    buf_clk cell_7100 ( .C ( clk ), .D ( signal_21792 ), .Q ( signal_21793 ) ) ;
    buf_clk cell_7108 ( .C ( clk ), .D ( signal_21800 ), .Q ( signal_21801 ) ) ;
    buf_clk cell_7146 ( .C ( clk ), .D ( signal_21838 ), .Q ( signal_21839 ) ) ;
    buf_clk cell_7154 ( .C ( clk ), .D ( signal_21846 ), .Q ( signal_21847 ) ) ;
    buf_clk cell_7162 ( .C ( clk ), .D ( signal_21854 ), .Q ( signal_21855 ) ) ;
    buf_clk cell_7170 ( .C ( clk ), .D ( signal_21862 ), .Q ( signal_21863 ) ) ;
    buf_clk cell_7178 ( .C ( clk ), .D ( signal_21870 ), .Q ( signal_21871 ) ) ;
    buf_clk cell_7186 ( .C ( clk ), .D ( signal_21878 ), .Q ( signal_21879 ) ) ;
    buf_clk cell_7194 ( .C ( clk ), .D ( signal_21886 ), .Q ( signal_21887 ) ) ;
    buf_clk cell_7202 ( .C ( clk ), .D ( signal_21894 ), .Q ( signal_21895 ) ) ;
    buf_clk cell_7210 ( .C ( clk ), .D ( signal_21902 ), .Q ( signal_21903 ) ) ;
    buf_clk cell_7218 ( .C ( clk ), .D ( signal_21910 ), .Q ( signal_21911 ) ) ;
    buf_clk cell_7226 ( .C ( clk ), .D ( signal_21918 ), .Q ( signal_21919 ) ) ;
    buf_clk cell_7234 ( .C ( clk ), .D ( signal_21926 ), .Q ( signal_21927 ) ) ;
    buf_clk cell_7242 ( .C ( clk ), .D ( signal_21934 ), .Q ( signal_21935 ) ) ;
    buf_clk cell_7250 ( .C ( clk ), .D ( signal_21942 ), .Q ( signal_21943 ) ) ;
    buf_clk cell_7258 ( .C ( clk ), .D ( signal_21950 ), .Q ( signal_21951 ) ) ;
    buf_clk cell_7268 ( .C ( clk ), .D ( signal_21960 ), .Q ( signal_21961 ) ) ;
    buf_clk cell_7278 ( .C ( clk ), .D ( signal_21970 ), .Q ( signal_21971 ) ) ;
    buf_clk cell_7288 ( .C ( clk ), .D ( signal_21980 ), .Q ( signal_21981 ) ) ;
    buf_clk cell_7298 ( .C ( clk ), .D ( signal_21990 ), .Q ( signal_21991 ) ) ;
    buf_clk cell_7308 ( .C ( clk ), .D ( signal_22000 ), .Q ( signal_22001 ) ) ;
    buf_clk cell_7316 ( .C ( clk ), .D ( signal_22008 ), .Q ( signal_22009 ) ) ;
    buf_clk cell_7324 ( .C ( clk ), .D ( signal_22016 ), .Q ( signal_22017 ) ) ;
    buf_clk cell_7332 ( .C ( clk ), .D ( signal_22024 ), .Q ( signal_22025 ) ) ;
    buf_clk cell_7340 ( .C ( clk ), .D ( signal_22032 ), .Q ( signal_22033 ) ) ;
    buf_clk cell_7348 ( .C ( clk ), .D ( signal_22040 ), .Q ( signal_22041 ) ) ;
    buf_clk cell_7356 ( .C ( clk ), .D ( signal_22048 ), .Q ( signal_22049 ) ) ;
    buf_clk cell_7364 ( .C ( clk ), .D ( signal_22056 ), .Q ( signal_22057 ) ) ;
    buf_clk cell_7372 ( .C ( clk ), .D ( signal_22064 ), .Q ( signal_22065 ) ) ;
    buf_clk cell_7380 ( .C ( clk ), .D ( signal_22072 ), .Q ( signal_22073 ) ) ;
    buf_clk cell_7388 ( .C ( clk ), .D ( signal_22080 ), .Q ( signal_22081 ) ) ;
    buf_clk cell_7406 ( .C ( clk ), .D ( signal_22098 ), .Q ( signal_22099 ) ) ;
    buf_clk cell_7414 ( .C ( clk ), .D ( signal_22106 ), .Q ( signal_22107 ) ) ;
    buf_clk cell_7422 ( .C ( clk ), .D ( signal_22114 ), .Q ( signal_22115 ) ) ;
    buf_clk cell_7430 ( .C ( clk ), .D ( signal_22122 ), .Q ( signal_22123 ) ) ;
    buf_clk cell_7438 ( .C ( clk ), .D ( signal_22130 ), .Q ( signal_22131 ) ) ;
    buf_clk cell_7446 ( .C ( clk ), .D ( signal_22138 ), .Q ( signal_22139 ) ) ;
    buf_clk cell_7454 ( .C ( clk ), .D ( signal_22146 ), .Q ( signal_22147 ) ) ;
    buf_clk cell_7462 ( .C ( clk ), .D ( signal_22154 ), .Q ( signal_22155 ) ) ;
    buf_clk cell_7470 ( .C ( clk ), .D ( signal_22162 ), .Q ( signal_22163 ) ) ;
    buf_clk cell_7478 ( .C ( clk ), .D ( signal_22170 ), .Q ( signal_22171 ) ) ;
    buf_clk cell_7486 ( .C ( clk ), .D ( signal_22178 ), .Q ( signal_22179 ) ) ;
    buf_clk cell_7494 ( .C ( clk ), .D ( signal_22186 ), .Q ( signal_22187 ) ) ;
    buf_clk cell_7502 ( .C ( clk ), .D ( signal_22194 ), .Q ( signal_22195 ) ) ;
    buf_clk cell_7510 ( .C ( clk ), .D ( signal_22202 ), .Q ( signal_22203 ) ) ;
    buf_clk cell_7518 ( .C ( clk ), .D ( signal_22210 ), .Q ( signal_22211 ) ) ;
    buf_clk cell_7696 ( .C ( clk ), .D ( signal_22388 ), .Q ( signal_22389 ) ) ;
    buf_clk cell_7706 ( .C ( clk ), .D ( signal_22398 ), .Q ( signal_22399 ) ) ;
    buf_clk cell_7716 ( .C ( clk ), .D ( signal_22408 ), .Q ( signal_22409 ) ) ;
    buf_clk cell_7726 ( .C ( clk ), .D ( signal_22418 ), .Q ( signal_22419 ) ) ;
    buf_clk cell_7736 ( .C ( clk ), .D ( signal_22428 ), .Q ( signal_22429 ) ) ;
    buf_clk cell_7826 ( .C ( clk ), .D ( signal_22518 ), .Q ( signal_22519 ) ) ;
    buf_clk cell_7836 ( .C ( clk ), .D ( signal_22528 ), .Q ( signal_22529 ) ) ;
    buf_clk cell_7846 ( .C ( clk ), .D ( signal_22538 ), .Q ( signal_22539 ) ) ;
    buf_clk cell_7856 ( .C ( clk ), .D ( signal_22548 ), .Q ( signal_22549 ) ) ;
    buf_clk cell_7866 ( .C ( clk ), .D ( signal_22558 ), .Q ( signal_22559 ) ) ;
    buf_clk cell_8836 ( .C ( clk ), .D ( signal_23528 ), .Q ( signal_23529 ) ) ;
    buf_clk cell_8850 ( .C ( clk ), .D ( signal_23542 ), .Q ( signal_23543 ) ) ;
    buf_clk cell_8864 ( .C ( clk ), .D ( signal_23556 ), .Q ( signal_23557 ) ) ;
    buf_clk cell_8878 ( .C ( clk ), .D ( signal_23570 ), .Q ( signal_23571 ) ) ;
    buf_clk cell_8892 ( .C ( clk ), .D ( signal_23584 ), .Q ( signal_23585 ) ) ;
    buf_clk cell_8946 ( .C ( clk ), .D ( signal_23638 ), .Q ( signal_23639 ) ) ;
    buf_clk cell_8960 ( .C ( clk ), .D ( signal_23652 ), .Q ( signal_23653 ) ) ;
    buf_clk cell_8974 ( .C ( clk ), .D ( signal_23666 ), .Q ( signal_23667 ) ) ;
    buf_clk cell_8988 ( .C ( clk ), .D ( signal_23680 ), .Q ( signal_23681 ) ) ;
    buf_clk cell_9002 ( .C ( clk ), .D ( signal_23694 ), .Q ( signal_23695 ) ) ;
    buf_clk cell_9146 ( .C ( clk ), .D ( signal_23838 ), .Q ( signal_23839 ) ) ;
    buf_clk cell_9162 ( .C ( clk ), .D ( signal_23854 ), .Q ( signal_23855 ) ) ;
    buf_clk cell_9178 ( .C ( clk ), .D ( signal_23870 ), .Q ( signal_23871 ) ) ;
    buf_clk cell_9194 ( .C ( clk ), .D ( signal_23886 ), .Q ( signal_23887 ) ) ;
    buf_clk cell_9210 ( .C ( clk ), .D ( signal_23902 ), .Q ( signal_23903 ) ) ;
    buf_clk cell_9246 ( .C ( clk ), .D ( signal_23938 ), .Q ( signal_23939 ) ) ;
    buf_clk cell_9262 ( .C ( clk ), .D ( signal_23954 ), .Q ( signal_23955 ) ) ;
    buf_clk cell_9278 ( .C ( clk ), .D ( signal_23970 ), .Q ( signal_23971 ) ) ;
    buf_clk cell_9294 ( .C ( clk ), .D ( signal_23986 ), .Q ( signal_23987 ) ) ;
    buf_clk cell_9310 ( .C ( clk ), .D ( signal_24002 ), .Q ( signal_24003 ) ) ;
    buf_clk cell_9636 ( .C ( clk ), .D ( signal_24328 ), .Q ( signal_24329 ) ) ;
    buf_clk cell_9654 ( .C ( clk ), .D ( signal_24346 ), .Q ( signal_24347 ) ) ;
    buf_clk cell_9672 ( .C ( clk ), .D ( signal_24364 ), .Q ( signal_24365 ) ) ;
    buf_clk cell_9690 ( .C ( clk ), .D ( signal_24382 ), .Q ( signal_24383 ) ) ;
    buf_clk cell_9708 ( .C ( clk ), .D ( signal_24400 ), .Q ( signal_24401 ) ) ;
    buf_clk cell_9886 ( .C ( clk ), .D ( signal_24578 ), .Q ( signal_24579 ) ) ;
    buf_clk cell_9906 ( .C ( clk ), .D ( signal_24598 ), .Q ( signal_24599 ) ) ;
    buf_clk cell_9926 ( .C ( clk ), .D ( signal_24618 ), .Q ( signal_24619 ) ) ;
    buf_clk cell_9946 ( .C ( clk ), .D ( signal_24638 ), .Q ( signal_24639 ) ) ;
    buf_clk cell_9966 ( .C ( clk ), .D ( signal_24658 ), .Q ( signal_24659 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_4895 ( .C ( clk ), .D ( signal_19379 ), .Q ( signal_19588 ) ) ;
    buf_clk cell_4897 ( .C ( clk ), .D ( signal_19381 ), .Q ( signal_19590 ) ) ;
    buf_clk cell_4899 ( .C ( clk ), .D ( signal_19383 ), .Q ( signal_19592 ) ) ;
    buf_clk cell_4901 ( .C ( clk ), .D ( signal_19385 ), .Q ( signal_19594 ) ) ;
    buf_clk cell_4903 ( .C ( clk ), .D ( signal_19387 ), .Q ( signal_19596 ) ) ;
    buf_clk cell_4909 ( .C ( clk ), .D ( signal_19601 ), .Q ( signal_19602 ) ) ;
    buf_clk cell_4915 ( .C ( clk ), .D ( signal_19607 ), .Q ( signal_19608 ) ) ;
    buf_clk cell_4921 ( .C ( clk ), .D ( signal_19613 ), .Q ( signal_19614 ) ) ;
    buf_clk cell_4927 ( .C ( clk ), .D ( signal_19619 ), .Q ( signal_19620 ) ) ;
    buf_clk cell_4933 ( .C ( clk ), .D ( signal_19625 ), .Q ( signal_19626 ) ) ;
    buf_clk cell_4939 ( .C ( clk ), .D ( signal_19631 ), .Q ( signal_19632 ) ) ;
    buf_clk cell_4945 ( .C ( clk ), .D ( signal_19637 ), .Q ( signal_19638 ) ) ;
    buf_clk cell_4951 ( .C ( clk ), .D ( signal_19643 ), .Q ( signal_19644 ) ) ;
    buf_clk cell_4957 ( .C ( clk ), .D ( signal_19649 ), .Q ( signal_19650 ) ) ;
    buf_clk cell_4963 ( .C ( clk ), .D ( signal_19655 ), .Q ( signal_19656 ) ) ;
    buf_clk cell_4969 ( .C ( clk ), .D ( signal_19661 ), .Q ( signal_19662 ) ) ;
    buf_clk cell_4975 ( .C ( clk ), .D ( signal_19667 ), .Q ( signal_19668 ) ) ;
    buf_clk cell_4981 ( .C ( clk ), .D ( signal_19673 ), .Q ( signal_19674 ) ) ;
    buf_clk cell_4987 ( .C ( clk ), .D ( signal_19679 ), .Q ( signal_19680 ) ) ;
    buf_clk cell_4993 ( .C ( clk ), .D ( signal_19685 ), .Q ( signal_19686 ) ) ;
    buf_clk cell_4997 ( .C ( clk ), .D ( signal_19689 ), .Q ( signal_19690 ) ) ;
    buf_clk cell_5001 ( .C ( clk ), .D ( signal_19693 ), .Q ( signal_19694 ) ) ;
    buf_clk cell_5005 ( .C ( clk ), .D ( signal_19697 ), .Q ( signal_19698 ) ) ;
    buf_clk cell_5009 ( .C ( clk ), .D ( signal_19701 ), .Q ( signal_19702 ) ) ;
    buf_clk cell_5013 ( .C ( clk ), .D ( signal_19705 ), .Q ( signal_19706 ) ) ;
    buf_clk cell_5019 ( .C ( clk ), .D ( signal_19711 ), .Q ( signal_19712 ) ) ;
    buf_clk cell_5025 ( .C ( clk ), .D ( signal_19717 ), .Q ( signal_19718 ) ) ;
    buf_clk cell_5031 ( .C ( clk ), .D ( signal_19723 ), .Q ( signal_19724 ) ) ;
    buf_clk cell_5037 ( .C ( clk ), .D ( signal_19729 ), .Q ( signal_19730 ) ) ;
    buf_clk cell_5043 ( .C ( clk ), .D ( signal_19735 ), .Q ( signal_19736 ) ) ;
    buf_clk cell_5047 ( .C ( clk ), .D ( signal_19739 ), .Q ( signal_19740 ) ) ;
    buf_clk cell_5051 ( .C ( clk ), .D ( signal_19743 ), .Q ( signal_19744 ) ) ;
    buf_clk cell_5055 ( .C ( clk ), .D ( signal_19747 ), .Q ( signal_19748 ) ) ;
    buf_clk cell_5059 ( .C ( clk ), .D ( signal_19751 ), .Q ( signal_19752 ) ) ;
    buf_clk cell_5063 ( .C ( clk ), .D ( signal_19755 ), .Q ( signal_19756 ) ) ;
    buf_clk cell_5067 ( .C ( clk ), .D ( signal_19759 ), .Q ( signal_19760 ) ) ;
    buf_clk cell_5071 ( .C ( clk ), .D ( signal_19763 ), .Q ( signal_19764 ) ) ;
    buf_clk cell_5075 ( .C ( clk ), .D ( signal_19767 ), .Q ( signal_19768 ) ) ;
    buf_clk cell_5079 ( .C ( clk ), .D ( signal_19771 ), .Q ( signal_19772 ) ) ;
    buf_clk cell_5083 ( .C ( clk ), .D ( signal_19775 ), .Q ( signal_19776 ) ) ;
    buf_clk cell_5087 ( .C ( clk ), .D ( signal_19779 ), .Q ( signal_19780 ) ) ;
    buf_clk cell_5091 ( .C ( clk ), .D ( signal_19783 ), .Q ( signal_19784 ) ) ;
    buf_clk cell_5095 ( .C ( clk ), .D ( signal_19787 ), .Q ( signal_19788 ) ) ;
    buf_clk cell_5099 ( .C ( clk ), .D ( signal_19791 ), .Q ( signal_19792 ) ) ;
    buf_clk cell_5103 ( .C ( clk ), .D ( signal_19795 ), .Q ( signal_19796 ) ) ;
    buf_clk cell_5107 ( .C ( clk ), .D ( signal_19799 ), .Q ( signal_19800 ) ) ;
    buf_clk cell_5111 ( .C ( clk ), .D ( signal_19803 ), .Q ( signal_19804 ) ) ;
    buf_clk cell_5115 ( .C ( clk ), .D ( signal_19807 ), .Q ( signal_19808 ) ) ;
    buf_clk cell_5119 ( .C ( clk ), .D ( signal_19811 ), .Q ( signal_19812 ) ) ;
    buf_clk cell_5123 ( .C ( clk ), .D ( signal_19815 ), .Q ( signal_19816 ) ) ;
    buf_clk cell_5127 ( .C ( clk ), .D ( signal_19819 ), .Q ( signal_19820 ) ) ;
    buf_clk cell_5131 ( .C ( clk ), .D ( signal_19823 ), .Q ( signal_19824 ) ) ;
    buf_clk cell_5135 ( .C ( clk ), .D ( signal_19827 ), .Q ( signal_19828 ) ) ;
    buf_clk cell_5139 ( .C ( clk ), .D ( signal_19831 ), .Q ( signal_19832 ) ) ;
    buf_clk cell_5143 ( .C ( clk ), .D ( signal_19835 ), .Q ( signal_19836 ) ) ;
    buf_clk cell_5149 ( .C ( clk ), .D ( signal_19841 ), .Q ( signal_19842 ) ) ;
    buf_clk cell_5155 ( .C ( clk ), .D ( signal_19847 ), .Q ( signal_19848 ) ) ;
    buf_clk cell_5161 ( .C ( clk ), .D ( signal_19853 ), .Q ( signal_19854 ) ) ;
    buf_clk cell_5167 ( .C ( clk ), .D ( signal_19859 ), .Q ( signal_19860 ) ) ;
    buf_clk cell_5173 ( .C ( clk ), .D ( signal_19865 ), .Q ( signal_19866 ) ) ;
    buf_clk cell_5177 ( .C ( clk ), .D ( signal_19869 ), .Q ( signal_19870 ) ) ;
    buf_clk cell_5181 ( .C ( clk ), .D ( signal_19873 ), .Q ( signal_19874 ) ) ;
    buf_clk cell_5185 ( .C ( clk ), .D ( signal_19877 ), .Q ( signal_19878 ) ) ;
    buf_clk cell_5189 ( .C ( clk ), .D ( signal_19881 ), .Q ( signal_19882 ) ) ;
    buf_clk cell_5193 ( .C ( clk ), .D ( signal_19885 ), .Q ( signal_19886 ) ) ;
    buf_clk cell_5195 ( .C ( clk ), .D ( signal_1999 ), .Q ( signal_19888 ) ) ;
    buf_clk cell_5197 ( .C ( clk ), .D ( signal_6652 ), .Q ( signal_19890 ) ) ;
    buf_clk cell_5199 ( .C ( clk ), .D ( signal_6653 ), .Q ( signal_19892 ) ) ;
    buf_clk cell_5201 ( .C ( clk ), .D ( signal_6654 ), .Q ( signal_19894 ) ) ;
    buf_clk cell_5203 ( .C ( clk ), .D ( signal_6655 ), .Q ( signal_19896 ) ) ;
    buf_clk cell_5205 ( .C ( clk ), .D ( signal_19149 ), .Q ( signal_19898 ) ) ;
    buf_clk cell_5207 ( .C ( clk ), .D ( signal_19151 ), .Q ( signal_19900 ) ) ;
    buf_clk cell_5209 ( .C ( clk ), .D ( signal_19153 ), .Q ( signal_19902 ) ) ;
    buf_clk cell_5211 ( .C ( clk ), .D ( signal_19155 ), .Q ( signal_19904 ) ) ;
    buf_clk cell_5213 ( .C ( clk ), .D ( signal_19157 ), .Q ( signal_19906 ) ) ;
    buf_clk cell_5215 ( .C ( clk ), .D ( signal_1811 ), .Q ( signal_19908 ) ) ;
    buf_clk cell_5217 ( .C ( clk ), .D ( signal_5900 ), .Q ( signal_19910 ) ) ;
    buf_clk cell_5219 ( .C ( clk ), .D ( signal_5901 ), .Q ( signal_19912 ) ) ;
    buf_clk cell_5221 ( .C ( clk ), .D ( signal_5902 ), .Q ( signal_19914 ) ) ;
    buf_clk cell_5223 ( .C ( clk ), .D ( signal_5903 ), .Q ( signal_19916 ) ) ;
    buf_clk cell_5225 ( .C ( clk ), .D ( signal_1980 ), .Q ( signal_19918 ) ) ;
    buf_clk cell_5227 ( .C ( clk ), .D ( signal_6576 ), .Q ( signal_19920 ) ) ;
    buf_clk cell_5229 ( .C ( clk ), .D ( signal_6577 ), .Q ( signal_19922 ) ) ;
    buf_clk cell_5231 ( .C ( clk ), .D ( signal_6578 ), .Q ( signal_19924 ) ) ;
    buf_clk cell_5233 ( .C ( clk ), .D ( signal_6579 ), .Q ( signal_19926 ) ) ;
    buf_clk cell_5235 ( .C ( clk ), .D ( signal_1983 ), .Q ( signal_19928 ) ) ;
    buf_clk cell_5237 ( .C ( clk ), .D ( signal_6588 ), .Q ( signal_19930 ) ) ;
    buf_clk cell_5239 ( .C ( clk ), .D ( signal_6589 ), .Q ( signal_19932 ) ) ;
    buf_clk cell_5241 ( .C ( clk ), .D ( signal_6590 ), .Q ( signal_19934 ) ) ;
    buf_clk cell_5243 ( .C ( clk ), .D ( signal_6591 ), .Q ( signal_19936 ) ) ;
    buf_clk cell_5247 ( .C ( clk ), .D ( signal_19939 ), .Q ( signal_19940 ) ) ;
    buf_clk cell_5251 ( .C ( clk ), .D ( signal_19943 ), .Q ( signal_19944 ) ) ;
    buf_clk cell_5255 ( .C ( clk ), .D ( signal_19947 ), .Q ( signal_19948 ) ) ;
    buf_clk cell_5259 ( .C ( clk ), .D ( signal_19951 ), .Q ( signal_19952 ) ) ;
    buf_clk cell_5263 ( .C ( clk ), .D ( signal_19955 ), .Q ( signal_19956 ) ) ;
    buf_clk cell_5265 ( .C ( clk ), .D ( signal_1965 ), .Q ( signal_19958 ) ) ;
    buf_clk cell_5267 ( .C ( clk ), .D ( signal_6516 ), .Q ( signal_19960 ) ) ;
    buf_clk cell_5269 ( .C ( clk ), .D ( signal_6517 ), .Q ( signal_19962 ) ) ;
    buf_clk cell_5271 ( .C ( clk ), .D ( signal_6518 ), .Q ( signal_19964 ) ) ;
    buf_clk cell_5273 ( .C ( clk ), .D ( signal_6519 ), .Q ( signal_19966 ) ) ;
    buf_clk cell_5275 ( .C ( clk ), .D ( signal_1968 ), .Q ( signal_19968 ) ) ;
    buf_clk cell_5277 ( .C ( clk ), .D ( signal_6528 ), .Q ( signal_19970 ) ) ;
    buf_clk cell_5279 ( .C ( clk ), .D ( signal_6529 ), .Q ( signal_19972 ) ) ;
    buf_clk cell_5281 ( .C ( clk ), .D ( signal_6530 ), .Q ( signal_19974 ) ) ;
    buf_clk cell_5283 ( .C ( clk ), .D ( signal_6531 ), .Q ( signal_19976 ) ) ;
    buf_clk cell_5285 ( .C ( clk ), .D ( signal_19259 ), .Q ( signal_19978 ) ) ;
    buf_clk cell_5287 ( .C ( clk ), .D ( signal_19261 ), .Q ( signal_19980 ) ) ;
    buf_clk cell_5289 ( .C ( clk ), .D ( signal_19263 ), .Q ( signal_19982 ) ) ;
    buf_clk cell_5291 ( .C ( clk ), .D ( signal_19265 ), .Q ( signal_19984 ) ) ;
    buf_clk cell_5293 ( .C ( clk ), .D ( signal_19267 ), .Q ( signal_19986 ) ) ;
    buf_clk cell_5299 ( .C ( clk ), .D ( signal_19991 ), .Q ( signal_19992 ) ) ;
    buf_clk cell_5305 ( .C ( clk ), .D ( signal_19997 ), .Q ( signal_19998 ) ) ;
    buf_clk cell_5311 ( .C ( clk ), .D ( signal_20003 ), .Q ( signal_20004 ) ) ;
    buf_clk cell_5317 ( .C ( clk ), .D ( signal_20009 ), .Q ( signal_20010 ) ) ;
    buf_clk cell_5323 ( .C ( clk ), .D ( signal_20015 ), .Q ( signal_20016 ) ) ;
    buf_clk cell_5325 ( .C ( clk ), .D ( signal_1970 ), .Q ( signal_20018 ) ) ;
    buf_clk cell_5327 ( .C ( clk ), .D ( signal_6536 ), .Q ( signal_20020 ) ) ;
    buf_clk cell_5329 ( .C ( clk ), .D ( signal_6537 ), .Q ( signal_20022 ) ) ;
    buf_clk cell_5331 ( .C ( clk ), .D ( signal_6538 ), .Q ( signal_20024 ) ) ;
    buf_clk cell_5333 ( .C ( clk ), .D ( signal_6539 ), .Q ( signal_20026 ) ) ;
    buf_clk cell_5337 ( .C ( clk ), .D ( signal_20029 ), .Q ( signal_20030 ) ) ;
    buf_clk cell_5341 ( .C ( clk ), .D ( signal_20033 ), .Q ( signal_20034 ) ) ;
    buf_clk cell_5345 ( .C ( clk ), .D ( signal_20037 ), .Q ( signal_20038 ) ) ;
    buf_clk cell_5349 ( .C ( clk ), .D ( signal_20041 ), .Q ( signal_20042 ) ) ;
    buf_clk cell_5353 ( .C ( clk ), .D ( signal_20045 ), .Q ( signal_20046 ) ) ;
    buf_clk cell_5355 ( .C ( clk ), .D ( signal_19081 ), .Q ( signal_20048 ) ) ;
    buf_clk cell_5357 ( .C ( clk ), .D ( signal_19085 ), .Q ( signal_20050 ) ) ;
    buf_clk cell_5359 ( .C ( clk ), .D ( signal_19089 ), .Q ( signal_20052 ) ) ;
    buf_clk cell_5361 ( .C ( clk ), .D ( signal_19093 ), .Q ( signal_20054 ) ) ;
    buf_clk cell_5363 ( .C ( clk ), .D ( signal_19097 ), .Q ( signal_20056 ) ) ;
    buf_clk cell_5365 ( .C ( clk ), .D ( signal_19279 ), .Q ( signal_20058 ) ) ;
    buf_clk cell_5367 ( .C ( clk ), .D ( signal_19281 ), .Q ( signal_20060 ) ) ;
    buf_clk cell_5369 ( .C ( clk ), .D ( signal_19283 ), .Q ( signal_20062 ) ) ;
    buf_clk cell_5371 ( .C ( clk ), .D ( signal_19285 ), .Q ( signal_20064 ) ) ;
    buf_clk cell_5373 ( .C ( clk ), .D ( signal_19287 ), .Q ( signal_20066 ) ) ;
    buf_clk cell_5379 ( .C ( clk ), .D ( signal_20071 ), .Q ( signal_20072 ) ) ;
    buf_clk cell_5385 ( .C ( clk ), .D ( signal_20077 ), .Q ( signal_20078 ) ) ;
    buf_clk cell_5391 ( .C ( clk ), .D ( signal_20083 ), .Q ( signal_20084 ) ) ;
    buf_clk cell_5397 ( .C ( clk ), .D ( signal_20089 ), .Q ( signal_20090 ) ) ;
    buf_clk cell_5403 ( .C ( clk ), .D ( signal_20095 ), .Q ( signal_20096 ) ) ;
    buf_clk cell_5407 ( .C ( clk ), .D ( signal_20099 ), .Q ( signal_20100 ) ) ;
    buf_clk cell_5411 ( .C ( clk ), .D ( signal_20103 ), .Q ( signal_20104 ) ) ;
    buf_clk cell_5415 ( .C ( clk ), .D ( signal_20107 ), .Q ( signal_20108 ) ) ;
    buf_clk cell_5419 ( .C ( clk ), .D ( signal_20111 ), .Q ( signal_20112 ) ) ;
    buf_clk cell_5423 ( .C ( clk ), .D ( signal_20115 ), .Q ( signal_20116 ) ) ;
    buf_clk cell_5425 ( .C ( clk ), .D ( signal_1755 ), .Q ( signal_20118 ) ) ;
    buf_clk cell_5427 ( .C ( clk ), .D ( signal_5676 ), .Q ( signal_20120 ) ) ;
    buf_clk cell_5429 ( .C ( clk ), .D ( signal_5677 ), .Q ( signal_20122 ) ) ;
    buf_clk cell_5431 ( .C ( clk ), .D ( signal_5678 ), .Q ( signal_20124 ) ) ;
    buf_clk cell_5433 ( .C ( clk ), .D ( signal_5679 ), .Q ( signal_20126 ) ) ;
    buf_clk cell_5435 ( .C ( clk ), .D ( signal_1987 ), .Q ( signal_20128 ) ) ;
    buf_clk cell_5437 ( .C ( clk ), .D ( signal_6604 ), .Q ( signal_20130 ) ) ;
    buf_clk cell_5439 ( .C ( clk ), .D ( signal_6605 ), .Q ( signal_20132 ) ) ;
    buf_clk cell_5441 ( .C ( clk ), .D ( signal_6606 ), .Q ( signal_20134 ) ) ;
    buf_clk cell_5443 ( .C ( clk ), .D ( signal_6607 ), .Q ( signal_20136 ) ) ;
    buf_clk cell_5447 ( .C ( clk ), .D ( signal_20139 ), .Q ( signal_20140 ) ) ;
    buf_clk cell_5451 ( .C ( clk ), .D ( signal_20143 ), .Q ( signal_20144 ) ) ;
    buf_clk cell_5455 ( .C ( clk ), .D ( signal_20147 ), .Q ( signal_20148 ) ) ;
    buf_clk cell_5459 ( .C ( clk ), .D ( signal_20151 ), .Q ( signal_20152 ) ) ;
    buf_clk cell_5463 ( .C ( clk ), .D ( signal_20155 ), .Q ( signal_20156 ) ) ;
    buf_clk cell_5467 ( .C ( clk ), .D ( signal_20159 ), .Q ( signal_20160 ) ) ;
    buf_clk cell_5471 ( .C ( clk ), .D ( signal_20163 ), .Q ( signal_20164 ) ) ;
    buf_clk cell_5475 ( .C ( clk ), .D ( signal_20167 ), .Q ( signal_20168 ) ) ;
    buf_clk cell_5479 ( .C ( clk ), .D ( signal_20171 ), .Q ( signal_20172 ) ) ;
    buf_clk cell_5483 ( .C ( clk ), .D ( signal_20175 ), .Q ( signal_20176 ) ) ;
    buf_clk cell_5487 ( .C ( clk ), .D ( signal_20179 ), .Q ( signal_20180 ) ) ;
    buf_clk cell_5491 ( .C ( clk ), .D ( signal_20183 ), .Q ( signal_20184 ) ) ;
    buf_clk cell_5495 ( .C ( clk ), .D ( signal_20187 ), .Q ( signal_20188 ) ) ;
    buf_clk cell_5499 ( .C ( clk ), .D ( signal_20191 ), .Q ( signal_20192 ) ) ;
    buf_clk cell_5503 ( .C ( clk ), .D ( signal_20195 ), .Q ( signal_20196 ) ) ;
    buf_clk cell_5505 ( .C ( clk ), .D ( signal_19211 ), .Q ( signal_20198 ) ) ;
    buf_clk cell_5507 ( .C ( clk ), .D ( signal_19215 ), .Q ( signal_20200 ) ) ;
    buf_clk cell_5509 ( .C ( clk ), .D ( signal_19219 ), .Q ( signal_20202 ) ) ;
    buf_clk cell_5511 ( .C ( clk ), .D ( signal_19223 ), .Q ( signal_20204 ) ) ;
    buf_clk cell_5513 ( .C ( clk ), .D ( signal_19227 ), .Q ( signal_20206 ) ) ;
    buf_clk cell_5519 ( .C ( clk ), .D ( signal_20211 ), .Q ( signal_20212 ) ) ;
    buf_clk cell_5525 ( .C ( clk ), .D ( signal_20217 ), .Q ( signal_20218 ) ) ;
    buf_clk cell_5531 ( .C ( clk ), .D ( signal_20223 ), .Q ( signal_20224 ) ) ;
    buf_clk cell_5537 ( .C ( clk ), .D ( signal_20229 ), .Q ( signal_20230 ) ) ;
    buf_clk cell_5543 ( .C ( clk ), .D ( signal_20235 ), .Q ( signal_20236 ) ) ;
    buf_clk cell_5547 ( .C ( clk ), .D ( signal_20239 ), .Q ( signal_20240 ) ) ;
    buf_clk cell_5551 ( .C ( clk ), .D ( signal_20243 ), .Q ( signal_20244 ) ) ;
    buf_clk cell_5555 ( .C ( clk ), .D ( signal_20247 ), .Q ( signal_20248 ) ) ;
    buf_clk cell_5559 ( .C ( clk ), .D ( signal_20251 ), .Q ( signal_20252 ) ) ;
    buf_clk cell_5563 ( .C ( clk ), .D ( signal_20255 ), .Q ( signal_20256 ) ) ;
    buf_clk cell_5569 ( .C ( clk ), .D ( signal_20261 ), .Q ( signal_20262 ) ) ;
    buf_clk cell_5575 ( .C ( clk ), .D ( signal_20267 ), .Q ( signal_20268 ) ) ;
    buf_clk cell_5581 ( .C ( clk ), .D ( signal_20273 ), .Q ( signal_20274 ) ) ;
    buf_clk cell_5587 ( .C ( clk ), .D ( signal_20279 ), .Q ( signal_20280 ) ) ;
    buf_clk cell_5593 ( .C ( clk ), .D ( signal_20285 ), .Q ( signal_20286 ) ) ;
    buf_clk cell_5597 ( .C ( clk ), .D ( signal_20289 ), .Q ( signal_20290 ) ) ;
    buf_clk cell_5601 ( .C ( clk ), .D ( signal_20293 ), .Q ( signal_20294 ) ) ;
    buf_clk cell_5605 ( .C ( clk ), .D ( signal_20297 ), .Q ( signal_20298 ) ) ;
    buf_clk cell_5609 ( .C ( clk ), .D ( signal_20301 ), .Q ( signal_20302 ) ) ;
    buf_clk cell_5613 ( .C ( clk ), .D ( signal_20305 ), .Q ( signal_20306 ) ) ;
    buf_clk cell_5617 ( .C ( clk ), .D ( signal_20309 ), .Q ( signal_20310 ) ) ;
    buf_clk cell_5621 ( .C ( clk ), .D ( signal_20313 ), .Q ( signal_20314 ) ) ;
    buf_clk cell_5625 ( .C ( clk ), .D ( signal_20317 ), .Q ( signal_20318 ) ) ;
    buf_clk cell_5629 ( .C ( clk ), .D ( signal_20321 ), .Q ( signal_20322 ) ) ;
    buf_clk cell_5633 ( .C ( clk ), .D ( signal_20325 ), .Q ( signal_20326 ) ) ;
    buf_clk cell_5637 ( .C ( clk ), .D ( signal_20329 ), .Q ( signal_20330 ) ) ;
    buf_clk cell_5641 ( .C ( clk ), .D ( signal_20333 ), .Q ( signal_20334 ) ) ;
    buf_clk cell_5645 ( .C ( clk ), .D ( signal_20337 ), .Q ( signal_20338 ) ) ;
    buf_clk cell_5649 ( .C ( clk ), .D ( signal_20341 ), .Q ( signal_20342 ) ) ;
    buf_clk cell_5653 ( .C ( clk ), .D ( signal_20345 ), .Q ( signal_20346 ) ) ;
    buf_clk cell_5655 ( .C ( clk ), .D ( signal_1966 ), .Q ( signal_20348 ) ) ;
    buf_clk cell_5657 ( .C ( clk ), .D ( signal_6520 ), .Q ( signal_20350 ) ) ;
    buf_clk cell_5659 ( .C ( clk ), .D ( signal_6521 ), .Q ( signal_20352 ) ) ;
    buf_clk cell_5661 ( .C ( clk ), .D ( signal_6522 ), .Q ( signal_20354 ) ) ;
    buf_clk cell_5663 ( .C ( clk ), .D ( signal_6523 ), .Q ( signal_20356 ) ) ;
    buf_clk cell_5667 ( .C ( clk ), .D ( signal_20359 ), .Q ( signal_20360 ) ) ;
    buf_clk cell_5671 ( .C ( clk ), .D ( signal_20363 ), .Q ( signal_20364 ) ) ;
    buf_clk cell_5675 ( .C ( clk ), .D ( signal_20367 ), .Q ( signal_20368 ) ) ;
    buf_clk cell_5679 ( .C ( clk ), .D ( signal_20371 ), .Q ( signal_20372 ) ) ;
    buf_clk cell_5683 ( .C ( clk ), .D ( signal_20375 ), .Q ( signal_20376 ) ) ;
    buf_clk cell_5687 ( .C ( clk ), .D ( signal_20379 ), .Q ( signal_20380 ) ) ;
    buf_clk cell_5691 ( .C ( clk ), .D ( signal_20383 ), .Q ( signal_20384 ) ) ;
    buf_clk cell_5695 ( .C ( clk ), .D ( signal_20387 ), .Q ( signal_20388 ) ) ;
    buf_clk cell_5699 ( .C ( clk ), .D ( signal_20391 ), .Q ( signal_20392 ) ) ;
    buf_clk cell_5703 ( .C ( clk ), .D ( signal_20395 ), .Q ( signal_20396 ) ) ;
    buf_clk cell_5709 ( .C ( clk ), .D ( signal_20401 ), .Q ( signal_20402 ) ) ;
    buf_clk cell_5715 ( .C ( clk ), .D ( signal_20407 ), .Q ( signal_20408 ) ) ;
    buf_clk cell_5721 ( .C ( clk ), .D ( signal_20413 ), .Q ( signal_20414 ) ) ;
    buf_clk cell_5727 ( .C ( clk ), .D ( signal_20419 ), .Q ( signal_20420 ) ) ;
    buf_clk cell_5733 ( .C ( clk ), .D ( signal_20425 ), .Q ( signal_20426 ) ) ;
    buf_clk cell_5735 ( .C ( clk ), .D ( signal_2011 ), .Q ( signal_20428 ) ) ;
    buf_clk cell_5737 ( .C ( clk ), .D ( signal_6700 ), .Q ( signal_20430 ) ) ;
    buf_clk cell_5739 ( .C ( clk ), .D ( signal_6701 ), .Q ( signal_20432 ) ) ;
    buf_clk cell_5741 ( .C ( clk ), .D ( signal_6702 ), .Q ( signal_20434 ) ) ;
    buf_clk cell_5743 ( .C ( clk ), .D ( signal_6703 ), .Q ( signal_20436 ) ) ;
    buf_clk cell_5745 ( .C ( clk ), .D ( signal_1843 ), .Q ( signal_20438 ) ) ;
    buf_clk cell_5747 ( .C ( clk ), .D ( signal_6028 ), .Q ( signal_20440 ) ) ;
    buf_clk cell_5749 ( .C ( clk ), .D ( signal_6029 ), .Q ( signal_20442 ) ) ;
    buf_clk cell_5751 ( .C ( clk ), .D ( signal_6030 ), .Q ( signal_20444 ) ) ;
    buf_clk cell_5753 ( .C ( clk ), .D ( signal_6031 ), .Q ( signal_20446 ) ) ;
    buf_clk cell_5757 ( .C ( clk ), .D ( signal_20449 ), .Q ( signal_20450 ) ) ;
    buf_clk cell_5761 ( .C ( clk ), .D ( signal_20453 ), .Q ( signal_20454 ) ) ;
    buf_clk cell_5765 ( .C ( clk ), .D ( signal_20457 ), .Q ( signal_20458 ) ) ;
    buf_clk cell_5769 ( .C ( clk ), .D ( signal_20461 ), .Q ( signal_20462 ) ) ;
    buf_clk cell_5773 ( .C ( clk ), .D ( signal_20465 ), .Q ( signal_20466 ) ) ;
    buf_clk cell_5779 ( .C ( clk ), .D ( signal_20471 ), .Q ( signal_20472 ) ) ;
    buf_clk cell_5785 ( .C ( clk ), .D ( signal_20477 ), .Q ( signal_20478 ) ) ;
    buf_clk cell_5791 ( .C ( clk ), .D ( signal_20483 ), .Q ( signal_20484 ) ) ;
    buf_clk cell_5797 ( .C ( clk ), .D ( signal_20489 ), .Q ( signal_20490 ) ) ;
    buf_clk cell_5803 ( .C ( clk ), .D ( signal_20495 ), .Q ( signal_20496 ) ) ;
    buf_clk cell_5809 ( .C ( clk ), .D ( signal_20501 ), .Q ( signal_20502 ) ) ;
    buf_clk cell_5815 ( .C ( clk ), .D ( signal_20507 ), .Q ( signal_20508 ) ) ;
    buf_clk cell_5821 ( .C ( clk ), .D ( signal_20513 ), .Q ( signal_20514 ) ) ;
    buf_clk cell_5827 ( .C ( clk ), .D ( signal_20519 ), .Q ( signal_20520 ) ) ;
    buf_clk cell_5833 ( .C ( clk ), .D ( signal_20525 ), .Q ( signal_20526 ) ) ;
    buf_clk cell_5839 ( .C ( clk ), .D ( signal_20531 ), .Q ( signal_20532 ) ) ;
    buf_clk cell_5845 ( .C ( clk ), .D ( signal_20537 ), .Q ( signal_20538 ) ) ;
    buf_clk cell_5851 ( .C ( clk ), .D ( signal_20543 ), .Q ( signal_20544 ) ) ;
    buf_clk cell_5857 ( .C ( clk ), .D ( signal_20549 ), .Q ( signal_20550 ) ) ;
    buf_clk cell_5863 ( .C ( clk ), .D ( signal_20555 ), .Q ( signal_20556 ) ) ;
    buf_clk cell_5867 ( .C ( clk ), .D ( signal_20559 ), .Q ( signal_20560 ) ) ;
    buf_clk cell_5871 ( .C ( clk ), .D ( signal_20563 ), .Q ( signal_20564 ) ) ;
    buf_clk cell_5875 ( .C ( clk ), .D ( signal_20567 ), .Q ( signal_20568 ) ) ;
    buf_clk cell_5879 ( .C ( clk ), .D ( signal_20571 ), .Q ( signal_20572 ) ) ;
    buf_clk cell_5883 ( .C ( clk ), .D ( signal_20575 ), .Q ( signal_20576 ) ) ;
    buf_clk cell_5885 ( .C ( clk ), .D ( signal_19191 ), .Q ( signal_20578 ) ) ;
    buf_clk cell_5887 ( .C ( clk ), .D ( signal_19195 ), .Q ( signal_20580 ) ) ;
    buf_clk cell_5889 ( .C ( clk ), .D ( signal_19199 ), .Q ( signal_20582 ) ) ;
    buf_clk cell_5891 ( .C ( clk ), .D ( signal_19203 ), .Q ( signal_20584 ) ) ;
    buf_clk cell_5893 ( .C ( clk ), .D ( signal_19207 ), .Q ( signal_20586 ) ) ;
    buf_clk cell_5895 ( .C ( clk ), .D ( signal_19241 ), .Q ( signal_20588 ) ) ;
    buf_clk cell_5897 ( .C ( clk ), .D ( signal_19245 ), .Q ( signal_20590 ) ) ;
    buf_clk cell_5899 ( .C ( clk ), .D ( signal_19249 ), .Q ( signal_20592 ) ) ;
    buf_clk cell_5901 ( .C ( clk ), .D ( signal_19253 ), .Q ( signal_20594 ) ) ;
    buf_clk cell_5903 ( .C ( clk ), .D ( signal_19257 ), .Q ( signal_20596 ) ) ;
    buf_clk cell_5909 ( .C ( clk ), .D ( signal_20601 ), .Q ( signal_20602 ) ) ;
    buf_clk cell_5917 ( .C ( clk ), .D ( signal_20609 ), .Q ( signal_20610 ) ) ;
    buf_clk cell_5925 ( .C ( clk ), .D ( signal_20617 ), .Q ( signal_20618 ) ) ;
    buf_clk cell_5933 ( .C ( clk ), .D ( signal_20625 ), .Q ( signal_20626 ) ) ;
    buf_clk cell_5941 ( .C ( clk ), .D ( signal_20633 ), .Q ( signal_20634 ) ) ;
    buf_clk cell_5945 ( .C ( clk ), .D ( signal_1758 ), .Q ( signal_20638 ) ) ;
    buf_clk cell_5949 ( .C ( clk ), .D ( signal_5688 ), .Q ( signal_20642 ) ) ;
    buf_clk cell_5953 ( .C ( clk ), .D ( signal_5689 ), .Q ( signal_20646 ) ) ;
    buf_clk cell_5957 ( .C ( clk ), .D ( signal_5690 ), .Q ( signal_20650 ) ) ;
    buf_clk cell_5961 ( .C ( clk ), .D ( signal_5691 ), .Q ( signal_20654 ) ) ;
    buf_clk cell_5967 ( .C ( clk ), .D ( signal_20659 ), .Q ( signal_20660 ) ) ;
    buf_clk cell_5973 ( .C ( clk ), .D ( signal_20665 ), .Q ( signal_20666 ) ) ;
    buf_clk cell_5979 ( .C ( clk ), .D ( signal_20671 ), .Q ( signal_20672 ) ) ;
    buf_clk cell_5985 ( .C ( clk ), .D ( signal_20677 ), .Q ( signal_20678 ) ) ;
    buf_clk cell_5991 ( .C ( clk ), .D ( signal_20683 ), .Q ( signal_20684 ) ) ;
    buf_clk cell_5997 ( .C ( clk ), .D ( signal_20689 ), .Q ( signal_20690 ) ) ;
    buf_clk cell_6003 ( .C ( clk ), .D ( signal_20695 ), .Q ( signal_20696 ) ) ;
    buf_clk cell_6009 ( .C ( clk ), .D ( signal_20701 ), .Q ( signal_20702 ) ) ;
    buf_clk cell_6015 ( .C ( clk ), .D ( signal_20707 ), .Q ( signal_20708 ) ) ;
    buf_clk cell_6021 ( .C ( clk ), .D ( signal_20713 ), .Q ( signal_20714 ) ) ;
    buf_clk cell_6025 ( .C ( clk ), .D ( signal_1762 ), .Q ( signal_20718 ) ) ;
    buf_clk cell_6029 ( .C ( clk ), .D ( signal_5704 ), .Q ( signal_20722 ) ) ;
    buf_clk cell_6033 ( .C ( clk ), .D ( signal_5705 ), .Q ( signal_20726 ) ) ;
    buf_clk cell_6037 ( .C ( clk ), .D ( signal_5706 ), .Q ( signal_20730 ) ) ;
    buf_clk cell_6041 ( .C ( clk ), .D ( signal_5707 ), .Q ( signal_20734 ) ) ;
    buf_clk cell_6047 ( .C ( clk ), .D ( signal_20739 ), .Q ( signal_20740 ) ) ;
    buf_clk cell_6053 ( .C ( clk ), .D ( signal_20745 ), .Q ( signal_20746 ) ) ;
    buf_clk cell_6059 ( .C ( clk ), .D ( signal_20751 ), .Q ( signal_20752 ) ) ;
    buf_clk cell_6065 ( .C ( clk ), .D ( signal_20757 ), .Q ( signal_20758 ) ) ;
    buf_clk cell_6071 ( .C ( clk ), .D ( signal_20763 ), .Q ( signal_20764 ) ) ;
    buf_clk cell_6075 ( .C ( clk ), .D ( signal_19041 ), .Q ( signal_20768 ) ) ;
    buf_clk cell_6079 ( .C ( clk ), .D ( signal_19045 ), .Q ( signal_20772 ) ) ;
    buf_clk cell_6083 ( .C ( clk ), .D ( signal_19049 ), .Q ( signal_20776 ) ) ;
    buf_clk cell_6087 ( .C ( clk ), .D ( signal_19053 ), .Q ( signal_20780 ) ) ;
    buf_clk cell_6091 ( .C ( clk ), .D ( signal_19057 ), .Q ( signal_20784 ) ) ;
    buf_clk cell_6095 ( .C ( clk ), .D ( signal_1845 ), .Q ( signal_20788 ) ) ;
    buf_clk cell_6099 ( .C ( clk ), .D ( signal_6036 ), .Q ( signal_20792 ) ) ;
    buf_clk cell_6103 ( .C ( clk ), .D ( signal_6037 ), .Q ( signal_20796 ) ) ;
    buf_clk cell_6107 ( .C ( clk ), .D ( signal_6038 ), .Q ( signal_20800 ) ) ;
    buf_clk cell_6111 ( .C ( clk ), .D ( signal_6039 ), .Q ( signal_20804 ) ) ;
    buf_clk cell_6137 ( .C ( clk ), .D ( signal_20829 ), .Q ( signal_20830 ) ) ;
    buf_clk cell_6143 ( .C ( clk ), .D ( signal_20835 ), .Q ( signal_20836 ) ) ;
    buf_clk cell_6149 ( .C ( clk ), .D ( signal_20841 ), .Q ( signal_20842 ) ) ;
    buf_clk cell_6155 ( .C ( clk ), .D ( signal_20847 ), .Q ( signal_20848 ) ) ;
    buf_clk cell_6161 ( .C ( clk ), .D ( signal_20853 ), .Q ( signal_20854 ) ) ;
    buf_clk cell_6167 ( .C ( clk ), .D ( signal_20859 ), .Q ( signal_20860 ) ) ;
    buf_clk cell_6173 ( .C ( clk ), .D ( signal_20865 ), .Q ( signal_20866 ) ) ;
    buf_clk cell_6179 ( .C ( clk ), .D ( signal_20871 ), .Q ( signal_20872 ) ) ;
    buf_clk cell_6185 ( .C ( clk ), .D ( signal_20877 ), .Q ( signal_20878 ) ) ;
    buf_clk cell_6191 ( .C ( clk ), .D ( signal_20883 ), .Q ( signal_20884 ) ) ;
    buf_clk cell_6197 ( .C ( clk ), .D ( signal_20889 ), .Q ( signal_20890 ) ) ;
    buf_clk cell_6203 ( .C ( clk ), .D ( signal_20895 ), .Q ( signal_20896 ) ) ;
    buf_clk cell_6209 ( .C ( clk ), .D ( signal_20901 ), .Q ( signal_20902 ) ) ;
    buf_clk cell_6215 ( .C ( clk ), .D ( signal_20907 ), .Q ( signal_20908 ) ) ;
    buf_clk cell_6221 ( .C ( clk ), .D ( signal_20913 ), .Q ( signal_20914 ) ) ;
    buf_clk cell_6235 ( .C ( clk ), .D ( signal_1810 ), .Q ( signal_20928 ) ) ;
    buf_clk cell_6239 ( .C ( clk ), .D ( signal_5896 ), .Q ( signal_20932 ) ) ;
    buf_clk cell_6243 ( .C ( clk ), .D ( signal_5897 ), .Q ( signal_20936 ) ) ;
    buf_clk cell_6247 ( .C ( clk ), .D ( signal_5898 ), .Q ( signal_20940 ) ) ;
    buf_clk cell_6251 ( .C ( clk ), .D ( signal_5899 ), .Q ( signal_20944 ) ) ;
    buf_clk cell_6257 ( .C ( clk ), .D ( signal_20949 ), .Q ( signal_20950 ) ) ;
    buf_clk cell_6263 ( .C ( clk ), .D ( signal_20955 ), .Q ( signal_20956 ) ) ;
    buf_clk cell_6269 ( .C ( clk ), .D ( signal_20961 ), .Q ( signal_20962 ) ) ;
    buf_clk cell_6275 ( .C ( clk ), .D ( signal_20967 ), .Q ( signal_20968 ) ) ;
    buf_clk cell_6281 ( .C ( clk ), .D ( signal_20973 ), .Q ( signal_20974 ) ) ;
    buf_clk cell_6297 ( .C ( clk ), .D ( signal_20989 ), .Q ( signal_20990 ) ) ;
    buf_clk cell_6303 ( .C ( clk ), .D ( signal_20995 ), .Q ( signal_20996 ) ) ;
    buf_clk cell_6309 ( .C ( clk ), .D ( signal_21001 ), .Q ( signal_21002 ) ) ;
    buf_clk cell_6315 ( .C ( clk ), .D ( signal_21007 ), .Q ( signal_21008 ) ) ;
    buf_clk cell_6321 ( .C ( clk ), .D ( signal_21013 ), .Q ( signal_21014 ) ) ;
    buf_clk cell_6339 ( .C ( clk ), .D ( signal_21031 ), .Q ( signal_21032 ) ) ;
    buf_clk cell_6347 ( .C ( clk ), .D ( signal_21039 ), .Q ( signal_21040 ) ) ;
    buf_clk cell_6355 ( .C ( clk ), .D ( signal_21047 ), .Q ( signal_21048 ) ) ;
    buf_clk cell_6363 ( .C ( clk ), .D ( signal_21055 ), .Q ( signal_21056 ) ) ;
    buf_clk cell_6371 ( .C ( clk ), .D ( signal_21063 ), .Q ( signal_21064 ) ) ;
    buf_clk cell_6375 ( .C ( clk ), .D ( signal_1814 ), .Q ( signal_21068 ) ) ;
    buf_clk cell_6379 ( .C ( clk ), .D ( signal_5912 ), .Q ( signal_21072 ) ) ;
    buf_clk cell_6383 ( .C ( clk ), .D ( signal_5913 ), .Q ( signal_21076 ) ) ;
    buf_clk cell_6387 ( .C ( clk ), .D ( signal_5914 ), .Q ( signal_21080 ) ) ;
    buf_clk cell_6391 ( .C ( clk ), .D ( signal_5915 ), .Q ( signal_21084 ) ) ;
    buf_clk cell_6395 ( .C ( clk ), .D ( signal_1820 ), .Q ( signal_21088 ) ) ;
    buf_clk cell_6399 ( .C ( clk ), .D ( signal_5936 ), .Q ( signal_21092 ) ) ;
    buf_clk cell_6403 ( .C ( clk ), .D ( signal_5937 ), .Q ( signal_21096 ) ) ;
    buf_clk cell_6407 ( .C ( clk ), .D ( signal_5938 ), .Q ( signal_21100 ) ) ;
    buf_clk cell_6411 ( .C ( clk ), .D ( signal_5939 ), .Q ( signal_21104 ) ) ;
    buf_clk cell_6417 ( .C ( clk ), .D ( signal_21109 ), .Q ( signal_21110 ) ) ;
    buf_clk cell_6423 ( .C ( clk ), .D ( signal_21115 ), .Q ( signal_21116 ) ) ;
    buf_clk cell_6429 ( .C ( clk ), .D ( signal_21121 ), .Q ( signal_21122 ) ) ;
    buf_clk cell_6435 ( .C ( clk ), .D ( signal_21127 ), .Q ( signal_21128 ) ) ;
    buf_clk cell_6441 ( .C ( clk ), .D ( signal_21133 ), .Q ( signal_21134 ) ) ;
    buf_clk cell_6447 ( .C ( clk ), .D ( signal_21139 ), .Q ( signal_21140 ) ) ;
    buf_clk cell_6453 ( .C ( clk ), .D ( signal_21145 ), .Q ( signal_21146 ) ) ;
    buf_clk cell_6459 ( .C ( clk ), .D ( signal_21151 ), .Q ( signal_21152 ) ) ;
    buf_clk cell_6465 ( .C ( clk ), .D ( signal_21157 ), .Q ( signal_21158 ) ) ;
    buf_clk cell_6471 ( .C ( clk ), .D ( signal_21163 ), .Q ( signal_21164 ) ) ;
    buf_clk cell_6475 ( .C ( clk ), .D ( signal_2006 ), .Q ( signal_21168 ) ) ;
    buf_clk cell_6479 ( .C ( clk ), .D ( signal_6680 ), .Q ( signal_21172 ) ) ;
    buf_clk cell_6483 ( .C ( clk ), .D ( signal_6681 ), .Q ( signal_21176 ) ) ;
    buf_clk cell_6487 ( .C ( clk ), .D ( signal_6682 ), .Q ( signal_21180 ) ) ;
    buf_clk cell_6491 ( .C ( clk ), .D ( signal_6683 ), .Q ( signal_21184 ) ) ;
    buf_clk cell_6499 ( .C ( clk ), .D ( signal_21191 ), .Q ( signal_21192 ) ) ;
    buf_clk cell_6507 ( .C ( clk ), .D ( signal_21199 ), .Q ( signal_21200 ) ) ;
    buf_clk cell_6515 ( .C ( clk ), .D ( signal_21207 ), .Q ( signal_21208 ) ) ;
    buf_clk cell_6523 ( .C ( clk ), .D ( signal_21215 ), .Q ( signal_21216 ) ) ;
    buf_clk cell_6531 ( .C ( clk ), .D ( signal_21223 ), .Q ( signal_21224 ) ) ;
    buf_clk cell_6537 ( .C ( clk ), .D ( signal_21229 ), .Q ( signal_21230 ) ) ;
    buf_clk cell_6543 ( .C ( clk ), .D ( signal_21235 ), .Q ( signal_21236 ) ) ;
    buf_clk cell_6549 ( .C ( clk ), .D ( signal_21241 ), .Q ( signal_21242 ) ) ;
    buf_clk cell_6555 ( .C ( clk ), .D ( signal_21247 ), .Q ( signal_21248 ) ) ;
    buf_clk cell_6561 ( .C ( clk ), .D ( signal_21253 ), .Q ( signal_21254 ) ) ;
    buf_clk cell_6567 ( .C ( clk ), .D ( signal_21259 ), .Q ( signal_21260 ) ) ;
    buf_clk cell_6573 ( .C ( clk ), .D ( signal_21265 ), .Q ( signal_21266 ) ) ;
    buf_clk cell_6579 ( .C ( clk ), .D ( signal_21271 ), .Q ( signal_21272 ) ) ;
    buf_clk cell_6585 ( .C ( clk ), .D ( signal_21277 ), .Q ( signal_21278 ) ) ;
    buf_clk cell_6591 ( .C ( clk ), .D ( signal_21283 ), .Q ( signal_21284 ) ) ;
    buf_clk cell_6617 ( .C ( clk ), .D ( signal_21309 ), .Q ( signal_21310 ) ) ;
    buf_clk cell_6623 ( .C ( clk ), .D ( signal_21315 ), .Q ( signal_21316 ) ) ;
    buf_clk cell_6629 ( .C ( clk ), .D ( signal_21321 ), .Q ( signal_21322 ) ) ;
    buf_clk cell_6635 ( .C ( clk ), .D ( signal_21327 ), .Q ( signal_21328 ) ) ;
    buf_clk cell_6641 ( .C ( clk ), .D ( signal_21333 ), .Q ( signal_21334 ) ) ;
    buf_clk cell_6667 ( .C ( clk ), .D ( signal_21359 ), .Q ( signal_21360 ) ) ;
    buf_clk cell_6673 ( .C ( clk ), .D ( signal_21365 ), .Q ( signal_21366 ) ) ;
    buf_clk cell_6679 ( .C ( clk ), .D ( signal_21371 ), .Q ( signal_21372 ) ) ;
    buf_clk cell_6685 ( .C ( clk ), .D ( signal_21377 ), .Q ( signal_21378 ) ) ;
    buf_clk cell_6691 ( .C ( clk ), .D ( signal_21383 ), .Q ( signal_21384 ) ) ;
    buf_clk cell_6697 ( .C ( clk ), .D ( signal_21389 ), .Q ( signal_21390 ) ) ;
    buf_clk cell_6703 ( .C ( clk ), .D ( signal_21395 ), .Q ( signal_21396 ) ) ;
    buf_clk cell_6709 ( .C ( clk ), .D ( signal_21401 ), .Q ( signal_21402 ) ) ;
    buf_clk cell_6715 ( .C ( clk ), .D ( signal_21407 ), .Q ( signal_21408 ) ) ;
    buf_clk cell_6721 ( .C ( clk ), .D ( signal_21413 ), .Q ( signal_21414 ) ) ;
    buf_clk cell_6725 ( .C ( clk ), .D ( signal_1818 ), .Q ( signal_21418 ) ) ;
    buf_clk cell_6729 ( .C ( clk ), .D ( signal_5928 ), .Q ( signal_21422 ) ) ;
    buf_clk cell_6733 ( .C ( clk ), .D ( signal_5929 ), .Q ( signal_21426 ) ) ;
    buf_clk cell_6737 ( .C ( clk ), .D ( signal_5930 ), .Q ( signal_21430 ) ) ;
    buf_clk cell_6741 ( .C ( clk ), .D ( signal_5931 ), .Q ( signal_21434 ) ) ;
    buf_clk cell_6749 ( .C ( clk ), .D ( signal_21441 ), .Q ( signal_21442 ) ) ;
    buf_clk cell_6759 ( .C ( clk ), .D ( signal_21451 ), .Q ( signal_21452 ) ) ;
    buf_clk cell_6769 ( .C ( clk ), .D ( signal_21461 ), .Q ( signal_21462 ) ) ;
    buf_clk cell_6779 ( .C ( clk ), .D ( signal_21471 ), .Q ( signal_21472 ) ) ;
    buf_clk cell_6789 ( .C ( clk ), .D ( signal_21481 ), .Q ( signal_21482 ) ) ;
    buf_clk cell_6795 ( .C ( clk ), .D ( signal_1988 ), .Q ( signal_21488 ) ) ;
    buf_clk cell_6801 ( .C ( clk ), .D ( signal_6608 ), .Q ( signal_21494 ) ) ;
    buf_clk cell_6807 ( .C ( clk ), .D ( signal_6609 ), .Q ( signal_21500 ) ) ;
    buf_clk cell_6813 ( .C ( clk ), .D ( signal_6610 ), .Q ( signal_21506 ) ) ;
    buf_clk cell_6819 ( .C ( clk ), .D ( signal_6611 ), .Q ( signal_21512 ) ) ;
    buf_clk cell_6827 ( .C ( clk ), .D ( signal_21519 ), .Q ( signal_21520 ) ) ;
    buf_clk cell_6835 ( .C ( clk ), .D ( signal_21527 ), .Q ( signal_21528 ) ) ;
    buf_clk cell_6843 ( .C ( clk ), .D ( signal_21535 ), .Q ( signal_21536 ) ) ;
    buf_clk cell_6851 ( .C ( clk ), .D ( signal_21543 ), .Q ( signal_21544 ) ) ;
    buf_clk cell_6859 ( .C ( clk ), .D ( signal_21551 ), .Q ( signal_21552 ) ) ;
    buf_clk cell_6867 ( .C ( clk ), .D ( signal_21559 ), .Q ( signal_21560 ) ) ;
    buf_clk cell_6875 ( .C ( clk ), .D ( signal_21567 ), .Q ( signal_21568 ) ) ;
    buf_clk cell_6883 ( .C ( clk ), .D ( signal_21575 ), .Q ( signal_21576 ) ) ;
    buf_clk cell_6891 ( .C ( clk ), .D ( signal_21583 ), .Q ( signal_21584 ) ) ;
    buf_clk cell_6899 ( .C ( clk ), .D ( signal_21591 ), .Q ( signal_21592 ) ) ;
    buf_clk cell_6989 ( .C ( clk ), .D ( signal_21681 ), .Q ( signal_21682 ) ) ;
    buf_clk cell_6999 ( .C ( clk ), .D ( signal_21691 ), .Q ( signal_21692 ) ) ;
    buf_clk cell_7009 ( .C ( clk ), .D ( signal_21701 ), .Q ( signal_21702 ) ) ;
    buf_clk cell_7019 ( .C ( clk ), .D ( signal_21711 ), .Q ( signal_21712 ) ) ;
    buf_clk cell_7029 ( .C ( clk ), .D ( signal_21721 ), .Q ( signal_21722 ) ) ;
    buf_clk cell_7035 ( .C ( clk ), .D ( signal_2016 ), .Q ( signal_21728 ) ) ;
    buf_clk cell_7041 ( .C ( clk ), .D ( signal_6720 ), .Q ( signal_21734 ) ) ;
    buf_clk cell_7047 ( .C ( clk ), .D ( signal_6721 ), .Q ( signal_21740 ) ) ;
    buf_clk cell_7053 ( .C ( clk ), .D ( signal_6722 ), .Q ( signal_21746 ) ) ;
    buf_clk cell_7059 ( .C ( clk ), .D ( signal_6723 ), .Q ( signal_21752 ) ) ;
    buf_clk cell_7077 ( .C ( clk ), .D ( signal_21769 ), .Q ( signal_21770 ) ) ;
    buf_clk cell_7085 ( .C ( clk ), .D ( signal_21777 ), .Q ( signal_21778 ) ) ;
    buf_clk cell_7093 ( .C ( clk ), .D ( signal_21785 ), .Q ( signal_21786 ) ) ;
    buf_clk cell_7101 ( .C ( clk ), .D ( signal_21793 ), .Q ( signal_21794 ) ) ;
    buf_clk cell_7109 ( .C ( clk ), .D ( signal_21801 ), .Q ( signal_21802 ) ) ;
    buf_clk cell_7115 ( .C ( clk ), .D ( signal_1979 ), .Q ( signal_21808 ) ) ;
    buf_clk cell_7121 ( .C ( clk ), .D ( signal_6572 ), .Q ( signal_21814 ) ) ;
    buf_clk cell_7127 ( .C ( clk ), .D ( signal_6573 ), .Q ( signal_21820 ) ) ;
    buf_clk cell_7133 ( .C ( clk ), .D ( signal_6574 ), .Q ( signal_21826 ) ) ;
    buf_clk cell_7139 ( .C ( clk ), .D ( signal_6575 ), .Q ( signal_21832 ) ) ;
    buf_clk cell_7147 ( .C ( clk ), .D ( signal_21839 ), .Q ( signal_21840 ) ) ;
    buf_clk cell_7155 ( .C ( clk ), .D ( signal_21847 ), .Q ( signal_21848 ) ) ;
    buf_clk cell_7163 ( .C ( clk ), .D ( signal_21855 ), .Q ( signal_21856 ) ) ;
    buf_clk cell_7171 ( .C ( clk ), .D ( signal_21863 ), .Q ( signal_21864 ) ) ;
    buf_clk cell_7179 ( .C ( clk ), .D ( signal_21871 ), .Q ( signal_21872 ) ) ;
    buf_clk cell_7187 ( .C ( clk ), .D ( signal_21879 ), .Q ( signal_21880 ) ) ;
    buf_clk cell_7195 ( .C ( clk ), .D ( signal_21887 ), .Q ( signal_21888 ) ) ;
    buf_clk cell_7203 ( .C ( clk ), .D ( signal_21895 ), .Q ( signal_21896 ) ) ;
    buf_clk cell_7211 ( .C ( clk ), .D ( signal_21903 ), .Q ( signal_21904 ) ) ;
    buf_clk cell_7219 ( .C ( clk ), .D ( signal_21911 ), .Q ( signal_21912 ) ) ;
    buf_clk cell_7227 ( .C ( clk ), .D ( signal_21919 ), .Q ( signal_21920 ) ) ;
    buf_clk cell_7235 ( .C ( clk ), .D ( signal_21927 ), .Q ( signal_21928 ) ) ;
    buf_clk cell_7243 ( .C ( clk ), .D ( signal_21935 ), .Q ( signal_21936 ) ) ;
    buf_clk cell_7251 ( .C ( clk ), .D ( signal_21943 ), .Q ( signal_21944 ) ) ;
    buf_clk cell_7259 ( .C ( clk ), .D ( signal_21951 ), .Q ( signal_21952 ) ) ;
    buf_clk cell_7269 ( .C ( clk ), .D ( signal_21961 ), .Q ( signal_21962 ) ) ;
    buf_clk cell_7279 ( .C ( clk ), .D ( signal_21971 ), .Q ( signal_21972 ) ) ;
    buf_clk cell_7289 ( .C ( clk ), .D ( signal_21981 ), .Q ( signal_21982 ) ) ;
    buf_clk cell_7299 ( .C ( clk ), .D ( signal_21991 ), .Q ( signal_21992 ) ) ;
    buf_clk cell_7309 ( .C ( clk ), .D ( signal_22001 ), .Q ( signal_22002 ) ) ;
    buf_clk cell_7317 ( .C ( clk ), .D ( signal_22009 ), .Q ( signal_22010 ) ) ;
    buf_clk cell_7325 ( .C ( clk ), .D ( signal_22017 ), .Q ( signal_22018 ) ) ;
    buf_clk cell_7333 ( .C ( clk ), .D ( signal_22025 ), .Q ( signal_22026 ) ) ;
    buf_clk cell_7341 ( .C ( clk ), .D ( signal_22033 ), .Q ( signal_22034 ) ) ;
    buf_clk cell_7349 ( .C ( clk ), .D ( signal_22041 ), .Q ( signal_22042 ) ) ;
    buf_clk cell_7357 ( .C ( clk ), .D ( signal_22049 ), .Q ( signal_22050 ) ) ;
    buf_clk cell_7365 ( .C ( clk ), .D ( signal_22057 ), .Q ( signal_22058 ) ) ;
    buf_clk cell_7373 ( .C ( clk ), .D ( signal_22065 ), .Q ( signal_22066 ) ) ;
    buf_clk cell_7381 ( .C ( clk ), .D ( signal_22073 ), .Q ( signal_22074 ) ) ;
    buf_clk cell_7389 ( .C ( clk ), .D ( signal_22081 ), .Q ( signal_22082 ) ) ;
    buf_clk cell_7407 ( .C ( clk ), .D ( signal_22099 ), .Q ( signal_22100 ) ) ;
    buf_clk cell_7415 ( .C ( clk ), .D ( signal_22107 ), .Q ( signal_22108 ) ) ;
    buf_clk cell_7423 ( .C ( clk ), .D ( signal_22115 ), .Q ( signal_22116 ) ) ;
    buf_clk cell_7431 ( .C ( clk ), .D ( signal_22123 ), .Q ( signal_22124 ) ) ;
    buf_clk cell_7439 ( .C ( clk ), .D ( signal_22131 ), .Q ( signal_22132 ) ) ;
    buf_clk cell_7447 ( .C ( clk ), .D ( signal_22139 ), .Q ( signal_22140 ) ) ;
    buf_clk cell_7455 ( .C ( clk ), .D ( signal_22147 ), .Q ( signal_22148 ) ) ;
    buf_clk cell_7463 ( .C ( clk ), .D ( signal_22155 ), .Q ( signal_22156 ) ) ;
    buf_clk cell_7471 ( .C ( clk ), .D ( signal_22163 ), .Q ( signal_22164 ) ) ;
    buf_clk cell_7479 ( .C ( clk ), .D ( signal_22171 ), .Q ( signal_22172 ) ) ;
    buf_clk cell_7487 ( .C ( clk ), .D ( signal_22179 ), .Q ( signal_22180 ) ) ;
    buf_clk cell_7495 ( .C ( clk ), .D ( signal_22187 ), .Q ( signal_22188 ) ) ;
    buf_clk cell_7503 ( .C ( clk ), .D ( signal_22195 ), .Q ( signal_22196 ) ) ;
    buf_clk cell_7511 ( .C ( clk ), .D ( signal_22203 ), .Q ( signal_22204 ) ) ;
    buf_clk cell_7519 ( .C ( clk ), .D ( signal_22211 ), .Q ( signal_22212 ) ) ;
    buf_clk cell_7555 ( .C ( clk ), .D ( signal_2030 ), .Q ( signal_22248 ) ) ;
    buf_clk cell_7563 ( .C ( clk ), .D ( signal_6776 ), .Q ( signal_22256 ) ) ;
    buf_clk cell_7571 ( .C ( clk ), .D ( signal_6777 ), .Q ( signal_22264 ) ) ;
    buf_clk cell_7579 ( .C ( clk ), .D ( signal_6778 ), .Q ( signal_22272 ) ) ;
    buf_clk cell_7587 ( .C ( clk ), .D ( signal_6779 ), .Q ( signal_22280 ) ) ;
    buf_clk cell_7655 ( .C ( clk ), .D ( signal_19559 ), .Q ( signal_22348 ) ) ;
    buf_clk cell_7663 ( .C ( clk ), .D ( signal_19561 ), .Q ( signal_22356 ) ) ;
    buf_clk cell_7671 ( .C ( clk ), .D ( signal_19563 ), .Q ( signal_22364 ) ) ;
    buf_clk cell_7679 ( .C ( clk ), .D ( signal_19565 ), .Q ( signal_22372 ) ) ;
    buf_clk cell_7687 ( .C ( clk ), .D ( signal_19567 ), .Q ( signal_22380 ) ) ;
    buf_clk cell_7697 ( .C ( clk ), .D ( signal_22389 ), .Q ( signal_22390 ) ) ;
    buf_clk cell_7707 ( .C ( clk ), .D ( signal_22399 ), .Q ( signal_22400 ) ) ;
    buf_clk cell_7717 ( .C ( clk ), .D ( signal_22409 ), .Q ( signal_22410 ) ) ;
    buf_clk cell_7727 ( .C ( clk ), .D ( signal_22419 ), .Q ( signal_22420 ) ) ;
    buf_clk cell_7737 ( .C ( clk ), .D ( signal_22429 ), .Q ( signal_22430 ) ) ;
    buf_clk cell_7785 ( .C ( clk ), .D ( signal_1982 ), .Q ( signal_22478 ) ) ;
    buf_clk cell_7793 ( .C ( clk ), .D ( signal_6584 ), .Q ( signal_22486 ) ) ;
    buf_clk cell_7801 ( .C ( clk ), .D ( signal_6585 ), .Q ( signal_22494 ) ) ;
    buf_clk cell_7809 ( .C ( clk ), .D ( signal_6586 ), .Q ( signal_22502 ) ) ;
    buf_clk cell_7817 ( .C ( clk ), .D ( signal_6587 ), .Q ( signal_22510 ) ) ;
    buf_clk cell_7827 ( .C ( clk ), .D ( signal_22519 ), .Q ( signal_22520 ) ) ;
    buf_clk cell_7837 ( .C ( clk ), .D ( signal_22529 ), .Q ( signal_22530 ) ) ;
    buf_clk cell_7847 ( .C ( clk ), .D ( signal_22539 ), .Q ( signal_22540 ) ) ;
    buf_clk cell_7857 ( .C ( clk ), .D ( signal_22549 ), .Q ( signal_22550 ) ) ;
    buf_clk cell_7867 ( .C ( clk ), .D ( signal_22559 ), .Q ( signal_22560 ) ) ;
    buf_clk cell_7875 ( .C ( clk ), .D ( signal_1967 ), .Q ( signal_22568 ) ) ;
    buf_clk cell_7883 ( .C ( clk ), .D ( signal_6524 ), .Q ( signal_22576 ) ) ;
    buf_clk cell_7891 ( .C ( clk ), .D ( signal_6525 ), .Q ( signal_22584 ) ) ;
    buf_clk cell_7899 ( .C ( clk ), .D ( signal_6526 ), .Q ( signal_22592 ) ) ;
    buf_clk cell_7907 ( .C ( clk ), .D ( signal_6527 ), .Q ( signal_22600 ) ) ;
    buf_clk cell_8275 ( .C ( clk ), .D ( signal_1978 ), .Q ( signal_22968 ) ) ;
    buf_clk cell_8285 ( .C ( clk ), .D ( signal_6568 ), .Q ( signal_22978 ) ) ;
    buf_clk cell_8295 ( .C ( clk ), .D ( signal_6569 ), .Q ( signal_22988 ) ) ;
    buf_clk cell_8305 ( .C ( clk ), .D ( signal_6570 ), .Q ( signal_22998 ) ) ;
    buf_clk cell_8315 ( .C ( clk ), .D ( signal_6571 ), .Q ( signal_23008 ) ) ;
    buf_clk cell_8715 ( .C ( clk ), .D ( signal_1736 ), .Q ( signal_23408 ) ) ;
    buf_clk cell_8727 ( .C ( clk ), .D ( signal_5600 ), .Q ( signal_23420 ) ) ;
    buf_clk cell_8739 ( .C ( clk ), .D ( signal_5601 ), .Q ( signal_23432 ) ) ;
    buf_clk cell_8751 ( .C ( clk ), .D ( signal_5602 ), .Q ( signal_23444 ) ) ;
    buf_clk cell_8763 ( .C ( clk ), .D ( signal_5603 ), .Q ( signal_23456 ) ) ;
    buf_clk cell_8837 ( .C ( clk ), .D ( signal_23529 ), .Q ( signal_23530 ) ) ;
    buf_clk cell_8851 ( .C ( clk ), .D ( signal_23543 ), .Q ( signal_23544 ) ) ;
    buf_clk cell_8865 ( .C ( clk ), .D ( signal_23557 ), .Q ( signal_23558 ) ) ;
    buf_clk cell_8879 ( .C ( clk ), .D ( signal_23571 ), .Q ( signal_23572 ) ) ;
    buf_clk cell_8893 ( .C ( clk ), .D ( signal_23585 ), .Q ( signal_23586 ) ) ;
    buf_clk cell_8947 ( .C ( clk ), .D ( signal_23639 ), .Q ( signal_23640 ) ) ;
    buf_clk cell_8961 ( .C ( clk ), .D ( signal_23653 ), .Q ( signal_23654 ) ) ;
    buf_clk cell_8975 ( .C ( clk ), .D ( signal_23667 ), .Q ( signal_23668 ) ) ;
    buf_clk cell_8989 ( .C ( clk ), .D ( signal_23681 ), .Q ( signal_23682 ) ) ;
    buf_clk cell_9003 ( .C ( clk ), .D ( signal_23695 ), .Q ( signal_23696 ) ) ;
    buf_clk cell_9147 ( .C ( clk ), .D ( signal_23839 ), .Q ( signal_23840 ) ) ;
    buf_clk cell_9163 ( .C ( clk ), .D ( signal_23855 ), .Q ( signal_23856 ) ) ;
    buf_clk cell_9179 ( .C ( clk ), .D ( signal_23871 ), .Q ( signal_23872 ) ) ;
    buf_clk cell_9195 ( .C ( clk ), .D ( signal_23887 ), .Q ( signal_23888 ) ) ;
    buf_clk cell_9211 ( .C ( clk ), .D ( signal_23903 ), .Q ( signal_23904 ) ) ;
    buf_clk cell_9247 ( .C ( clk ), .D ( signal_23939 ), .Q ( signal_23940 ) ) ;
    buf_clk cell_9263 ( .C ( clk ), .D ( signal_23955 ), .Q ( signal_23956 ) ) ;
    buf_clk cell_9279 ( .C ( clk ), .D ( signal_23971 ), .Q ( signal_23972 ) ) ;
    buf_clk cell_9295 ( .C ( clk ), .D ( signal_23987 ), .Q ( signal_23988 ) ) ;
    buf_clk cell_9311 ( .C ( clk ), .D ( signal_24003 ), .Q ( signal_24004 ) ) ;
    buf_clk cell_9555 ( .C ( clk ), .D ( signal_1783 ), .Q ( signal_24248 ) ) ;
    buf_clk cell_9571 ( .C ( clk ), .D ( signal_5788 ), .Q ( signal_24264 ) ) ;
    buf_clk cell_9587 ( .C ( clk ), .D ( signal_5789 ), .Q ( signal_24280 ) ) ;
    buf_clk cell_9603 ( .C ( clk ), .D ( signal_5790 ), .Q ( signal_24296 ) ) ;
    buf_clk cell_9619 ( .C ( clk ), .D ( signal_5791 ), .Q ( signal_24312 ) ) ;
    buf_clk cell_9637 ( .C ( clk ), .D ( signal_24329 ), .Q ( signal_24330 ) ) ;
    buf_clk cell_9655 ( .C ( clk ), .D ( signal_24347 ), .Q ( signal_24348 ) ) ;
    buf_clk cell_9673 ( .C ( clk ), .D ( signal_24365 ), .Q ( signal_24366 ) ) ;
    buf_clk cell_9691 ( .C ( clk ), .D ( signal_24383 ), .Q ( signal_24384 ) ) ;
    buf_clk cell_9709 ( .C ( clk ), .D ( signal_24401 ), .Q ( signal_24402 ) ) ;
    buf_clk cell_9887 ( .C ( clk ), .D ( signal_24579 ), .Q ( signal_24580 ) ) ;
    buf_clk cell_9907 ( .C ( clk ), .D ( signal_24599 ), .Q ( signal_24600 ) ) ;
    buf_clk cell_9927 ( .C ( clk ), .D ( signal_24619 ), .Q ( signal_24620 ) ) ;
    buf_clk cell_9947 ( .C ( clk ), .D ( signal_24639 ), .Q ( signal_24640 ) ) ;
    buf_clk cell_9967 ( .C ( clk ), .D ( signal_24659 ), .Q ( signal_24660 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1819 ( .a ({signal_18667, signal_18665, signal_18663, signal_18661, signal_18659}), .b ({signal_5407, signal_5406, signal_5405, signal_5404, signal_1687}), .clk ( clk ), .r ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810]}), .c ({signal_5995, signal_5994, signal_5993, signal_5992, signal_1834}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1834 ( .a ({signal_18677, signal_18675, signal_18673, signal_18671, signal_18669}), .b ({signal_5499, signal_5498, signal_5497, signal_5496, signal_1710}), .clk ( clk ), .r ({Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .c ({signal_6055, signal_6054, signal_6053, signal_6052, signal_1849}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1872 ( .a ({signal_5995, signal_5994, signal_5993, signal_5992, signal_1834}), .b ({signal_6207, signal_6206, signal_6205, signal_6204, signal_1887}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1875 ( .a ({signal_6055, signal_6054, signal_6053, signal_6052, signal_1849}), .b ({signal_6219, signal_6218, signal_6217, signal_6216, signal_1890}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1893 ( .a ({signal_18697, signal_18693, signal_18689, signal_18685, signal_18681}), .b ({signal_5579, signal_5578, signal_5577, signal_5576, signal_1730}), .clk ( clk ), .r ({Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830]}), .c ({signal_6291, signal_6290, signal_6289, signal_6288, signal_1908}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1902 ( .a ({signal_5727, signal_5726, signal_5725, signal_5724, signal_1767}), .b ({signal_5803, signal_5802, signal_5801, signal_5800, signal_1786}), .clk ( clk ), .r ({Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840]}), .c ({signal_6327, signal_6326, signal_6325, signal_6324, signal_1917}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1904 ( .a ({signal_18697, signal_18693, signal_18689, signal_18685, signal_18681}), .b ({signal_5619, signal_5618, signal_5617, signal_5616, signal_1740}), .clk ( clk ), .r ({Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850]}), .c ({signal_6335, signal_6334, signal_6333, signal_6332, signal_1919}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1911 ( .a ({signal_5819, signal_5818, signal_5817, signal_5816, signal_1790}), .b ({signal_18707, signal_18705, signal_18703, signal_18701, signal_18699}), .clk ( clk ), .r ({Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860]}), .c ({signal_6363, signal_6362, signal_6361, signal_6360, signal_1926}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1912 ( .a ({signal_18727, signal_18723, signal_18719, signal_18715, signal_18711}), .b ({signal_5827, signal_5826, signal_5825, signal_5824, signal_1792}), .clk ( clk ), .r ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870]}), .c ({signal_6367, signal_6366, signal_6365, signal_6364, signal_1927}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1918 ( .a ({signal_18747, signal_18743, signal_18739, signal_18735, signal_18731}), .b ({signal_5875, signal_5874, signal_5873, signal_5872, signal_1804}), .clk ( clk ), .r ({Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .c ({signal_6391, signal_6390, signal_6389, signal_6388, signal_1933}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1921 ( .a ({signal_18767, signal_18763, signal_18759, signal_18755, signal_18751}), .b ({signal_5883, signal_5882, signal_5881, signal_5880, signal_1806}), .clk ( clk ), .r ({Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890]}), .c ({signal_6403, signal_6402, signal_6401, signal_6400, signal_1936}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1922 ( .a ({signal_5891, signal_5890, signal_5889, signal_5888, signal_1808}), .b ({signal_5895, signal_5894, signal_5893, signal_5892, signal_1809}), .clk ( clk ), .r ({Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900]}), .c ({signal_6407, signal_6406, signal_6405, signal_6404, signal_1937}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1924 ( .a ({signal_18807, signal_18799, signal_18791, signal_18783, signal_18775}), .b ({signal_5667, signal_5666, signal_5665, signal_5664, signal_1752}), .clk ( clk ), .r ({Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910]}), .c ({signal_6415, signal_6414, signal_6413, signal_6412, signal_1939}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1925 ( .a ({signal_18817, signal_18815, signal_18813, signal_18811, signal_18809}), .b ({signal_5919, signal_5918, signal_5917, signal_5916, signal_1815}), .clk ( clk ), .r ({Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920]}), .c ({signal_6419, signal_6418, signal_6417, signal_6416, signal_1940}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1926 ( .a ({signal_18827, signal_18825, signal_18823, signal_18821, signal_18819}), .b ({signal_5671, signal_5670, signal_5669, signal_5668, signal_1753}), .clk ( clk ), .r ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930]}), .c ({signal_6423, signal_6422, signal_6421, signal_6420, signal_1941}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1928 ( .a ({signal_18847, signal_18843, signal_18839, signal_18835, signal_18831}), .b ({signal_5935, signal_5934, signal_5933, signal_5932, signal_1819}), .clk ( clk ), .r ({Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .c ({signal_6431, signal_6430, signal_6429, signal_6428, signal_1943}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1929 ( .a ({signal_5815, signal_5814, signal_5813, signal_5812, signal_1789}), .b ({signal_18857, signal_18855, signal_18853, signal_18851, signal_18849}), .clk ( clk ), .r ({Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950]}), .c ({signal_6435, signal_6434, signal_6433, signal_6432, signal_1944}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1930 ( .a ({signal_5683, signal_5682, signal_5681, signal_5680, signal_1756}), .b ({signal_5687, signal_5686, signal_5685, signal_5684, signal_1757}), .clk ( clk ), .r ({Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960]}), .c ({signal_6439, signal_6438, signal_6437, signal_6436, signal_1945}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1931 ( .a ({signal_18867, signal_18865, signal_18863, signal_18861, signal_18859}), .b ({signal_5695, signal_5694, signal_5693, signal_5692, signal_1759}), .clk ( clk ), .r ({Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970]}), .c ({signal_6443, signal_6442, signal_6441, signal_6440, signal_1946}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1933 ( .a ({signal_18887, signal_18883, signal_18879, signal_18875, signal_18871}), .b ({signal_5967, signal_5966, signal_5965, signal_5964, signal_1827}), .clk ( clk ), .r ({Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980]}), .c ({signal_6451, signal_6450, signal_6449, signal_6448, signal_1948}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1934 ( .a ({signal_18897, signal_18895, signal_18893, signal_18891, signal_18889}), .b ({signal_5991, signal_5990, signal_5989, signal_5988, signal_1833}), .clk ( clk ), .r ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990]}), .c ({signal_6455, signal_6454, signal_6453, signal_6452, signal_1949}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1935 ( .a ({signal_18907, signal_18905, signal_18903, signal_18901, signal_18899}), .b ({signal_5999, signal_5998, signal_5997, signal_5996, signal_1835}), .clk ( clk ), .r ({Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .c ({signal_6459, signal_6458, signal_6457, signal_6456, signal_1950}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1936 ( .a ({signal_5703, signal_5702, signal_5701, signal_5700, signal_1761}), .b ({signal_6003, signal_6002, signal_6001, signal_6000, signal_1836}), .clk ( clk ), .r ({Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010]}), .c ({signal_6463, signal_6462, signal_6461, signal_6460, signal_1951}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1937 ( .a ({signal_18917, signal_18915, signal_18913, signal_18911, signal_18909}), .b ({signal_5679, signal_5678, signal_5677, signal_5676, signal_1755}), .clk ( clk ), .r ({Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020]}), .c ({signal_6467, signal_6466, signal_6465, signal_6464, signal_1952}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1938 ( .a ({signal_18927, signal_18925, signal_18923, signal_18921, signal_18919}), .b ({signal_6007, signal_6006, signal_6005, signal_6004, signal_1837}), .clk ( clk ), .r ({Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030]}), .c ({signal_6471, signal_6470, signal_6469, signal_6468, signal_1953}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1939 ( .a ({signal_18937, signal_18935, signal_18933, signal_18931, signal_18929}), .b ({signal_6011, signal_6010, signal_6009, signal_6008, signal_1838}), .clk ( clk ), .r ({Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040]}), .c ({signal_6475, signal_6474, signal_6473, signal_6472, signal_1954}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1940 ( .a ({signal_18957, signal_18953, signal_18949, signal_18945, signal_18941}), .b ({signal_6019, signal_6018, signal_6017, signal_6016, signal_1840}), .clk ( clk ), .r ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050]}), .c ({signal_6479, signal_6478, signal_6477, signal_6476, signal_1955}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1941 ( .a ({signal_18967, signal_18965, signal_18963, signal_18961, signal_18959}), .b ({signal_5711, signal_5710, signal_5709, signal_5708, signal_1763}), .clk ( clk ), .r ({Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .c ({signal_6483, signal_6482, signal_6481, signal_6480, signal_1956}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1942 ( .a ({signal_18977, signal_18975, signal_18973, signal_18971, signal_18969}), .b ({signal_6023, signal_6022, signal_6021, signal_6020, signal_1841}), .clk ( clk ), .r ({Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070]}), .c ({signal_6487, signal_6486, signal_6485, signal_6484, signal_1957}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1943 ( .a ({signal_5871, signal_5870, signal_5869, signal_5868, signal_1803}), .b ({signal_18987, signal_18985, signal_18983, signal_18981, signal_18979}), .clk ( clk ), .r ({Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080]}), .c ({signal_6491, signal_6490, signal_6489, signal_6488, signal_1958}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1945 ( .a ({signal_5959, signal_5958, signal_5957, signal_5956, signal_1825}), .b ({signal_6043, signal_6042, signal_6041, signal_6040, signal_1846}), .clk ( clk ), .r ({Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090]}), .c ({signal_6499, signal_6498, signal_6497, signal_6496, signal_1960}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1946 ( .a ({signal_18997, signal_18995, signal_18993, signal_18991, signal_18989}), .b ({signal_5719, signal_5718, signal_5717, signal_5716, signal_1765}), .clk ( clk ), .r ({Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100]}), .c ({signal_6503, signal_6502, signal_6501, signal_6500, signal_1961}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1947 ( .a ({signal_5843, signal_5842, signal_5841, signal_5840, signal_1796}), .b ({signal_6047, signal_6046, signal_6045, signal_6044, signal_1847}), .clk ( clk ), .r ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110]}), .c ({signal_6507, signal_6506, signal_6505, signal_6504, signal_1962}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1961 ( .a ({signal_6291, signal_6290, signal_6289, signal_6288, signal_1908}), .b ({signal_6563, signal_6562, signal_6561, signal_6560, signal_1976}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1969 ( .a ({signal_6327, signal_6326, signal_6325, signal_6324, signal_1917}), .b ({signal_6595, signal_6594, signal_6593, signal_6592, signal_1984}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1971 ( .a ({signal_6335, signal_6334, signal_6333, signal_6332, signal_1919}), .b ({signal_6603, signal_6602, signal_6601, signal_6600, signal_1986}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1978 ( .a ({signal_6367, signal_6366, signal_6365, signal_6364, signal_1927}), .b ({signal_6631, signal_6630, signal_6629, signal_6628, signal_1993}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1986 ( .a ({signal_6403, signal_6402, signal_6401, signal_6400, signal_1936}), .b ({signal_6663, signal_6662, signal_6661, signal_6660, signal_2001}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1987 ( .a ({signal_6407, signal_6406, signal_6405, signal_6404, signal_1937}), .b ({signal_6667, signal_6666, signal_6665, signal_6664, signal_2002}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1989 ( .a ({signal_6415, signal_6414, signal_6413, signal_6412, signal_1939}), .b ({signal_6675, signal_6674, signal_6673, signal_6672, signal_2004}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1992 ( .a ({signal_6455, signal_6454, signal_6453, signal_6452, signal_1949}), .b ({signal_6687, signal_6686, signal_6685, signal_6684, signal_2007}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1993 ( .a ({signal_6463, signal_6462, signal_6461, signal_6460, signal_1951}), .b ({signal_6691, signal_6690, signal_6689, signal_6688, signal_2008}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1994 ( .a ({signal_6487, signal_6486, signal_6485, signal_6484, signal_1957}), .b ({signal_6695, signal_6694, signal_6693, signal_6692, signal_2009}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1995 ( .a ({signal_6491, signal_6490, signal_6489, signal_6488, signal_1958}), .b ({signal_6699, signal_6698, signal_6697, signal_6696, signal_2010}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1997 ( .a ({signal_6499, signal_6498, signal_6497, signal_6496, signal_1960}), .b ({signal_6707, signal_6706, signal_6705, signal_6704, signal_2012}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_1998 ( .a ({signal_6507, signal_6506, signal_6505, signal_6504, signal_1962}), .b ({signal_6711, signal_6710, signal_6709, signal_6708, signal_2013}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_1999 ( .a ({signal_6087, signal_6086, signal_6085, signal_6084, signal_1857}), .b ({signal_19017, signal_19013, signal_19009, signal_19005, signal_19001}), .clk ( clk ), .r ({Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .c ({signal_6715, signal_6714, signal_6713, signal_6712, signal_2014}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2002 ( .a ({signal_19027, signal_19025, signal_19023, signal_19021, signal_19019}), .b ({signal_5755, signal_5754, signal_5753, signal_5752, signal_1774}), .clk ( clk ), .r ({Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130]}), .c ({signal_6727, signal_6726, signal_6725, signal_6724, signal_2017}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2007 ( .a ({signal_19037, signal_19035, signal_19033, signal_19031, signal_19029}), .b ({signal_6235, signal_6234, signal_6233, signal_6232, signal_1894}), .clk ( clk ), .r ({Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140]}), .c ({signal_6747, signal_6746, signal_6745, signal_6744, signal_2022}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2009 ( .a ({signal_19057, signal_19053, signal_19049, signal_19045, signal_19041}), .b ({signal_6243, signal_6242, signal_6241, signal_6240, signal_1896}), .clk ( clk ), .r ({Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150]}), .c ({signal_6755, signal_6754, signal_6753, signal_6752, signal_2024}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2010 ( .a ({signal_19077, signal_19073, signal_19069, signal_19065, signal_19061}), .b ({signal_6255, signal_6254, signal_6253, signal_6252, signal_1899}), .clk ( clk ), .r ({Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160]}), .c ({signal_6759, signal_6758, signal_6757, signal_6756, signal_2025}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2013 ( .a ({signal_19097, signal_19093, signal_19089, signal_19085, signal_19081}), .b ({signal_6131, signal_6130, signal_6129, signal_6128, signal_1868}), .clk ( clk ), .r ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170]}), .c ({signal_6771, signal_6770, signal_6769, signal_6768, signal_2028}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2016 ( .a ({signal_19117, signal_19113, signal_19109, signal_19105, signal_19101}), .b ({signal_6155, signal_6154, signal_6153, signal_6152, signal_1874}), .clk ( clk ), .r ({Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .c ({signal_6783, signal_6782, signal_6781, signal_6780, signal_2031}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2017 ( .a ({signal_19127, signal_19125, signal_19123, signal_19121, signal_19119}), .b ({signal_6159, signal_6158, signal_6157, signal_6156, signal_1875}), .clk ( clk ), .r ({Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190]}), .c ({signal_6787, signal_6786, signal_6785, signal_6784, signal_2032}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2018 ( .a ({signal_19137, signal_19135, signal_19133, signal_19131, signal_19129}), .b ({signal_6163, signal_6162, signal_6161, signal_6160, signal_1876}), .clk ( clk ), .r ({Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200]}), .c ({signal_6791, signal_6790, signal_6789, signal_6788, signal_2033}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2019 ( .a ({signal_19147, signal_19145, signal_19143, signal_19141, signal_19139}), .b ({signal_5911, signal_5910, signal_5909, signal_5908, signal_1813}), .clk ( clk ), .r ({Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210]}), .c ({signal_6795, signal_6794, signal_6793, signal_6792, signal_2034}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2020 ( .a ({signal_19157, signal_19155, signal_19153, signal_19151, signal_19149}), .b ({signal_6167, signal_6166, signal_6165, signal_6164, signal_1877}), .clk ( clk ), .r ({Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220]}), .c ({signal_6799, signal_6798, signal_6797, signal_6796, signal_2035}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2021 ( .a ({signal_19167, signal_19165, signal_19163, signal_19161, signal_19159}), .b ({signal_6171, signal_6170, signal_6169, signal_6168, signal_1878}), .clk ( clk ), .r ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230]}), .c ({signal_6803, signal_6802, signal_6801, signal_6800, signal_2036}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2022 ( .a ({signal_19187, signal_19183, signal_19179, signal_19175, signal_19171}), .b ({signal_6175, signal_6174, signal_6173, signal_6172, signal_1879}), .clk ( clk ), .r ({Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .c ({signal_6807, signal_6806, signal_6805, signal_6804, signal_2037}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2023 ( .a ({signal_19207, signal_19203, signal_19199, signal_19195, signal_19191}), .b ({signal_6179, signal_6178, signal_6177, signal_6176, signal_1880}), .clk ( clk ), .r ({Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250]}), .c ({signal_6811, signal_6810, signal_6809, signal_6808, signal_2038}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2024 ( .a ({signal_19227, signal_19223, signal_19219, signal_19215, signal_19211}), .b ({signal_6183, signal_6182, signal_6181, signal_6180, signal_1881}), .clk ( clk ), .r ({Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260]}), .c ({signal_6815, signal_6814, signal_6813, signal_6812, signal_2039}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2025 ( .a ({signal_19237, signal_19235, signal_19233, signal_19231, signal_19229}), .b ({signal_6187, signal_6186, signal_6185, signal_6184, signal_1882}), .clk ( clk ), .r ({Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270]}), .c ({signal_6819, signal_6818, signal_6817, signal_6816, signal_2040}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2026 ( .a ({signal_5963, signal_5962, signal_5961, signal_5960, signal_1826}), .b ({signal_6323, signal_6322, signal_6321, signal_6320, signal_1916}), .clk ( clk ), .r ({Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280]}), .c ({signal_6823, signal_6822, signal_6821, signal_6820, signal_2041}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2028 ( .a ({signal_19257, signal_19253, signal_19249, signal_19245, signal_19241}), .b ({signal_6191, signal_6190, signal_6189, signal_6188, signal_1883}), .clk ( clk ), .r ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290]}), .c ({signal_6831, signal_6830, signal_6829, signal_6828, signal_2043}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2029 ( .a ({signal_19267, signal_19265, signal_19263, signal_19261, signal_19259}), .b ({signal_6195, signal_6194, signal_6193, signal_6192, signal_1884}), .clk ( clk ), .r ({Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .c ({signal_6835, signal_6834, signal_6833, signal_6832, signal_2044}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2030 ( .a ({signal_19277, signal_19275, signal_19273, signal_19271, signal_19269}), .b ({signal_5979, signal_5978, signal_5977, signal_5976, signal_1830}), .clk ( clk ), .r ({Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310]}), .c ({signal_6839, signal_6838, signal_6837, signal_6836, signal_2045}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2031 ( .a ({signal_19287, signal_19285, signal_19283, signal_19281, signal_19279}), .b ({signal_6203, signal_6202, signal_6201, signal_6200, signal_1886}), .clk ( clk ), .r ({Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320]}), .c ({signal_6843, signal_6842, signal_6841, signal_6840, signal_2046}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2033 ( .a ({signal_19297, signal_19295, signal_19293, signal_19291, signal_19289}), .b ({signal_6015, signal_6014, signal_6013, signal_6012, signal_1839}), .clk ( clk ), .r ({Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330]}), .c ({signal_6851, signal_6850, signal_6849, signal_6848, signal_2048}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2034 ( .a ({signal_19307, signal_19305, signal_19303, signal_19301, signal_19299}), .b ({signal_5931, signal_5930, signal_5929, signal_5928, signal_1818}), .clk ( clk ), .r ({Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340]}), .c ({signal_6855, signal_6854, signal_6853, signal_6852, signal_2049}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2035 ( .a ({signal_19327, signal_19323, signal_19319, signal_19315, signal_19311}), .b ({signal_6211, signal_6210, signal_6209, signal_6208, signal_1888}), .clk ( clk ), .r ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350]}), .c ({signal_6859, signal_6858, signal_6857, signal_6856, signal_2050}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2036 ( .a ({signal_19057, signal_19053, signal_19049, signal_19045, signal_19041}), .b ({signal_6215, signal_6214, signal_6213, signal_6212, signal_1889}), .clk ( clk ), .r ({Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .c ({signal_6863, signal_6862, signal_6861, signal_6860, signal_2051}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2046 ( .a ({signal_6715, signal_6714, signal_6713, signal_6712, signal_2014}), .b ({signal_6903, signal_6902, signal_6901, signal_6900, signal_2061}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2047 ( .a ({signal_6727, signal_6726, signal_6725, signal_6724, signal_2017}), .b ({signal_6907, signal_6906, signal_6905, signal_6904, signal_2062}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2049 ( .a ({signal_6747, signal_6746, signal_6745, signal_6744, signal_2022}), .b ({signal_6915, signal_6914, signal_6913, signal_6912, signal_2064}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2050 ( .a ({signal_6755, signal_6754, signal_6753, signal_6752, signal_2024}), .b ({signal_6919, signal_6918, signal_6917, signal_6916, signal_2065}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2051 ( .a ({signal_6759, signal_6758, signal_6757, signal_6756, signal_2025}), .b ({signal_6923, signal_6922, signal_6921, signal_6920, signal_2066}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2053 ( .a ({signal_6771, signal_6770, signal_6769, signal_6768, signal_2028}), .b ({signal_6931, signal_6930, signal_6929, signal_6928, signal_2068}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2054 ( .a ({signal_6783, signal_6782, signal_6781, signal_6780, signal_2031}), .b ({signal_6935, signal_6934, signal_6933, signal_6932, signal_2069}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2055 ( .a ({signal_6787, signal_6786, signal_6785, signal_6784, signal_2032}), .b ({signal_6939, signal_6938, signal_6937, signal_6936, signal_2070}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2056 ( .a ({signal_6791, signal_6790, signal_6789, signal_6788, signal_2033}), .b ({signal_6943, signal_6942, signal_6941, signal_6940, signal_2071}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2057 ( .a ({signal_6795, signal_6794, signal_6793, signal_6792, signal_2034}), .b ({signal_6947, signal_6946, signal_6945, signal_6944, signal_2072}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2058 ( .a ({signal_6799, signal_6798, signal_6797, signal_6796, signal_2035}), .b ({signal_6951, signal_6950, signal_6949, signal_6948, signal_2073}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2059 ( .a ({signal_6803, signal_6802, signal_6801, signal_6800, signal_2036}), .b ({signal_6955, signal_6954, signal_6953, signal_6952, signal_2074}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2060 ( .a ({signal_6807, signal_6806, signal_6805, signal_6804, signal_2037}), .b ({signal_6959, signal_6958, signal_6957, signal_6956, signal_2075}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2061 ( .a ({signal_6811, signal_6810, signal_6809, signal_6808, signal_2038}), .b ({signal_6963, signal_6962, signal_6961, signal_6960, signal_2076}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2062 ( .a ({signal_6815, signal_6814, signal_6813, signal_6812, signal_2039}), .b ({signal_6967, signal_6966, signal_6965, signal_6964, signal_2077}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2063 ( .a ({signal_6823, signal_6822, signal_6821, signal_6820, signal_2041}), .b ({signal_6971, signal_6970, signal_6969, signal_6968, signal_2078}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2065 ( .a ({signal_6831, signal_6830, signal_6829, signal_6828, signal_2043}), .b ({signal_6979, signal_6978, signal_6977, signal_6976, signal_2080}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2066 ( .a ({signal_6835, signal_6834, signal_6833, signal_6832, signal_2044}), .b ({signal_6983, signal_6982, signal_6981, signal_6980, signal_2081}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2067 ( .a ({signal_6843, signal_6842, signal_6841, signal_6840, signal_2046}), .b ({signal_6987, signal_6986, signal_6985, signal_6984, signal_2082}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2069 ( .a ({signal_6851, signal_6850, signal_6849, signal_6848, signal_2048}), .b ({signal_6995, signal_6994, signal_6993, signal_6992, signal_2084}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2070 ( .a ({signal_6859, signal_6858, signal_6857, signal_6856, signal_2050}), .b ({signal_6999, signal_6998, signal_6997, signal_6996, signal_2085}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2071 ( .a ({signal_6863, signal_6862, signal_6861, signal_6860, signal_2051}), .b ({signal_7003, signal_7002, signal_7001, signal_7000, signal_2086}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2074 ( .a ({signal_6567, signal_6566, signal_6565, signal_6564, signal_1977}), .b ({signal_19347, signal_19343, signal_19339, signal_19335, signal_19331}), .clk ( clk ), .r ({Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370]}), .c ({signal_7015, signal_7014, signal_7013, signal_7012, signal_2089}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2075 ( .a ({signal_19357, signal_19355, signal_19353, signal_19351, signal_19349}), .b ({signal_6515, signal_6514, signal_6513, signal_6512, signal_1964}), .clk ( clk ), .r ({Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380]}), .c ({signal_7019, signal_7018, signal_7017, signal_7016, signal_2090}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2076 ( .a ({signal_19377, signal_19373, signal_19369, signal_19365, signal_19361}), .b ({signal_6719, signal_6718, signal_6717, signal_6716, signal_2015}), .clk ( clk ), .r ({Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390]}), .c ({signal_7023, signal_7022, signal_7021, signal_7020, signal_2091}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2077 ( .a ({signal_19387, signal_19385, signal_19383, signal_19381, signal_19379}), .b ({signal_6535, signal_6534, signal_6533, signal_6532, signal_1969}), .clk ( clk ), .r ({Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400]}), .c ({signal_7027, signal_7026, signal_7025, signal_7024, signal_2092}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2078 ( .a ({signal_6511, signal_6510, signal_6509, signal_6508, signal_1963}), .b ({signal_19397, signal_19395, signal_19393, signal_19391, signal_19389}), .clk ( clk ), .r ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410]}), .c ({signal_7031, signal_7030, signal_7029, signal_7028, signal_2093}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2079 ( .a ({signal_6551, signal_6550, signal_6549, signal_6548, signal_1973}), .b ({signal_6555, signal_6554, signal_6553, signal_6552, signal_1974}), .clk ( clk ), .r ({Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .c ({signal_7035, signal_7034, signal_7033, signal_7032, signal_2094}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2080 ( .a ({signal_19417, signal_19413, signal_19409, signal_19405, signal_19401}), .b ({signal_6731, signal_6730, signal_6729, signal_6728, signal_2018}), .clk ( clk ), .r ({Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430]}), .c ({signal_7039, signal_7038, signal_7037, signal_7036, signal_2095}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2081 ( .a ({signal_19437, signal_19433, signal_19429, signal_19425, signal_19421}), .b ({signal_6739, signal_6738, signal_6737, signal_6736, signal_2020}), .clk ( clk ), .r ({Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440]}), .c ({signal_7043, signal_7042, signal_7041, signal_7040, signal_2096}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2082 ( .a ({signal_19457, signal_19453, signal_19449, signal_19445, signal_19441}), .b ({signal_6743, signal_6742, signal_6741, signal_6740, signal_2021}), .clk ( clk ), .r ({Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450]}), .c ({signal_7047, signal_7046, signal_7045, signal_7044, signal_2097}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2083 ( .a ({signal_19467, signal_19465, signal_19463, signal_19461, signal_19459}), .b ({signal_6583, signal_6582, signal_6581, signal_6580, signal_1981}), .clk ( clk ), .r ({Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460]}), .c ({signal_7051, signal_7050, signal_7049, signal_7048, signal_2098}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2085 ( .a ({signal_19487, signal_19483, signal_19479, signal_19475, signal_19471}), .b ({signal_6599, signal_6598, signal_6597, signal_6596, signal_1985}), .clk ( clk ), .r ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470]}), .c ({signal_7059, signal_7058, signal_7057, signal_7056, signal_2100}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2086 ( .a ({signal_19507, signal_19503, signal_19499, signal_19495, signal_19491}), .b ({signal_6751, signal_6750, signal_6749, signal_6748, signal_2023}), .clk ( clk ), .r ({Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .c ({signal_7063, signal_7062, signal_7061, signal_7060, signal_2101}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2087 ( .a ({signal_6223, signal_6222, signal_6221, signal_6220, signal_1891}), .b ({signal_6615, signal_6614, signal_6613, signal_6612, signal_1989}), .clk ( clk ), .r ({Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490]}), .c ({signal_7067, signal_7066, signal_7065, signal_7064, signal_2102}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2088 ( .a ({signal_6619, signal_6618, signal_6617, signal_6616, signal_1990}), .b ({signal_6623, signal_6622, signal_6621, signal_6620, signal_1991}), .clk ( clk ), .r ({Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500]}), .c ({signal_7071, signal_7070, signal_7069, signal_7068, signal_2103}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2089 ( .a ({signal_19517, signal_19515, signal_19513, signal_19511, signal_19509}), .b ({signal_6627, signal_6626, signal_6625, signal_6624, signal_1992}), .clk ( clk ), .r ({Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510]}), .c ({signal_7075, signal_7074, signal_7073, signal_7072, signal_2104}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2091 ( .a ({signal_6767, signal_6766, signal_6765, signal_6764, signal_2027}), .b ({signal_6199, signal_6198, signal_6197, signal_6196, signal_1885}), .clk ( clk ), .r ({Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520]}), .c ({signal_7083, signal_7082, signal_7081, signal_7080, signal_2106}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2092 ( .a ({signal_19537, signal_19533, signal_19529, signal_19525, signal_19521}), .b ({signal_6635, signal_6634, signal_6633, signal_6632, signal_1994}), .clk ( clk ), .r ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530]}), .c ({signal_7087, signal_7086, signal_7085, signal_7084, signal_2107}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2093 ( .a ({signal_19547, signal_19545, signal_19543, signal_19541, signal_19539}), .b ({signal_6639, signal_6638, signal_6637, signal_6636, signal_1995}), .clk ( clk ), .r ({Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .c ({signal_7091, signal_7090, signal_7089, signal_7088, signal_2108}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2094 ( .a ({signal_5867, signal_5866, signal_5865, signal_5864, signal_1802}), .b ({signal_6643, signal_6642, signal_6641, signal_6640, signal_1996}), .clk ( clk ), .r ({Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550]}), .c ({signal_7095, signal_7094, signal_7093, signal_7092, signal_2109}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2095 ( .a ({signal_6543, signal_6542, signal_6541, signal_6540, signal_1971}), .b ({signal_6647, signal_6646, signal_6645, signal_6644, signal_1997}), .clk ( clk ), .r ({Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560]}), .c ({signal_7099, signal_7098, signal_7097, signal_7096, signal_2110}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2096 ( .a ({signal_5683, signal_5682, signal_5681, signal_5680, signal_1756}), .b ({signal_6651, signal_6650, signal_6649, signal_6648, signal_1998}), .clk ( clk ), .r ({Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570]}), .c ({signal_7103, signal_7102, signal_7101, signal_7100, signal_2111}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2097 ( .a ({signal_6547, signal_6546, signal_6545, signal_6544, signal_1972}), .b ({signal_18857, signal_18855, signal_18853, signal_18851, signal_18849}), .clk ( clk ), .r ({Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580]}), .c ({signal_7107, signal_7106, signal_7105, signal_7104, signal_2112}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2099 ( .a ({signal_5451, signal_5450, signal_5449, signal_5448, signal_1698}), .b ({signal_6659, signal_6658, signal_6657, signal_6656, signal_2000}), .clk ( clk ), .r ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590]}), .c ({signal_7115, signal_7114, signal_7113, signal_7112, signal_2114}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2101 ( .a ({signal_6559, signal_6558, signal_6557, signal_6556, signal_1975}), .b ({signal_6671, signal_6670, signal_6669, signal_6668, signal_2003}), .clk ( clk ), .r ({Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .c ({signal_7123, signal_7122, signal_7121, signal_7120, signal_2116}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2104 ( .a ({signal_19557, signal_19555, signal_19553, signal_19551, signal_19549}), .b ({signal_6679, signal_6678, signal_6677, signal_6676, signal_2005}), .clk ( clk ), .r ({Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610]}), .c ({signal_7135, signal_7134, signal_7133, signal_7132, signal_2119}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2110 ( .a ({signal_6775, signal_6774, signal_6773, signal_6772, signal_2029}), .b ({signal_6051, signal_6050, signal_6049, signal_6048, signal_1848}), .clk ( clk ), .r ({Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620]}), .c ({signal_7159, signal_7158, signal_7157, signal_7156, signal_2125}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2124 ( .a ({signal_7015, signal_7014, signal_7013, signal_7012, signal_2089}), .b ({signal_7215, signal_7214, signal_7213, signal_7212, signal_2139}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2125 ( .a ({signal_7023, signal_7022, signal_7021, signal_7020, signal_2091}), .b ({signal_7219, signal_7218, signal_7217, signal_7216, signal_2140}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2126 ( .a ({signal_7027, signal_7026, signal_7025, signal_7024, signal_2092}), .b ({signal_7223, signal_7222, signal_7221, signal_7220, signal_2141}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2127 ( .a ({signal_7043, signal_7042, signal_7041, signal_7040, signal_2096}), .b ({signal_7227, signal_7226, signal_7225, signal_7224, signal_2142}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2128 ( .a ({signal_7047, signal_7046, signal_7045, signal_7044, signal_2097}), .b ({signal_7231, signal_7230, signal_7229, signal_7228, signal_2143}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2130 ( .a ({signal_7063, signal_7062, signal_7061, signal_7060, signal_2101}), .b ({signal_7239, signal_7238, signal_7237, signal_7236, signal_2145}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2133 ( .a ({signal_7135, signal_7134, signal_7133, signal_7132, signal_2119}), .b ({signal_7251, signal_7250, signal_7249, signal_7248, signal_2148}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2135 ( .a ({signal_7159, signal_7158, signal_7157, signal_7156, signal_2125}), .b ({signal_7259, signal_7258, signal_7257, signal_7256, signal_2150}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2144 ( .a ({signal_19567, signal_19565, signal_19563, signal_19561, signal_19559}), .b ({signal_6911, signal_6910, signal_6909, signal_6908, signal_2063}), .clk ( clk ), .r ({Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630]}), .c ({signal_7295, signal_7294, signal_7293, signal_7292, signal_2159}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2148 ( .a ({signal_19587, signal_19583, signal_19579, signal_19575, signal_19571}), .b ({signal_6927, signal_6926, signal_6925, signal_6924, signal_2067}), .clk ( clk ), .r ({Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640]}), .c ({signal_7311, signal_7310, signal_7309, signal_7308, signal_2163}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2185 ( .a ({signal_7295, signal_7294, signal_7293, signal_7292, signal_2159}), .b ({signal_7459, signal_7458, signal_7457, signal_7456, signal_2200}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2186 ( .a ({signal_7311, signal_7310, signal_7309, signal_7308, signal_2163}), .b ({signal_7463, signal_7462, signal_7461, signal_7460, signal_2201}) ) ;
    buf_clk cell_4896 ( .C ( clk ), .D ( signal_19588 ), .Q ( signal_19589 ) ) ;
    buf_clk cell_4898 ( .C ( clk ), .D ( signal_19590 ), .Q ( signal_19591 ) ) ;
    buf_clk cell_4900 ( .C ( clk ), .D ( signal_19592 ), .Q ( signal_19593 ) ) ;
    buf_clk cell_4902 ( .C ( clk ), .D ( signal_19594 ), .Q ( signal_19595 ) ) ;
    buf_clk cell_4904 ( .C ( clk ), .D ( signal_19596 ), .Q ( signal_19597 ) ) ;
    buf_clk cell_4910 ( .C ( clk ), .D ( signal_19602 ), .Q ( signal_19603 ) ) ;
    buf_clk cell_4916 ( .C ( clk ), .D ( signal_19608 ), .Q ( signal_19609 ) ) ;
    buf_clk cell_4922 ( .C ( clk ), .D ( signal_19614 ), .Q ( signal_19615 ) ) ;
    buf_clk cell_4928 ( .C ( clk ), .D ( signal_19620 ), .Q ( signal_19621 ) ) ;
    buf_clk cell_4934 ( .C ( clk ), .D ( signal_19626 ), .Q ( signal_19627 ) ) ;
    buf_clk cell_4940 ( .C ( clk ), .D ( signal_19632 ), .Q ( signal_19633 ) ) ;
    buf_clk cell_4946 ( .C ( clk ), .D ( signal_19638 ), .Q ( signal_19639 ) ) ;
    buf_clk cell_4952 ( .C ( clk ), .D ( signal_19644 ), .Q ( signal_19645 ) ) ;
    buf_clk cell_4958 ( .C ( clk ), .D ( signal_19650 ), .Q ( signal_19651 ) ) ;
    buf_clk cell_4964 ( .C ( clk ), .D ( signal_19656 ), .Q ( signal_19657 ) ) ;
    buf_clk cell_4970 ( .C ( clk ), .D ( signal_19662 ), .Q ( signal_19663 ) ) ;
    buf_clk cell_4976 ( .C ( clk ), .D ( signal_19668 ), .Q ( signal_19669 ) ) ;
    buf_clk cell_4982 ( .C ( clk ), .D ( signal_19674 ), .Q ( signal_19675 ) ) ;
    buf_clk cell_4988 ( .C ( clk ), .D ( signal_19680 ), .Q ( signal_19681 ) ) ;
    buf_clk cell_4994 ( .C ( clk ), .D ( signal_19686 ), .Q ( signal_19687 ) ) ;
    buf_clk cell_4998 ( .C ( clk ), .D ( signal_19690 ), .Q ( signal_19691 ) ) ;
    buf_clk cell_5002 ( .C ( clk ), .D ( signal_19694 ), .Q ( signal_19695 ) ) ;
    buf_clk cell_5006 ( .C ( clk ), .D ( signal_19698 ), .Q ( signal_19699 ) ) ;
    buf_clk cell_5010 ( .C ( clk ), .D ( signal_19702 ), .Q ( signal_19703 ) ) ;
    buf_clk cell_5014 ( .C ( clk ), .D ( signal_19706 ), .Q ( signal_19707 ) ) ;
    buf_clk cell_5020 ( .C ( clk ), .D ( signal_19712 ), .Q ( signal_19713 ) ) ;
    buf_clk cell_5026 ( .C ( clk ), .D ( signal_19718 ), .Q ( signal_19719 ) ) ;
    buf_clk cell_5032 ( .C ( clk ), .D ( signal_19724 ), .Q ( signal_19725 ) ) ;
    buf_clk cell_5038 ( .C ( clk ), .D ( signal_19730 ), .Q ( signal_19731 ) ) ;
    buf_clk cell_5044 ( .C ( clk ), .D ( signal_19736 ), .Q ( signal_19737 ) ) ;
    buf_clk cell_5048 ( .C ( clk ), .D ( signal_19740 ), .Q ( signal_19741 ) ) ;
    buf_clk cell_5052 ( .C ( clk ), .D ( signal_19744 ), .Q ( signal_19745 ) ) ;
    buf_clk cell_5056 ( .C ( clk ), .D ( signal_19748 ), .Q ( signal_19749 ) ) ;
    buf_clk cell_5060 ( .C ( clk ), .D ( signal_19752 ), .Q ( signal_19753 ) ) ;
    buf_clk cell_5064 ( .C ( clk ), .D ( signal_19756 ), .Q ( signal_19757 ) ) ;
    buf_clk cell_5068 ( .C ( clk ), .D ( signal_19760 ), .Q ( signal_19761 ) ) ;
    buf_clk cell_5072 ( .C ( clk ), .D ( signal_19764 ), .Q ( signal_19765 ) ) ;
    buf_clk cell_5076 ( .C ( clk ), .D ( signal_19768 ), .Q ( signal_19769 ) ) ;
    buf_clk cell_5080 ( .C ( clk ), .D ( signal_19772 ), .Q ( signal_19773 ) ) ;
    buf_clk cell_5084 ( .C ( clk ), .D ( signal_19776 ), .Q ( signal_19777 ) ) ;
    buf_clk cell_5088 ( .C ( clk ), .D ( signal_19780 ), .Q ( signal_19781 ) ) ;
    buf_clk cell_5092 ( .C ( clk ), .D ( signal_19784 ), .Q ( signal_19785 ) ) ;
    buf_clk cell_5096 ( .C ( clk ), .D ( signal_19788 ), .Q ( signal_19789 ) ) ;
    buf_clk cell_5100 ( .C ( clk ), .D ( signal_19792 ), .Q ( signal_19793 ) ) ;
    buf_clk cell_5104 ( .C ( clk ), .D ( signal_19796 ), .Q ( signal_19797 ) ) ;
    buf_clk cell_5108 ( .C ( clk ), .D ( signal_19800 ), .Q ( signal_19801 ) ) ;
    buf_clk cell_5112 ( .C ( clk ), .D ( signal_19804 ), .Q ( signal_19805 ) ) ;
    buf_clk cell_5116 ( .C ( clk ), .D ( signal_19808 ), .Q ( signal_19809 ) ) ;
    buf_clk cell_5120 ( .C ( clk ), .D ( signal_19812 ), .Q ( signal_19813 ) ) ;
    buf_clk cell_5124 ( .C ( clk ), .D ( signal_19816 ), .Q ( signal_19817 ) ) ;
    buf_clk cell_5128 ( .C ( clk ), .D ( signal_19820 ), .Q ( signal_19821 ) ) ;
    buf_clk cell_5132 ( .C ( clk ), .D ( signal_19824 ), .Q ( signal_19825 ) ) ;
    buf_clk cell_5136 ( .C ( clk ), .D ( signal_19828 ), .Q ( signal_19829 ) ) ;
    buf_clk cell_5140 ( .C ( clk ), .D ( signal_19832 ), .Q ( signal_19833 ) ) ;
    buf_clk cell_5144 ( .C ( clk ), .D ( signal_19836 ), .Q ( signal_19837 ) ) ;
    buf_clk cell_5150 ( .C ( clk ), .D ( signal_19842 ), .Q ( signal_19843 ) ) ;
    buf_clk cell_5156 ( .C ( clk ), .D ( signal_19848 ), .Q ( signal_19849 ) ) ;
    buf_clk cell_5162 ( .C ( clk ), .D ( signal_19854 ), .Q ( signal_19855 ) ) ;
    buf_clk cell_5168 ( .C ( clk ), .D ( signal_19860 ), .Q ( signal_19861 ) ) ;
    buf_clk cell_5174 ( .C ( clk ), .D ( signal_19866 ), .Q ( signal_19867 ) ) ;
    buf_clk cell_5178 ( .C ( clk ), .D ( signal_19870 ), .Q ( signal_19871 ) ) ;
    buf_clk cell_5182 ( .C ( clk ), .D ( signal_19874 ), .Q ( signal_19875 ) ) ;
    buf_clk cell_5186 ( .C ( clk ), .D ( signal_19878 ), .Q ( signal_19879 ) ) ;
    buf_clk cell_5190 ( .C ( clk ), .D ( signal_19882 ), .Q ( signal_19883 ) ) ;
    buf_clk cell_5194 ( .C ( clk ), .D ( signal_19886 ), .Q ( signal_19887 ) ) ;
    buf_clk cell_5196 ( .C ( clk ), .D ( signal_19888 ), .Q ( signal_19889 ) ) ;
    buf_clk cell_5198 ( .C ( clk ), .D ( signal_19890 ), .Q ( signal_19891 ) ) ;
    buf_clk cell_5200 ( .C ( clk ), .D ( signal_19892 ), .Q ( signal_19893 ) ) ;
    buf_clk cell_5202 ( .C ( clk ), .D ( signal_19894 ), .Q ( signal_19895 ) ) ;
    buf_clk cell_5204 ( .C ( clk ), .D ( signal_19896 ), .Q ( signal_19897 ) ) ;
    buf_clk cell_5206 ( .C ( clk ), .D ( signal_19898 ), .Q ( signal_19899 ) ) ;
    buf_clk cell_5208 ( .C ( clk ), .D ( signal_19900 ), .Q ( signal_19901 ) ) ;
    buf_clk cell_5210 ( .C ( clk ), .D ( signal_19902 ), .Q ( signal_19903 ) ) ;
    buf_clk cell_5212 ( .C ( clk ), .D ( signal_19904 ), .Q ( signal_19905 ) ) ;
    buf_clk cell_5214 ( .C ( clk ), .D ( signal_19906 ), .Q ( signal_19907 ) ) ;
    buf_clk cell_5216 ( .C ( clk ), .D ( signal_19908 ), .Q ( signal_19909 ) ) ;
    buf_clk cell_5218 ( .C ( clk ), .D ( signal_19910 ), .Q ( signal_19911 ) ) ;
    buf_clk cell_5220 ( .C ( clk ), .D ( signal_19912 ), .Q ( signal_19913 ) ) ;
    buf_clk cell_5222 ( .C ( clk ), .D ( signal_19914 ), .Q ( signal_19915 ) ) ;
    buf_clk cell_5224 ( .C ( clk ), .D ( signal_19916 ), .Q ( signal_19917 ) ) ;
    buf_clk cell_5226 ( .C ( clk ), .D ( signal_19918 ), .Q ( signal_19919 ) ) ;
    buf_clk cell_5228 ( .C ( clk ), .D ( signal_19920 ), .Q ( signal_19921 ) ) ;
    buf_clk cell_5230 ( .C ( clk ), .D ( signal_19922 ), .Q ( signal_19923 ) ) ;
    buf_clk cell_5232 ( .C ( clk ), .D ( signal_19924 ), .Q ( signal_19925 ) ) ;
    buf_clk cell_5234 ( .C ( clk ), .D ( signal_19926 ), .Q ( signal_19927 ) ) ;
    buf_clk cell_5236 ( .C ( clk ), .D ( signal_19928 ), .Q ( signal_19929 ) ) ;
    buf_clk cell_5238 ( .C ( clk ), .D ( signal_19930 ), .Q ( signal_19931 ) ) ;
    buf_clk cell_5240 ( .C ( clk ), .D ( signal_19932 ), .Q ( signal_19933 ) ) ;
    buf_clk cell_5242 ( .C ( clk ), .D ( signal_19934 ), .Q ( signal_19935 ) ) ;
    buf_clk cell_5244 ( .C ( clk ), .D ( signal_19936 ), .Q ( signal_19937 ) ) ;
    buf_clk cell_5248 ( .C ( clk ), .D ( signal_19940 ), .Q ( signal_19941 ) ) ;
    buf_clk cell_5252 ( .C ( clk ), .D ( signal_19944 ), .Q ( signal_19945 ) ) ;
    buf_clk cell_5256 ( .C ( clk ), .D ( signal_19948 ), .Q ( signal_19949 ) ) ;
    buf_clk cell_5260 ( .C ( clk ), .D ( signal_19952 ), .Q ( signal_19953 ) ) ;
    buf_clk cell_5264 ( .C ( clk ), .D ( signal_19956 ), .Q ( signal_19957 ) ) ;
    buf_clk cell_5266 ( .C ( clk ), .D ( signal_19958 ), .Q ( signal_19959 ) ) ;
    buf_clk cell_5268 ( .C ( clk ), .D ( signal_19960 ), .Q ( signal_19961 ) ) ;
    buf_clk cell_5270 ( .C ( clk ), .D ( signal_19962 ), .Q ( signal_19963 ) ) ;
    buf_clk cell_5272 ( .C ( clk ), .D ( signal_19964 ), .Q ( signal_19965 ) ) ;
    buf_clk cell_5274 ( .C ( clk ), .D ( signal_19966 ), .Q ( signal_19967 ) ) ;
    buf_clk cell_5276 ( .C ( clk ), .D ( signal_19968 ), .Q ( signal_19969 ) ) ;
    buf_clk cell_5278 ( .C ( clk ), .D ( signal_19970 ), .Q ( signal_19971 ) ) ;
    buf_clk cell_5280 ( .C ( clk ), .D ( signal_19972 ), .Q ( signal_19973 ) ) ;
    buf_clk cell_5282 ( .C ( clk ), .D ( signal_19974 ), .Q ( signal_19975 ) ) ;
    buf_clk cell_5284 ( .C ( clk ), .D ( signal_19976 ), .Q ( signal_19977 ) ) ;
    buf_clk cell_5286 ( .C ( clk ), .D ( signal_19978 ), .Q ( signal_19979 ) ) ;
    buf_clk cell_5288 ( .C ( clk ), .D ( signal_19980 ), .Q ( signal_19981 ) ) ;
    buf_clk cell_5290 ( .C ( clk ), .D ( signal_19982 ), .Q ( signal_19983 ) ) ;
    buf_clk cell_5292 ( .C ( clk ), .D ( signal_19984 ), .Q ( signal_19985 ) ) ;
    buf_clk cell_5294 ( .C ( clk ), .D ( signal_19986 ), .Q ( signal_19987 ) ) ;
    buf_clk cell_5300 ( .C ( clk ), .D ( signal_19992 ), .Q ( signal_19993 ) ) ;
    buf_clk cell_5306 ( .C ( clk ), .D ( signal_19998 ), .Q ( signal_19999 ) ) ;
    buf_clk cell_5312 ( .C ( clk ), .D ( signal_20004 ), .Q ( signal_20005 ) ) ;
    buf_clk cell_5318 ( .C ( clk ), .D ( signal_20010 ), .Q ( signal_20011 ) ) ;
    buf_clk cell_5324 ( .C ( clk ), .D ( signal_20016 ), .Q ( signal_20017 ) ) ;
    buf_clk cell_5326 ( .C ( clk ), .D ( signal_20018 ), .Q ( signal_20019 ) ) ;
    buf_clk cell_5328 ( .C ( clk ), .D ( signal_20020 ), .Q ( signal_20021 ) ) ;
    buf_clk cell_5330 ( .C ( clk ), .D ( signal_20022 ), .Q ( signal_20023 ) ) ;
    buf_clk cell_5332 ( .C ( clk ), .D ( signal_20024 ), .Q ( signal_20025 ) ) ;
    buf_clk cell_5334 ( .C ( clk ), .D ( signal_20026 ), .Q ( signal_20027 ) ) ;
    buf_clk cell_5338 ( .C ( clk ), .D ( signal_20030 ), .Q ( signal_20031 ) ) ;
    buf_clk cell_5342 ( .C ( clk ), .D ( signal_20034 ), .Q ( signal_20035 ) ) ;
    buf_clk cell_5346 ( .C ( clk ), .D ( signal_20038 ), .Q ( signal_20039 ) ) ;
    buf_clk cell_5350 ( .C ( clk ), .D ( signal_20042 ), .Q ( signal_20043 ) ) ;
    buf_clk cell_5354 ( .C ( clk ), .D ( signal_20046 ), .Q ( signal_20047 ) ) ;
    buf_clk cell_5356 ( .C ( clk ), .D ( signal_20048 ), .Q ( signal_20049 ) ) ;
    buf_clk cell_5358 ( .C ( clk ), .D ( signal_20050 ), .Q ( signal_20051 ) ) ;
    buf_clk cell_5360 ( .C ( clk ), .D ( signal_20052 ), .Q ( signal_20053 ) ) ;
    buf_clk cell_5362 ( .C ( clk ), .D ( signal_20054 ), .Q ( signal_20055 ) ) ;
    buf_clk cell_5364 ( .C ( clk ), .D ( signal_20056 ), .Q ( signal_20057 ) ) ;
    buf_clk cell_5366 ( .C ( clk ), .D ( signal_20058 ), .Q ( signal_20059 ) ) ;
    buf_clk cell_5368 ( .C ( clk ), .D ( signal_20060 ), .Q ( signal_20061 ) ) ;
    buf_clk cell_5370 ( .C ( clk ), .D ( signal_20062 ), .Q ( signal_20063 ) ) ;
    buf_clk cell_5372 ( .C ( clk ), .D ( signal_20064 ), .Q ( signal_20065 ) ) ;
    buf_clk cell_5374 ( .C ( clk ), .D ( signal_20066 ), .Q ( signal_20067 ) ) ;
    buf_clk cell_5380 ( .C ( clk ), .D ( signal_20072 ), .Q ( signal_20073 ) ) ;
    buf_clk cell_5386 ( .C ( clk ), .D ( signal_20078 ), .Q ( signal_20079 ) ) ;
    buf_clk cell_5392 ( .C ( clk ), .D ( signal_20084 ), .Q ( signal_20085 ) ) ;
    buf_clk cell_5398 ( .C ( clk ), .D ( signal_20090 ), .Q ( signal_20091 ) ) ;
    buf_clk cell_5404 ( .C ( clk ), .D ( signal_20096 ), .Q ( signal_20097 ) ) ;
    buf_clk cell_5408 ( .C ( clk ), .D ( signal_20100 ), .Q ( signal_20101 ) ) ;
    buf_clk cell_5412 ( .C ( clk ), .D ( signal_20104 ), .Q ( signal_20105 ) ) ;
    buf_clk cell_5416 ( .C ( clk ), .D ( signal_20108 ), .Q ( signal_20109 ) ) ;
    buf_clk cell_5420 ( .C ( clk ), .D ( signal_20112 ), .Q ( signal_20113 ) ) ;
    buf_clk cell_5424 ( .C ( clk ), .D ( signal_20116 ), .Q ( signal_20117 ) ) ;
    buf_clk cell_5426 ( .C ( clk ), .D ( signal_20118 ), .Q ( signal_20119 ) ) ;
    buf_clk cell_5428 ( .C ( clk ), .D ( signal_20120 ), .Q ( signal_20121 ) ) ;
    buf_clk cell_5430 ( .C ( clk ), .D ( signal_20122 ), .Q ( signal_20123 ) ) ;
    buf_clk cell_5432 ( .C ( clk ), .D ( signal_20124 ), .Q ( signal_20125 ) ) ;
    buf_clk cell_5434 ( .C ( clk ), .D ( signal_20126 ), .Q ( signal_20127 ) ) ;
    buf_clk cell_5436 ( .C ( clk ), .D ( signal_20128 ), .Q ( signal_20129 ) ) ;
    buf_clk cell_5438 ( .C ( clk ), .D ( signal_20130 ), .Q ( signal_20131 ) ) ;
    buf_clk cell_5440 ( .C ( clk ), .D ( signal_20132 ), .Q ( signal_20133 ) ) ;
    buf_clk cell_5442 ( .C ( clk ), .D ( signal_20134 ), .Q ( signal_20135 ) ) ;
    buf_clk cell_5444 ( .C ( clk ), .D ( signal_20136 ), .Q ( signal_20137 ) ) ;
    buf_clk cell_5448 ( .C ( clk ), .D ( signal_20140 ), .Q ( signal_20141 ) ) ;
    buf_clk cell_5452 ( .C ( clk ), .D ( signal_20144 ), .Q ( signal_20145 ) ) ;
    buf_clk cell_5456 ( .C ( clk ), .D ( signal_20148 ), .Q ( signal_20149 ) ) ;
    buf_clk cell_5460 ( .C ( clk ), .D ( signal_20152 ), .Q ( signal_20153 ) ) ;
    buf_clk cell_5464 ( .C ( clk ), .D ( signal_20156 ), .Q ( signal_20157 ) ) ;
    buf_clk cell_5468 ( .C ( clk ), .D ( signal_20160 ), .Q ( signal_20161 ) ) ;
    buf_clk cell_5472 ( .C ( clk ), .D ( signal_20164 ), .Q ( signal_20165 ) ) ;
    buf_clk cell_5476 ( .C ( clk ), .D ( signal_20168 ), .Q ( signal_20169 ) ) ;
    buf_clk cell_5480 ( .C ( clk ), .D ( signal_20172 ), .Q ( signal_20173 ) ) ;
    buf_clk cell_5484 ( .C ( clk ), .D ( signal_20176 ), .Q ( signal_20177 ) ) ;
    buf_clk cell_5488 ( .C ( clk ), .D ( signal_20180 ), .Q ( signal_20181 ) ) ;
    buf_clk cell_5492 ( .C ( clk ), .D ( signal_20184 ), .Q ( signal_20185 ) ) ;
    buf_clk cell_5496 ( .C ( clk ), .D ( signal_20188 ), .Q ( signal_20189 ) ) ;
    buf_clk cell_5500 ( .C ( clk ), .D ( signal_20192 ), .Q ( signal_20193 ) ) ;
    buf_clk cell_5504 ( .C ( clk ), .D ( signal_20196 ), .Q ( signal_20197 ) ) ;
    buf_clk cell_5506 ( .C ( clk ), .D ( signal_20198 ), .Q ( signal_20199 ) ) ;
    buf_clk cell_5508 ( .C ( clk ), .D ( signal_20200 ), .Q ( signal_20201 ) ) ;
    buf_clk cell_5510 ( .C ( clk ), .D ( signal_20202 ), .Q ( signal_20203 ) ) ;
    buf_clk cell_5512 ( .C ( clk ), .D ( signal_20204 ), .Q ( signal_20205 ) ) ;
    buf_clk cell_5514 ( .C ( clk ), .D ( signal_20206 ), .Q ( signal_20207 ) ) ;
    buf_clk cell_5520 ( .C ( clk ), .D ( signal_20212 ), .Q ( signal_20213 ) ) ;
    buf_clk cell_5526 ( .C ( clk ), .D ( signal_20218 ), .Q ( signal_20219 ) ) ;
    buf_clk cell_5532 ( .C ( clk ), .D ( signal_20224 ), .Q ( signal_20225 ) ) ;
    buf_clk cell_5538 ( .C ( clk ), .D ( signal_20230 ), .Q ( signal_20231 ) ) ;
    buf_clk cell_5544 ( .C ( clk ), .D ( signal_20236 ), .Q ( signal_20237 ) ) ;
    buf_clk cell_5548 ( .C ( clk ), .D ( signal_20240 ), .Q ( signal_20241 ) ) ;
    buf_clk cell_5552 ( .C ( clk ), .D ( signal_20244 ), .Q ( signal_20245 ) ) ;
    buf_clk cell_5556 ( .C ( clk ), .D ( signal_20248 ), .Q ( signal_20249 ) ) ;
    buf_clk cell_5560 ( .C ( clk ), .D ( signal_20252 ), .Q ( signal_20253 ) ) ;
    buf_clk cell_5564 ( .C ( clk ), .D ( signal_20256 ), .Q ( signal_20257 ) ) ;
    buf_clk cell_5570 ( .C ( clk ), .D ( signal_20262 ), .Q ( signal_20263 ) ) ;
    buf_clk cell_5576 ( .C ( clk ), .D ( signal_20268 ), .Q ( signal_20269 ) ) ;
    buf_clk cell_5582 ( .C ( clk ), .D ( signal_20274 ), .Q ( signal_20275 ) ) ;
    buf_clk cell_5588 ( .C ( clk ), .D ( signal_20280 ), .Q ( signal_20281 ) ) ;
    buf_clk cell_5594 ( .C ( clk ), .D ( signal_20286 ), .Q ( signal_20287 ) ) ;
    buf_clk cell_5598 ( .C ( clk ), .D ( signal_20290 ), .Q ( signal_20291 ) ) ;
    buf_clk cell_5602 ( .C ( clk ), .D ( signal_20294 ), .Q ( signal_20295 ) ) ;
    buf_clk cell_5606 ( .C ( clk ), .D ( signal_20298 ), .Q ( signal_20299 ) ) ;
    buf_clk cell_5610 ( .C ( clk ), .D ( signal_20302 ), .Q ( signal_20303 ) ) ;
    buf_clk cell_5614 ( .C ( clk ), .D ( signal_20306 ), .Q ( signal_20307 ) ) ;
    buf_clk cell_5618 ( .C ( clk ), .D ( signal_20310 ), .Q ( signal_20311 ) ) ;
    buf_clk cell_5622 ( .C ( clk ), .D ( signal_20314 ), .Q ( signal_20315 ) ) ;
    buf_clk cell_5626 ( .C ( clk ), .D ( signal_20318 ), .Q ( signal_20319 ) ) ;
    buf_clk cell_5630 ( .C ( clk ), .D ( signal_20322 ), .Q ( signal_20323 ) ) ;
    buf_clk cell_5634 ( .C ( clk ), .D ( signal_20326 ), .Q ( signal_20327 ) ) ;
    buf_clk cell_5638 ( .C ( clk ), .D ( signal_20330 ), .Q ( signal_20331 ) ) ;
    buf_clk cell_5642 ( .C ( clk ), .D ( signal_20334 ), .Q ( signal_20335 ) ) ;
    buf_clk cell_5646 ( .C ( clk ), .D ( signal_20338 ), .Q ( signal_20339 ) ) ;
    buf_clk cell_5650 ( .C ( clk ), .D ( signal_20342 ), .Q ( signal_20343 ) ) ;
    buf_clk cell_5654 ( .C ( clk ), .D ( signal_20346 ), .Q ( signal_20347 ) ) ;
    buf_clk cell_5656 ( .C ( clk ), .D ( signal_20348 ), .Q ( signal_20349 ) ) ;
    buf_clk cell_5658 ( .C ( clk ), .D ( signal_20350 ), .Q ( signal_20351 ) ) ;
    buf_clk cell_5660 ( .C ( clk ), .D ( signal_20352 ), .Q ( signal_20353 ) ) ;
    buf_clk cell_5662 ( .C ( clk ), .D ( signal_20354 ), .Q ( signal_20355 ) ) ;
    buf_clk cell_5664 ( .C ( clk ), .D ( signal_20356 ), .Q ( signal_20357 ) ) ;
    buf_clk cell_5668 ( .C ( clk ), .D ( signal_20360 ), .Q ( signal_20361 ) ) ;
    buf_clk cell_5672 ( .C ( clk ), .D ( signal_20364 ), .Q ( signal_20365 ) ) ;
    buf_clk cell_5676 ( .C ( clk ), .D ( signal_20368 ), .Q ( signal_20369 ) ) ;
    buf_clk cell_5680 ( .C ( clk ), .D ( signal_20372 ), .Q ( signal_20373 ) ) ;
    buf_clk cell_5684 ( .C ( clk ), .D ( signal_20376 ), .Q ( signal_20377 ) ) ;
    buf_clk cell_5688 ( .C ( clk ), .D ( signal_20380 ), .Q ( signal_20381 ) ) ;
    buf_clk cell_5692 ( .C ( clk ), .D ( signal_20384 ), .Q ( signal_20385 ) ) ;
    buf_clk cell_5696 ( .C ( clk ), .D ( signal_20388 ), .Q ( signal_20389 ) ) ;
    buf_clk cell_5700 ( .C ( clk ), .D ( signal_20392 ), .Q ( signal_20393 ) ) ;
    buf_clk cell_5704 ( .C ( clk ), .D ( signal_20396 ), .Q ( signal_20397 ) ) ;
    buf_clk cell_5710 ( .C ( clk ), .D ( signal_20402 ), .Q ( signal_20403 ) ) ;
    buf_clk cell_5716 ( .C ( clk ), .D ( signal_20408 ), .Q ( signal_20409 ) ) ;
    buf_clk cell_5722 ( .C ( clk ), .D ( signal_20414 ), .Q ( signal_20415 ) ) ;
    buf_clk cell_5728 ( .C ( clk ), .D ( signal_20420 ), .Q ( signal_20421 ) ) ;
    buf_clk cell_5734 ( .C ( clk ), .D ( signal_20426 ), .Q ( signal_20427 ) ) ;
    buf_clk cell_5736 ( .C ( clk ), .D ( signal_20428 ), .Q ( signal_20429 ) ) ;
    buf_clk cell_5738 ( .C ( clk ), .D ( signal_20430 ), .Q ( signal_20431 ) ) ;
    buf_clk cell_5740 ( .C ( clk ), .D ( signal_20432 ), .Q ( signal_20433 ) ) ;
    buf_clk cell_5742 ( .C ( clk ), .D ( signal_20434 ), .Q ( signal_20435 ) ) ;
    buf_clk cell_5744 ( .C ( clk ), .D ( signal_20436 ), .Q ( signal_20437 ) ) ;
    buf_clk cell_5746 ( .C ( clk ), .D ( signal_20438 ), .Q ( signal_20439 ) ) ;
    buf_clk cell_5748 ( .C ( clk ), .D ( signal_20440 ), .Q ( signal_20441 ) ) ;
    buf_clk cell_5750 ( .C ( clk ), .D ( signal_20442 ), .Q ( signal_20443 ) ) ;
    buf_clk cell_5752 ( .C ( clk ), .D ( signal_20444 ), .Q ( signal_20445 ) ) ;
    buf_clk cell_5754 ( .C ( clk ), .D ( signal_20446 ), .Q ( signal_20447 ) ) ;
    buf_clk cell_5758 ( .C ( clk ), .D ( signal_20450 ), .Q ( signal_20451 ) ) ;
    buf_clk cell_5762 ( .C ( clk ), .D ( signal_20454 ), .Q ( signal_20455 ) ) ;
    buf_clk cell_5766 ( .C ( clk ), .D ( signal_20458 ), .Q ( signal_20459 ) ) ;
    buf_clk cell_5770 ( .C ( clk ), .D ( signal_20462 ), .Q ( signal_20463 ) ) ;
    buf_clk cell_5774 ( .C ( clk ), .D ( signal_20466 ), .Q ( signal_20467 ) ) ;
    buf_clk cell_5780 ( .C ( clk ), .D ( signal_20472 ), .Q ( signal_20473 ) ) ;
    buf_clk cell_5786 ( .C ( clk ), .D ( signal_20478 ), .Q ( signal_20479 ) ) ;
    buf_clk cell_5792 ( .C ( clk ), .D ( signal_20484 ), .Q ( signal_20485 ) ) ;
    buf_clk cell_5798 ( .C ( clk ), .D ( signal_20490 ), .Q ( signal_20491 ) ) ;
    buf_clk cell_5804 ( .C ( clk ), .D ( signal_20496 ), .Q ( signal_20497 ) ) ;
    buf_clk cell_5810 ( .C ( clk ), .D ( signal_20502 ), .Q ( signal_20503 ) ) ;
    buf_clk cell_5816 ( .C ( clk ), .D ( signal_20508 ), .Q ( signal_20509 ) ) ;
    buf_clk cell_5822 ( .C ( clk ), .D ( signal_20514 ), .Q ( signal_20515 ) ) ;
    buf_clk cell_5828 ( .C ( clk ), .D ( signal_20520 ), .Q ( signal_20521 ) ) ;
    buf_clk cell_5834 ( .C ( clk ), .D ( signal_20526 ), .Q ( signal_20527 ) ) ;
    buf_clk cell_5840 ( .C ( clk ), .D ( signal_20532 ), .Q ( signal_20533 ) ) ;
    buf_clk cell_5846 ( .C ( clk ), .D ( signal_20538 ), .Q ( signal_20539 ) ) ;
    buf_clk cell_5852 ( .C ( clk ), .D ( signal_20544 ), .Q ( signal_20545 ) ) ;
    buf_clk cell_5858 ( .C ( clk ), .D ( signal_20550 ), .Q ( signal_20551 ) ) ;
    buf_clk cell_5864 ( .C ( clk ), .D ( signal_20556 ), .Q ( signal_20557 ) ) ;
    buf_clk cell_5868 ( .C ( clk ), .D ( signal_20560 ), .Q ( signal_20561 ) ) ;
    buf_clk cell_5872 ( .C ( clk ), .D ( signal_20564 ), .Q ( signal_20565 ) ) ;
    buf_clk cell_5876 ( .C ( clk ), .D ( signal_20568 ), .Q ( signal_20569 ) ) ;
    buf_clk cell_5880 ( .C ( clk ), .D ( signal_20572 ), .Q ( signal_20573 ) ) ;
    buf_clk cell_5884 ( .C ( clk ), .D ( signal_20576 ), .Q ( signal_20577 ) ) ;
    buf_clk cell_5886 ( .C ( clk ), .D ( signal_20578 ), .Q ( signal_20579 ) ) ;
    buf_clk cell_5888 ( .C ( clk ), .D ( signal_20580 ), .Q ( signal_20581 ) ) ;
    buf_clk cell_5890 ( .C ( clk ), .D ( signal_20582 ), .Q ( signal_20583 ) ) ;
    buf_clk cell_5892 ( .C ( clk ), .D ( signal_20584 ), .Q ( signal_20585 ) ) ;
    buf_clk cell_5894 ( .C ( clk ), .D ( signal_20586 ), .Q ( signal_20587 ) ) ;
    buf_clk cell_5896 ( .C ( clk ), .D ( signal_20588 ), .Q ( signal_20589 ) ) ;
    buf_clk cell_5898 ( .C ( clk ), .D ( signal_20590 ), .Q ( signal_20591 ) ) ;
    buf_clk cell_5900 ( .C ( clk ), .D ( signal_20592 ), .Q ( signal_20593 ) ) ;
    buf_clk cell_5902 ( .C ( clk ), .D ( signal_20594 ), .Q ( signal_20595 ) ) ;
    buf_clk cell_5904 ( .C ( clk ), .D ( signal_20596 ), .Q ( signal_20597 ) ) ;
    buf_clk cell_5910 ( .C ( clk ), .D ( signal_20602 ), .Q ( signal_20603 ) ) ;
    buf_clk cell_5918 ( .C ( clk ), .D ( signal_20610 ), .Q ( signal_20611 ) ) ;
    buf_clk cell_5926 ( .C ( clk ), .D ( signal_20618 ), .Q ( signal_20619 ) ) ;
    buf_clk cell_5934 ( .C ( clk ), .D ( signal_20626 ), .Q ( signal_20627 ) ) ;
    buf_clk cell_5942 ( .C ( clk ), .D ( signal_20634 ), .Q ( signal_20635 ) ) ;
    buf_clk cell_5946 ( .C ( clk ), .D ( signal_20638 ), .Q ( signal_20639 ) ) ;
    buf_clk cell_5950 ( .C ( clk ), .D ( signal_20642 ), .Q ( signal_20643 ) ) ;
    buf_clk cell_5954 ( .C ( clk ), .D ( signal_20646 ), .Q ( signal_20647 ) ) ;
    buf_clk cell_5958 ( .C ( clk ), .D ( signal_20650 ), .Q ( signal_20651 ) ) ;
    buf_clk cell_5962 ( .C ( clk ), .D ( signal_20654 ), .Q ( signal_20655 ) ) ;
    buf_clk cell_5968 ( .C ( clk ), .D ( signal_20660 ), .Q ( signal_20661 ) ) ;
    buf_clk cell_5974 ( .C ( clk ), .D ( signal_20666 ), .Q ( signal_20667 ) ) ;
    buf_clk cell_5980 ( .C ( clk ), .D ( signal_20672 ), .Q ( signal_20673 ) ) ;
    buf_clk cell_5986 ( .C ( clk ), .D ( signal_20678 ), .Q ( signal_20679 ) ) ;
    buf_clk cell_5992 ( .C ( clk ), .D ( signal_20684 ), .Q ( signal_20685 ) ) ;
    buf_clk cell_5998 ( .C ( clk ), .D ( signal_20690 ), .Q ( signal_20691 ) ) ;
    buf_clk cell_6004 ( .C ( clk ), .D ( signal_20696 ), .Q ( signal_20697 ) ) ;
    buf_clk cell_6010 ( .C ( clk ), .D ( signal_20702 ), .Q ( signal_20703 ) ) ;
    buf_clk cell_6016 ( .C ( clk ), .D ( signal_20708 ), .Q ( signal_20709 ) ) ;
    buf_clk cell_6022 ( .C ( clk ), .D ( signal_20714 ), .Q ( signal_20715 ) ) ;
    buf_clk cell_6026 ( .C ( clk ), .D ( signal_20718 ), .Q ( signal_20719 ) ) ;
    buf_clk cell_6030 ( .C ( clk ), .D ( signal_20722 ), .Q ( signal_20723 ) ) ;
    buf_clk cell_6034 ( .C ( clk ), .D ( signal_20726 ), .Q ( signal_20727 ) ) ;
    buf_clk cell_6038 ( .C ( clk ), .D ( signal_20730 ), .Q ( signal_20731 ) ) ;
    buf_clk cell_6042 ( .C ( clk ), .D ( signal_20734 ), .Q ( signal_20735 ) ) ;
    buf_clk cell_6048 ( .C ( clk ), .D ( signal_20740 ), .Q ( signal_20741 ) ) ;
    buf_clk cell_6054 ( .C ( clk ), .D ( signal_20746 ), .Q ( signal_20747 ) ) ;
    buf_clk cell_6060 ( .C ( clk ), .D ( signal_20752 ), .Q ( signal_20753 ) ) ;
    buf_clk cell_6066 ( .C ( clk ), .D ( signal_20758 ), .Q ( signal_20759 ) ) ;
    buf_clk cell_6072 ( .C ( clk ), .D ( signal_20764 ), .Q ( signal_20765 ) ) ;
    buf_clk cell_6076 ( .C ( clk ), .D ( signal_20768 ), .Q ( signal_20769 ) ) ;
    buf_clk cell_6080 ( .C ( clk ), .D ( signal_20772 ), .Q ( signal_20773 ) ) ;
    buf_clk cell_6084 ( .C ( clk ), .D ( signal_20776 ), .Q ( signal_20777 ) ) ;
    buf_clk cell_6088 ( .C ( clk ), .D ( signal_20780 ), .Q ( signal_20781 ) ) ;
    buf_clk cell_6092 ( .C ( clk ), .D ( signal_20784 ), .Q ( signal_20785 ) ) ;
    buf_clk cell_6096 ( .C ( clk ), .D ( signal_20788 ), .Q ( signal_20789 ) ) ;
    buf_clk cell_6100 ( .C ( clk ), .D ( signal_20792 ), .Q ( signal_20793 ) ) ;
    buf_clk cell_6104 ( .C ( clk ), .D ( signal_20796 ), .Q ( signal_20797 ) ) ;
    buf_clk cell_6108 ( .C ( clk ), .D ( signal_20800 ), .Q ( signal_20801 ) ) ;
    buf_clk cell_6112 ( .C ( clk ), .D ( signal_20804 ), .Q ( signal_20805 ) ) ;
    buf_clk cell_6138 ( .C ( clk ), .D ( signal_20830 ), .Q ( signal_20831 ) ) ;
    buf_clk cell_6144 ( .C ( clk ), .D ( signal_20836 ), .Q ( signal_20837 ) ) ;
    buf_clk cell_6150 ( .C ( clk ), .D ( signal_20842 ), .Q ( signal_20843 ) ) ;
    buf_clk cell_6156 ( .C ( clk ), .D ( signal_20848 ), .Q ( signal_20849 ) ) ;
    buf_clk cell_6162 ( .C ( clk ), .D ( signal_20854 ), .Q ( signal_20855 ) ) ;
    buf_clk cell_6168 ( .C ( clk ), .D ( signal_20860 ), .Q ( signal_20861 ) ) ;
    buf_clk cell_6174 ( .C ( clk ), .D ( signal_20866 ), .Q ( signal_20867 ) ) ;
    buf_clk cell_6180 ( .C ( clk ), .D ( signal_20872 ), .Q ( signal_20873 ) ) ;
    buf_clk cell_6186 ( .C ( clk ), .D ( signal_20878 ), .Q ( signal_20879 ) ) ;
    buf_clk cell_6192 ( .C ( clk ), .D ( signal_20884 ), .Q ( signal_20885 ) ) ;
    buf_clk cell_6198 ( .C ( clk ), .D ( signal_20890 ), .Q ( signal_20891 ) ) ;
    buf_clk cell_6204 ( .C ( clk ), .D ( signal_20896 ), .Q ( signal_20897 ) ) ;
    buf_clk cell_6210 ( .C ( clk ), .D ( signal_20902 ), .Q ( signal_20903 ) ) ;
    buf_clk cell_6216 ( .C ( clk ), .D ( signal_20908 ), .Q ( signal_20909 ) ) ;
    buf_clk cell_6222 ( .C ( clk ), .D ( signal_20914 ), .Q ( signal_20915 ) ) ;
    buf_clk cell_6236 ( .C ( clk ), .D ( signal_20928 ), .Q ( signal_20929 ) ) ;
    buf_clk cell_6240 ( .C ( clk ), .D ( signal_20932 ), .Q ( signal_20933 ) ) ;
    buf_clk cell_6244 ( .C ( clk ), .D ( signal_20936 ), .Q ( signal_20937 ) ) ;
    buf_clk cell_6248 ( .C ( clk ), .D ( signal_20940 ), .Q ( signal_20941 ) ) ;
    buf_clk cell_6252 ( .C ( clk ), .D ( signal_20944 ), .Q ( signal_20945 ) ) ;
    buf_clk cell_6258 ( .C ( clk ), .D ( signal_20950 ), .Q ( signal_20951 ) ) ;
    buf_clk cell_6264 ( .C ( clk ), .D ( signal_20956 ), .Q ( signal_20957 ) ) ;
    buf_clk cell_6270 ( .C ( clk ), .D ( signal_20962 ), .Q ( signal_20963 ) ) ;
    buf_clk cell_6276 ( .C ( clk ), .D ( signal_20968 ), .Q ( signal_20969 ) ) ;
    buf_clk cell_6282 ( .C ( clk ), .D ( signal_20974 ), .Q ( signal_20975 ) ) ;
    buf_clk cell_6298 ( .C ( clk ), .D ( signal_20990 ), .Q ( signal_20991 ) ) ;
    buf_clk cell_6304 ( .C ( clk ), .D ( signal_20996 ), .Q ( signal_20997 ) ) ;
    buf_clk cell_6310 ( .C ( clk ), .D ( signal_21002 ), .Q ( signal_21003 ) ) ;
    buf_clk cell_6316 ( .C ( clk ), .D ( signal_21008 ), .Q ( signal_21009 ) ) ;
    buf_clk cell_6322 ( .C ( clk ), .D ( signal_21014 ), .Q ( signal_21015 ) ) ;
    buf_clk cell_6340 ( .C ( clk ), .D ( signal_21032 ), .Q ( signal_21033 ) ) ;
    buf_clk cell_6348 ( .C ( clk ), .D ( signal_21040 ), .Q ( signal_21041 ) ) ;
    buf_clk cell_6356 ( .C ( clk ), .D ( signal_21048 ), .Q ( signal_21049 ) ) ;
    buf_clk cell_6364 ( .C ( clk ), .D ( signal_21056 ), .Q ( signal_21057 ) ) ;
    buf_clk cell_6372 ( .C ( clk ), .D ( signal_21064 ), .Q ( signal_21065 ) ) ;
    buf_clk cell_6376 ( .C ( clk ), .D ( signal_21068 ), .Q ( signal_21069 ) ) ;
    buf_clk cell_6380 ( .C ( clk ), .D ( signal_21072 ), .Q ( signal_21073 ) ) ;
    buf_clk cell_6384 ( .C ( clk ), .D ( signal_21076 ), .Q ( signal_21077 ) ) ;
    buf_clk cell_6388 ( .C ( clk ), .D ( signal_21080 ), .Q ( signal_21081 ) ) ;
    buf_clk cell_6392 ( .C ( clk ), .D ( signal_21084 ), .Q ( signal_21085 ) ) ;
    buf_clk cell_6396 ( .C ( clk ), .D ( signal_21088 ), .Q ( signal_21089 ) ) ;
    buf_clk cell_6400 ( .C ( clk ), .D ( signal_21092 ), .Q ( signal_21093 ) ) ;
    buf_clk cell_6404 ( .C ( clk ), .D ( signal_21096 ), .Q ( signal_21097 ) ) ;
    buf_clk cell_6408 ( .C ( clk ), .D ( signal_21100 ), .Q ( signal_21101 ) ) ;
    buf_clk cell_6412 ( .C ( clk ), .D ( signal_21104 ), .Q ( signal_21105 ) ) ;
    buf_clk cell_6418 ( .C ( clk ), .D ( signal_21110 ), .Q ( signal_21111 ) ) ;
    buf_clk cell_6424 ( .C ( clk ), .D ( signal_21116 ), .Q ( signal_21117 ) ) ;
    buf_clk cell_6430 ( .C ( clk ), .D ( signal_21122 ), .Q ( signal_21123 ) ) ;
    buf_clk cell_6436 ( .C ( clk ), .D ( signal_21128 ), .Q ( signal_21129 ) ) ;
    buf_clk cell_6442 ( .C ( clk ), .D ( signal_21134 ), .Q ( signal_21135 ) ) ;
    buf_clk cell_6448 ( .C ( clk ), .D ( signal_21140 ), .Q ( signal_21141 ) ) ;
    buf_clk cell_6454 ( .C ( clk ), .D ( signal_21146 ), .Q ( signal_21147 ) ) ;
    buf_clk cell_6460 ( .C ( clk ), .D ( signal_21152 ), .Q ( signal_21153 ) ) ;
    buf_clk cell_6466 ( .C ( clk ), .D ( signal_21158 ), .Q ( signal_21159 ) ) ;
    buf_clk cell_6472 ( .C ( clk ), .D ( signal_21164 ), .Q ( signal_21165 ) ) ;
    buf_clk cell_6476 ( .C ( clk ), .D ( signal_21168 ), .Q ( signal_21169 ) ) ;
    buf_clk cell_6480 ( .C ( clk ), .D ( signal_21172 ), .Q ( signal_21173 ) ) ;
    buf_clk cell_6484 ( .C ( clk ), .D ( signal_21176 ), .Q ( signal_21177 ) ) ;
    buf_clk cell_6488 ( .C ( clk ), .D ( signal_21180 ), .Q ( signal_21181 ) ) ;
    buf_clk cell_6492 ( .C ( clk ), .D ( signal_21184 ), .Q ( signal_21185 ) ) ;
    buf_clk cell_6500 ( .C ( clk ), .D ( signal_21192 ), .Q ( signal_21193 ) ) ;
    buf_clk cell_6508 ( .C ( clk ), .D ( signal_21200 ), .Q ( signal_21201 ) ) ;
    buf_clk cell_6516 ( .C ( clk ), .D ( signal_21208 ), .Q ( signal_21209 ) ) ;
    buf_clk cell_6524 ( .C ( clk ), .D ( signal_21216 ), .Q ( signal_21217 ) ) ;
    buf_clk cell_6532 ( .C ( clk ), .D ( signal_21224 ), .Q ( signal_21225 ) ) ;
    buf_clk cell_6538 ( .C ( clk ), .D ( signal_21230 ), .Q ( signal_21231 ) ) ;
    buf_clk cell_6544 ( .C ( clk ), .D ( signal_21236 ), .Q ( signal_21237 ) ) ;
    buf_clk cell_6550 ( .C ( clk ), .D ( signal_21242 ), .Q ( signal_21243 ) ) ;
    buf_clk cell_6556 ( .C ( clk ), .D ( signal_21248 ), .Q ( signal_21249 ) ) ;
    buf_clk cell_6562 ( .C ( clk ), .D ( signal_21254 ), .Q ( signal_21255 ) ) ;
    buf_clk cell_6568 ( .C ( clk ), .D ( signal_21260 ), .Q ( signal_21261 ) ) ;
    buf_clk cell_6574 ( .C ( clk ), .D ( signal_21266 ), .Q ( signal_21267 ) ) ;
    buf_clk cell_6580 ( .C ( clk ), .D ( signal_21272 ), .Q ( signal_21273 ) ) ;
    buf_clk cell_6586 ( .C ( clk ), .D ( signal_21278 ), .Q ( signal_21279 ) ) ;
    buf_clk cell_6592 ( .C ( clk ), .D ( signal_21284 ), .Q ( signal_21285 ) ) ;
    buf_clk cell_6618 ( .C ( clk ), .D ( signal_21310 ), .Q ( signal_21311 ) ) ;
    buf_clk cell_6624 ( .C ( clk ), .D ( signal_21316 ), .Q ( signal_21317 ) ) ;
    buf_clk cell_6630 ( .C ( clk ), .D ( signal_21322 ), .Q ( signal_21323 ) ) ;
    buf_clk cell_6636 ( .C ( clk ), .D ( signal_21328 ), .Q ( signal_21329 ) ) ;
    buf_clk cell_6642 ( .C ( clk ), .D ( signal_21334 ), .Q ( signal_21335 ) ) ;
    buf_clk cell_6668 ( .C ( clk ), .D ( signal_21360 ), .Q ( signal_21361 ) ) ;
    buf_clk cell_6674 ( .C ( clk ), .D ( signal_21366 ), .Q ( signal_21367 ) ) ;
    buf_clk cell_6680 ( .C ( clk ), .D ( signal_21372 ), .Q ( signal_21373 ) ) ;
    buf_clk cell_6686 ( .C ( clk ), .D ( signal_21378 ), .Q ( signal_21379 ) ) ;
    buf_clk cell_6692 ( .C ( clk ), .D ( signal_21384 ), .Q ( signal_21385 ) ) ;
    buf_clk cell_6698 ( .C ( clk ), .D ( signal_21390 ), .Q ( signal_21391 ) ) ;
    buf_clk cell_6704 ( .C ( clk ), .D ( signal_21396 ), .Q ( signal_21397 ) ) ;
    buf_clk cell_6710 ( .C ( clk ), .D ( signal_21402 ), .Q ( signal_21403 ) ) ;
    buf_clk cell_6716 ( .C ( clk ), .D ( signal_21408 ), .Q ( signal_21409 ) ) ;
    buf_clk cell_6722 ( .C ( clk ), .D ( signal_21414 ), .Q ( signal_21415 ) ) ;
    buf_clk cell_6726 ( .C ( clk ), .D ( signal_21418 ), .Q ( signal_21419 ) ) ;
    buf_clk cell_6730 ( .C ( clk ), .D ( signal_21422 ), .Q ( signal_21423 ) ) ;
    buf_clk cell_6734 ( .C ( clk ), .D ( signal_21426 ), .Q ( signal_21427 ) ) ;
    buf_clk cell_6738 ( .C ( clk ), .D ( signal_21430 ), .Q ( signal_21431 ) ) ;
    buf_clk cell_6742 ( .C ( clk ), .D ( signal_21434 ), .Q ( signal_21435 ) ) ;
    buf_clk cell_6750 ( .C ( clk ), .D ( signal_21442 ), .Q ( signal_21443 ) ) ;
    buf_clk cell_6760 ( .C ( clk ), .D ( signal_21452 ), .Q ( signal_21453 ) ) ;
    buf_clk cell_6770 ( .C ( clk ), .D ( signal_21462 ), .Q ( signal_21463 ) ) ;
    buf_clk cell_6780 ( .C ( clk ), .D ( signal_21472 ), .Q ( signal_21473 ) ) ;
    buf_clk cell_6790 ( .C ( clk ), .D ( signal_21482 ), .Q ( signal_21483 ) ) ;
    buf_clk cell_6796 ( .C ( clk ), .D ( signal_21488 ), .Q ( signal_21489 ) ) ;
    buf_clk cell_6802 ( .C ( clk ), .D ( signal_21494 ), .Q ( signal_21495 ) ) ;
    buf_clk cell_6808 ( .C ( clk ), .D ( signal_21500 ), .Q ( signal_21501 ) ) ;
    buf_clk cell_6814 ( .C ( clk ), .D ( signal_21506 ), .Q ( signal_21507 ) ) ;
    buf_clk cell_6820 ( .C ( clk ), .D ( signal_21512 ), .Q ( signal_21513 ) ) ;
    buf_clk cell_6828 ( .C ( clk ), .D ( signal_21520 ), .Q ( signal_21521 ) ) ;
    buf_clk cell_6836 ( .C ( clk ), .D ( signal_21528 ), .Q ( signal_21529 ) ) ;
    buf_clk cell_6844 ( .C ( clk ), .D ( signal_21536 ), .Q ( signal_21537 ) ) ;
    buf_clk cell_6852 ( .C ( clk ), .D ( signal_21544 ), .Q ( signal_21545 ) ) ;
    buf_clk cell_6860 ( .C ( clk ), .D ( signal_21552 ), .Q ( signal_21553 ) ) ;
    buf_clk cell_6868 ( .C ( clk ), .D ( signal_21560 ), .Q ( signal_21561 ) ) ;
    buf_clk cell_6876 ( .C ( clk ), .D ( signal_21568 ), .Q ( signal_21569 ) ) ;
    buf_clk cell_6884 ( .C ( clk ), .D ( signal_21576 ), .Q ( signal_21577 ) ) ;
    buf_clk cell_6892 ( .C ( clk ), .D ( signal_21584 ), .Q ( signal_21585 ) ) ;
    buf_clk cell_6900 ( .C ( clk ), .D ( signal_21592 ), .Q ( signal_21593 ) ) ;
    buf_clk cell_6990 ( .C ( clk ), .D ( signal_21682 ), .Q ( signal_21683 ) ) ;
    buf_clk cell_7000 ( .C ( clk ), .D ( signal_21692 ), .Q ( signal_21693 ) ) ;
    buf_clk cell_7010 ( .C ( clk ), .D ( signal_21702 ), .Q ( signal_21703 ) ) ;
    buf_clk cell_7020 ( .C ( clk ), .D ( signal_21712 ), .Q ( signal_21713 ) ) ;
    buf_clk cell_7030 ( .C ( clk ), .D ( signal_21722 ), .Q ( signal_21723 ) ) ;
    buf_clk cell_7036 ( .C ( clk ), .D ( signal_21728 ), .Q ( signal_21729 ) ) ;
    buf_clk cell_7042 ( .C ( clk ), .D ( signal_21734 ), .Q ( signal_21735 ) ) ;
    buf_clk cell_7048 ( .C ( clk ), .D ( signal_21740 ), .Q ( signal_21741 ) ) ;
    buf_clk cell_7054 ( .C ( clk ), .D ( signal_21746 ), .Q ( signal_21747 ) ) ;
    buf_clk cell_7060 ( .C ( clk ), .D ( signal_21752 ), .Q ( signal_21753 ) ) ;
    buf_clk cell_7078 ( .C ( clk ), .D ( signal_21770 ), .Q ( signal_21771 ) ) ;
    buf_clk cell_7086 ( .C ( clk ), .D ( signal_21778 ), .Q ( signal_21779 ) ) ;
    buf_clk cell_7094 ( .C ( clk ), .D ( signal_21786 ), .Q ( signal_21787 ) ) ;
    buf_clk cell_7102 ( .C ( clk ), .D ( signal_21794 ), .Q ( signal_21795 ) ) ;
    buf_clk cell_7110 ( .C ( clk ), .D ( signal_21802 ), .Q ( signal_21803 ) ) ;
    buf_clk cell_7116 ( .C ( clk ), .D ( signal_21808 ), .Q ( signal_21809 ) ) ;
    buf_clk cell_7122 ( .C ( clk ), .D ( signal_21814 ), .Q ( signal_21815 ) ) ;
    buf_clk cell_7128 ( .C ( clk ), .D ( signal_21820 ), .Q ( signal_21821 ) ) ;
    buf_clk cell_7134 ( .C ( clk ), .D ( signal_21826 ), .Q ( signal_21827 ) ) ;
    buf_clk cell_7140 ( .C ( clk ), .D ( signal_21832 ), .Q ( signal_21833 ) ) ;
    buf_clk cell_7148 ( .C ( clk ), .D ( signal_21840 ), .Q ( signal_21841 ) ) ;
    buf_clk cell_7156 ( .C ( clk ), .D ( signal_21848 ), .Q ( signal_21849 ) ) ;
    buf_clk cell_7164 ( .C ( clk ), .D ( signal_21856 ), .Q ( signal_21857 ) ) ;
    buf_clk cell_7172 ( .C ( clk ), .D ( signal_21864 ), .Q ( signal_21865 ) ) ;
    buf_clk cell_7180 ( .C ( clk ), .D ( signal_21872 ), .Q ( signal_21873 ) ) ;
    buf_clk cell_7188 ( .C ( clk ), .D ( signal_21880 ), .Q ( signal_21881 ) ) ;
    buf_clk cell_7196 ( .C ( clk ), .D ( signal_21888 ), .Q ( signal_21889 ) ) ;
    buf_clk cell_7204 ( .C ( clk ), .D ( signal_21896 ), .Q ( signal_21897 ) ) ;
    buf_clk cell_7212 ( .C ( clk ), .D ( signal_21904 ), .Q ( signal_21905 ) ) ;
    buf_clk cell_7220 ( .C ( clk ), .D ( signal_21912 ), .Q ( signal_21913 ) ) ;
    buf_clk cell_7228 ( .C ( clk ), .D ( signal_21920 ), .Q ( signal_21921 ) ) ;
    buf_clk cell_7236 ( .C ( clk ), .D ( signal_21928 ), .Q ( signal_21929 ) ) ;
    buf_clk cell_7244 ( .C ( clk ), .D ( signal_21936 ), .Q ( signal_21937 ) ) ;
    buf_clk cell_7252 ( .C ( clk ), .D ( signal_21944 ), .Q ( signal_21945 ) ) ;
    buf_clk cell_7260 ( .C ( clk ), .D ( signal_21952 ), .Q ( signal_21953 ) ) ;
    buf_clk cell_7270 ( .C ( clk ), .D ( signal_21962 ), .Q ( signal_21963 ) ) ;
    buf_clk cell_7280 ( .C ( clk ), .D ( signal_21972 ), .Q ( signal_21973 ) ) ;
    buf_clk cell_7290 ( .C ( clk ), .D ( signal_21982 ), .Q ( signal_21983 ) ) ;
    buf_clk cell_7300 ( .C ( clk ), .D ( signal_21992 ), .Q ( signal_21993 ) ) ;
    buf_clk cell_7310 ( .C ( clk ), .D ( signal_22002 ), .Q ( signal_22003 ) ) ;
    buf_clk cell_7318 ( .C ( clk ), .D ( signal_22010 ), .Q ( signal_22011 ) ) ;
    buf_clk cell_7326 ( .C ( clk ), .D ( signal_22018 ), .Q ( signal_22019 ) ) ;
    buf_clk cell_7334 ( .C ( clk ), .D ( signal_22026 ), .Q ( signal_22027 ) ) ;
    buf_clk cell_7342 ( .C ( clk ), .D ( signal_22034 ), .Q ( signal_22035 ) ) ;
    buf_clk cell_7350 ( .C ( clk ), .D ( signal_22042 ), .Q ( signal_22043 ) ) ;
    buf_clk cell_7358 ( .C ( clk ), .D ( signal_22050 ), .Q ( signal_22051 ) ) ;
    buf_clk cell_7366 ( .C ( clk ), .D ( signal_22058 ), .Q ( signal_22059 ) ) ;
    buf_clk cell_7374 ( .C ( clk ), .D ( signal_22066 ), .Q ( signal_22067 ) ) ;
    buf_clk cell_7382 ( .C ( clk ), .D ( signal_22074 ), .Q ( signal_22075 ) ) ;
    buf_clk cell_7390 ( .C ( clk ), .D ( signal_22082 ), .Q ( signal_22083 ) ) ;
    buf_clk cell_7408 ( .C ( clk ), .D ( signal_22100 ), .Q ( signal_22101 ) ) ;
    buf_clk cell_7416 ( .C ( clk ), .D ( signal_22108 ), .Q ( signal_22109 ) ) ;
    buf_clk cell_7424 ( .C ( clk ), .D ( signal_22116 ), .Q ( signal_22117 ) ) ;
    buf_clk cell_7432 ( .C ( clk ), .D ( signal_22124 ), .Q ( signal_22125 ) ) ;
    buf_clk cell_7440 ( .C ( clk ), .D ( signal_22132 ), .Q ( signal_22133 ) ) ;
    buf_clk cell_7448 ( .C ( clk ), .D ( signal_22140 ), .Q ( signal_22141 ) ) ;
    buf_clk cell_7456 ( .C ( clk ), .D ( signal_22148 ), .Q ( signal_22149 ) ) ;
    buf_clk cell_7464 ( .C ( clk ), .D ( signal_22156 ), .Q ( signal_22157 ) ) ;
    buf_clk cell_7472 ( .C ( clk ), .D ( signal_22164 ), .Q ( signal_22165 ) ) ;
    buf_clk cell_7480 ( .C ( clk ), .D ( signal_22172 ), .Q ( signal_22173 ) ) ;
    buf_clk cell_7488 ( .C ( clk ), .D ( signal_22180 ), .Q ( signal_22181 ) ) ;
    buf_clk cell_7496 ( .C ( clk ), .D ( signal_22188 ), .Q ( signal_22189 ) ) ;
    buf_clk cell_7504 ( .C ( clk ), .D ( signal_22196 ), .Q ( signal_22197 ) ) ;
    buf_clk cell_7512 ( .C ( clk ), .D ( signal_22204 ), .Q ( signal_22205 ) ) ;
    buf_clk cell_7520 ( .C ( clk ), .D ( signal_22212 ), .Q ( signal_22213 ) ) ;
    buf_clk cell_7556 ( .C ( clk ), .D ( signal_22248 ), .Q ( signal_22249 ) ) ;
    buf_clk cell_7564 ( .C ( clk ), .D ( signal_22256 ), .Q ( signal_22257 ) ) ;
    buf_clk cell_7572 ( .C ( clk ), .D ( signal_22264 ), .Q ( signal_22265 ) ) ;
    buf_clk cell_7580 ( .C ( clk ), .D ( signal_22272 ), .Q ( signal_22273 ) ) ;
    buf_clk cell_7588 ( .C ( clk ), .D ( signal_22280 ), .Q ( signal_22281 ) ) ;
    buf_clk cell_7656 ( .C ( clk ), .D ( signal_22348 ), .Q ( signal_22349 ) ) ;
    buf_clk cell_7664 ( .C ( clk ), .D ( signal_22356 ), .Q ( signal_22357 ) ) ;
    buf_clk cell_7672 ( .C ( clk ), .D ( signal_22364 ), .Q ( signal_22365 ) ) ;
    buf_clk cell_7680 ( .C ( clk ), .D ( signal_22372 ), .Q ( signal_22373 ) ) ;
    buf_clk cell_7688 ( .C ( clk ), .D ( signal_22380 ), .Q ( signal_22381 ) ) ;
    buf_clk cell_7698 ( .C ( clk ), .D ( signal_22390 ), .Q ( signal_22391 ) ) ;
    buf_clk cell_7708 ( .C ( clk ), .D ( signal_22400 ), .Q ( signal_22401 ) ) ;
    buf_clk cell_7718 ( .C ( clk ), .D ( signal_22410 ), .Q ( signal_22411 ) ) ;
    buf_clk cell_7728 ( .C ( clk ), .D ( signal_22420 ), .Q ( signal_22421 ) ) ;
    buf_clk cell_7738 ( .C ( clk ), .D ( signal_22430 ), .Q ( signal_22431 ) ) ;
    buf_clk cell_7786 ( .C ( clk ), .D ( signal_22478 ), .Q ( signal_22479 ) ) ;
    buf_clk cell_7794 ( .C ( clk ), .D ( signal_22486 ), .Q ( signal_22487 ) ) ;
    buf_clk cell_7802 ( .C ( clk ), .D ( signal_22494 ), .Q ( signal_22495 ) ) ;
    buf_clk cell_7810 ( .C ( clk ), .D ( signal_22502 ), .Q ( signal_22503 ) ) ;
    buf_clk cell_7818 ( .C ( clk ), .D ( signal_22510 ), .Q ( signal_22511 ) ) ;
    buf_clk cell_7828 ( .C ( clk ), .D ( signal_22520 ), .Q ( signal_22521 ) ) ;
    buf_clk cell_7838 ( .C ( clk ), .D ( signal_22530 ), .Q ( signal_22531 ) ) ;
    buf_clk cell_7848 ( .C ( clk ), .D ( signal_22540 ), .Q ( signal_22541 ) ) ;
    buf_clk cell_7858 ( .C ( clk ), .D ( signal_22550 ), .Q ( signal_22551 ) ) ;
    buf_clk cell_7868 ( .C ( clk ), .D ( signal_22560 ), .Q ( signal_22561 ) ) ;
    buf_clk cell_7876 ( .C ( clk ), .D ( signal_22568 ), .Q ( signal_22569 ) ) ;
    buf_clk cell_7884 ( .C ( clk ), .D ( signal_22576 ), .Q ( signal_22577 ) ) ;
    buf_clk cell_7892 ( .C ( clk ), .D ( signal_22584 ), .Q ( signal_22585 ) ) ;
    buf_clk cell_7900 ( .C ( clk ), .D ( signal_22592 ), .Q ( signal_22593 ) ) ;
    buf_clk cell_7908 ( .C ( clk ), .D ( signal_22600 ), .Q ( signal_22601 ) ) ;
    buf_clk cell_8276 ( .C ( clk ), .D ( signal_22968 ), .Q ( signal_22969 ) ) ;
    buf_clk cell_8286 ( .C ( clk ), .D ( signal_22978 ), .Q ( signal_22979 ) ) ;
    buf_clk cell_8296 ( .C ( clk ), .D ( signal_22988 ), .Q ( signal_22989 ) ) ;
    buf_clk cell_8306 ( .C ( clk ), .D ( signal_22998 ), .Q ( signal_22999 ) ) ;
    buf_clk cell_8316 ( .C ( clk ), .D ( signal_23008 ), .Q ( signal_23009 ) ) ;
    buf_clk cell_8716 ( .C ( clk ), .D ( signal_23408 ), .Q ( signal_23409 ) ) ;
    buf_clk cell_8728 ( .C ( clk ), .D ( signal_23420 ), .Q ( signal_23421 ) ) ;
    buf_clk cell_8740 ( .C ( clk ), .D ( signal_23432 ), .Q ( signal_23433 ) ) ;
    buf_clk cell_8752 ( .C ( clk ), .D ( signal_23444 ), .Q ( signal_23445 ) ) ;
    buf_clk cell_8764 ( .C ( clk ), .D ( signal_23456 ), .Q ( signal_23457 ) ) ;
    buf_clk cell_8838 ( .C ( clk ), .D ( signal_23530 ), .Q ( signal_23531 ) ) ;
    buf_clk cell_8852 ( .C ( clk ), .D ( signal_23544 ), .Q ( signal_23545 ) ) ;
    buf_clk cell_8866 ( .C ( clk ), .D ( signal_23558 ), .Q ( signal_23559 ) ) ;
    buf_clk cell_8880 ( .C ( clk ), .D ( signal_23572 ), .Q ( signal_23573 ) ) ;
    buf_clk cell_8894 ( .C ( clk ), .D ( signal_23586 ), .Q ( signal_23587 ) ) ;
    buf_clk cell_8948 ( .C ( clk ), .D ( signal_23640 ), .Q ( signal_23641 ) ) ;
    buf_clk cell_8962 ( .C ( clk ), .D ( signal_23654 ), .Q ( signal_23655 ) ) ;
    buf_clk cell_8976 ( .C ( clk ), .D ( signal_23668 ), .Q ( signal_23669 ) ) ;
    buf_clk cell_8990 ( .C ( clk ), .D ( signal_23682 ), .Q ( signal_23683 ) ) ;
    buf_clk cell_9004 ( .C ( clk ), .D ( signal_23696 ), .Q ( signal_23697 ) ) ;
    buf_clk cell_9148 ( .C ( clk ), .D ( signal_23840 ), .Q ( signal_23841 ) ) ;
    buf_clk cell_9164 ( .C ( clk ), .D ( signal_23856 ), .Q ( signal_23857 ) ) ;
    buf_clk cell_9180 ( .C ( clk ), .D ( signal_23872 ), .Q ( signal_23873 ) ) ;
    buf_clk cell_9196 ( .C ( clk ), .D ( signal_23888 ), .Q ( signal_23889 ) ) ;
    buf_clk cell_9212 ( .C ( clk ), .D ( signal_23904 ), .Q ( signal_23905 ) ) ;
    buf_clk cell_9248 ( .C ( clk ), .D ( signal_23940 ), .Q ( signal_23941 ) ) ;
    buf_clk cell_9264 ( .C ( clk ), .D ( signal_23956 ), .Q ( signal_23957 ) ) ;
    buf_clk cell_9280 ( .C ( clk ), .D ( signal_23972 ), .Q ( signal_23973 ) ) ;
    buf_clk cell_9296 ( .C ( clk ), .D ( signal_23988 ), .Q ( signal_23989 ) ) ;
    buf_clk cell_9312 ( .C ( clk ), .D ( signal_24004 ), .Q ( signal_24005 ) ) ;
    buf_clk cell_9556 ( .C ( clk ), .D ( signal_24248 ), .Q ( signal_24249 ) ) ;
    buf_clk cell_9572 ( .C ( clk ), .D ( signal_24264 ), .Q ( signal_24265 ) ) ;
    buf_clk cell_9588 ( .C ( clk ), .D ( signal_24280 ), .Q ( signal_24281 ) ) ;
    buf_clk cell_9604 ( .C ( clk ), .D ( signal_24296 ), .Q ( signal_24297 ) ) ;
    buf_clk cell_9620 ( .C ( clk ), .D ( signal_24312 ), .Q ( signal_24313 ) ) ;
    buf_clk cell_9638 ( .C ( clk ), .D ( signal_24330 ), .Q ( signal_24331 ) ) ;
    buf_clk cell_9656 ( .C ( clk ), .D ( signal_24348 ), .Q ( signal_24349 ) ) ;
    buf_clk cell_9674 ( .C ( clk ), .D ( signal_24366 ), .Q ( signal_24367 ) ) ;
    buf_clk cell_9692 ( .C ( clk ), .D ( signal_24384 ), .Q ( signal_24385 ) ) ;
    buf_clk cell_9710 ( .C ( clk ), .D ( signal_24402 ), .Q ( signal_24403 ) ) ;
    buf_clk cell_9888 ( .C ( clk ), .D ( signal_24580 ), .Q ( signal_24581 ) ) ;
    buf_clk cell_9908 ( .C ( clk ), .D ( signal_24600 ), .Q ( signal_24601 ) ) ;
    buf_clk cell_9928 ( .C ( clk ), .D ( signal_24620 ), .Q ( signal_24621 ) ) ;
    buf_clk cell_9948 ( .C ( clk ), .D ( signal_24640 ), .Q ( signal_24641 ) ) ;
    buf_clk cell_9968 ( .C ( clk ), .D ( signal_24660 ), .Q ( signal_24661 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_5911 ( .C ( clk ), .D ( signal_20603 ), .Q ( signal_20604 ) ) ;
    buf_clk cell_5919 ( .C ( clk ), .D ( signal_20611 ), .Q ( signal_20612 ) ) ;
    buf_clk cell_5927 ( .C ( clk ), .D ( signal_20619 ), .Q ( signal_20620 ) ) ;
    buf_clk cell_5935 ( .C ( clk ), .D ( signal_20627 ), .Q ( signal_20628 ) ) ;
    buf_clk cell_5943 ( .C ( clk ), .D ( signal_20635 ), .Q ( signal_20636 ) ) ;
    buf_clk cell_5947 ( .C ( clk ), .D ( signal_20639 ), .Q ( signal_20640 ) ) ;
    buf_clk cell_5951 ( .C ( clk ), .D ( signal_20643 ), .Q ( signal_20644 ) ) ;
    buf_clk cell_5955 ( .C ( clk ), .D ( signal_20647 ), .Q ( signal_20648 ) ) ;
    buf_clk cell_5959 ( .C ( clk ), .D ( signal_20651 ), .Q ( signal_20652 ) ) ;
    buf_clk cell_5963 ( .C ( clk ), .D ( signal_20655 ), .Q ( signal_20656 ) ) ;
    buf_clk cell_5969 ( .C ( clk ), .D ( signal_20661 ), .Q ( signal_20662 ) ) ;
    buf_clk cell_5975 ( .C ( clk ), .D ( signal_20667 ), .Q ( signal_20668 ) ) ;
    buf_clk cell_5981 ( .C ( clk ), .D ( signal_20673 ), .Q ( signal_20674 ) ) ;
    buf_clk cell_5987 ( .C ( clk ), .D ( signal_20679 ), .Q ( signal_20680 ) ) ;
    buf_clk cell_5993 ( .C ( clk ), .D ( signal_20685 ), .Q ( signal_20686 ) ) ;
    buf_clk cell_5999 ( .C ( clk ), .D ( signal_20691 ), .Q ( signal_20692 ) ) ;
    buf_clk cell_6005 ( .C ( clk ), .D ( signal_20697 ), .Q ( signal_20698 ) ) ;
    buf_clk cell_6011 ( .C ( clk ), .D ( signal_20703 ), .Q ( signal_20704 ) ) ;
    buf_clk cell_6017 ( .C ( clk ), .D ( signal_20709 ), .Q ( signal_20710 ) ) ;
    buf_clk cell_6023 ( .C ( clk ), .D ( signal_20715 ), .Q ( signal_20716 ) ) ;
    buf_clk cell_6027 ( .C ( clk ), .D ( signal_20719 ), .Q ( signal_20720 ) ) ;
    buf_clk cell_6031 ( .C ( clk ), .D ( signal_20723 ), .Q ( signal_20724 ) ) ;
    buf_clk cell_6035 ( .C ( clk ), .D ( signal_20727 ), .Q ( signal_20728 ) ) ;
    buf_clk cell_6039 ( .C ( clk ), .D ( signal_20731 ), .Q ( signal_20732 ) ) ;
    buf_clk cell_6043 ( .C ( clk ), .D ( signal_20735 ), .Q ( signal_20736 ) ) ;
    buf_clk cell_6049 ( .C ( clk ), .D ( signal_20741 ), .Q ( signal_20742 ) ) ;
    buf_clk cell_6055 ( .C ( clk ), .D ( signal_20747 ), .Q ( signal_20748 ) ) ;
    buf_clk cell_6061 ( .C ( clk ), .D ( signal_20753 ), .Q ( signal_20754 ) ) ;
    buf_clk cell_6067 ( .C ( clk ), .D ( signal_20759 ), .Q ( signal_20760 ) ) ;
    buf_clk cell_6073 ( .C ( clk ), .D ( signal_20765 ), .Q ( signal_20766 ) ) ;
    buf_clk cell_6077 ( .C ( clk ), .D ( signal_20769 ), .Q ( signal_20770 ) ) ;
    buf_clk cell_6081 ( .C ( clk ), .D ( signal_20773 ), .Q ( signal_20774 ) ) ;
    buf_clk cell_6085 ( .C ( clk ), .D ( signal_20777 ), .Q ( signal_20778 ) ) ;
    buf_clk cell_6089 ( .C ( clk ), .D ( signal_20781 ), .Q ( signal_20782 ) ) ;
    buf_clk cell_6093 ( .C ( clk ), .D ( signal_20785 ), .Q ( signal_20786 ) ) ;
    buf_clk cell_6097 ( .C ( clk ), .D ( signal_20789 ), .Q ( signal_20790 ) ) ;
    buf_clk cell_6101 ( .C ( clk ), .D ( signal_20793 ), .Q ( signal_20794 ) ) ;
    buf_clk cell_6105 ( .C ( clk ), .D ( signal_20797 ), .Q ( signal_20798 ) ) ;
    buf_clk cell_6109 ( .C ( clk ), .D ( signal_20801 ), .Q ( signal_20802 ) ) ;
    buf_clk cell_6113 ( .C ( clk ), .D ( signal_20805 ), .Q ( signal_20806 ) ) ;
    buf_clk cell_6115 ( .C ( clk ), .D ( signal_2071 ), .Q ( signal_20808 ) ) ;
    buf_clk cell_6117 ( .C ( clk ), .D ( signal_6940 ), .Q ( signal_20810 ) ) ;
    buf_clk cell_6119 ( .C ( clk ), .D ( signal_6941 ), .Q ( signal_20812 ) ) ;
    buf_clk cell_6121 ( .C ( clk ), .D ( signal_6942 ), .Q ( signal_20814 ) ) ;
    buf_clk cell_6123 ( .C ( clk ), .D ( signal_6943 ), .Q ( signal_20816 ) ) ;
    buf_clk cell_6125 ( .C ( clk ), .D ( signal_20199 ), .Q ( signal_20818 ) ) ;
    buf_clk cell_6127 ( .C ( clk ), .D ( signal_20201 ), .Q ( signal_20820 ) ) ;
    buf_clk cell_6129 ( .C ( clk ), .D ( signal_20203 ), .Q ( signal_20822 ) ) ;
    buf_clk cell_6131 ( .C ( clk ), .D ( signal_20205 ), .Q ( signal_20824 ) ) ;
    buf_clk cell_6133 ( .C ( clk ), .D ( signal_20207 ), .Q ( signal_20826 ) ) ;
    buf_clk cell_6139 ( .C ( clk ), .D ( signal_20831 ), .Q ( signal_20832 ) ) ;
    buf_clk cell_6145 ( .C ( clk ), .D ( signal_20837 ), .Q ( signal_20838 ) ) ;
    buf_clk cell_6151 ( .C ( clk ), .D ( signal_20843 ), .Q ( signal_20844 ) ) ;
    buf_clk cell_6157 ( .C ( clk ), .D ( signal_20849 ), .Q ( signal_20850 ) ) ;
    buf_clk cell_6163 ( .C ( clk ), .D ( signal_20855 ), .Q ( signal_20856 ) ) ;
    buf_clk cell_6169 ( .C ( clk ), .D ( signal_20861 ), .Q ( signal_20862 ) ) ;
    buf_clk cell_6175 ( .C ( clk ), .D ( signal_20867 ), .Q ( signal_20868 ) ) ;
    buf_clk cell_6181 ( .C ( clk ), .D ( signal_20873 ), .Q ( signal_20874 ) ) ;
    buf_clk cell_6187 ( .C ( clk ), .D ( signal_20879 ), .Q ( signal_20880 ) ) ;
    buf_clk cell_6193 ( .C ( clk ), .D ( signal_20885 ), .Q ( signal_20886 ) ) ;
    buf_clk cell_6199 ( .C ( clk ), .D ( signal_20891 ), .Q ( signal_20892 ) ) ;
    buf_clk cell_6205 ( .C ( clk ), .D ( signal_20897 ), .Q ( signal_20898 ) ) ;
    buf_clk cell_6211 ( .C ( clk ), .D ( signal_20903 ), .Q ( signal_20904 ) ) ;
    buf_clk cell_6217 ( .C ( clk ), .D ( signal_20909 ), .Q ( signal_20910 ) ) ;
    buf_clk cell_6223 ( .C ( clk ), .D ( signal_20915 ), .Q ( signal_20916 ) ) ;
    buf_clk cell_6225 ( .C ( clk ), .D ( signal_19871 ), .Q ( signal_20918 ) ) ;
    buf_clk cell_6227 ( .C ( clk ), .D ( signal_19875 ), .Q ( signal_20920 ) ) ;
    buf_clk cell_6229 ( .C ( clk ), .D ( signal_19879 ), .Q ( signal_20922 ) ) ;
    buf_clk cell_6231 ( .C ( clk ), .D ( signal_19883 ), .Q ( signal_20924 ) ) ;
    buf_clk cell_6233 ( .C ( clk ), .D ( signal_19887 ), .Q ( signal_20926 ) ) ;
    buf_clk cell_6237 ( .C ( clk ), .D ( signal_20929 ), .Q ( signal_20930 ) ) ;
    buf_clk cell_6241 ( .C ( clk ), .D ( signal_20933 ), .Q ( signal_20934 ) ) ;
    buf_clk cell_6245 ( .C ( clk ), .D ( signal_20937 ), .Q ( signal_20938 ) ) ;
    buf_clk cell_6249 ( .C ( clk ), .D ( signal_20941 ), .Q ( signal_20942 ) ) ;
    buf_clk cell_6253 ( .C ( clk ), .D ( signal_20945 ), .Q ( signal_20946 ) ) ;
    buf_clk cell_6259 ( .C ( clk ), .D ( signal_20951 ), .Q ( signal_20952 ) ) ;
    buf_clk cell_6265 ( .C ( clk ), .D ( signal_20957 ), .Q ( signal_20958 ) ) ;
    buf_clk cell_6271 ( .C ( clk ), .D ( signal_20963 ), .Q ( signal_20964 ) ) ;
    buf_clk cell_6277 ( .C ( clk ), .D ( signal_20969 ), .Q ( signal_20970 ) ) ;
    buf_clk cell_6283 ( .C ( clk ), .D ( signal_20975 ), .Q ( signal_20976 ) ) ;
    buf_clk cell_6285 ( .C ( clk ), .D ( signal_2081 ), .Q ( signal_20978 ) ) ;
    buf_clk cell_6287 ( .C ( clk ), .D ( signal_6980 ), .Q ( signal_20980 ) ) ;
    buf_clk cell_6289 ( .C ( clk ), .D ( signal_6981 ), .Q ( signal_20982 ) ) ;
    buf_clk cell_6291 ( .C ( clk ), .D ( signal_6982 ), .Q ( signal_20984 ) ) ;
    buf_clk cell_6293 ( .C ( clk ), .D ( signal_6983 ), .Q ( signal_20986 ) ) ;
    buf_clk cell_6299 ( .C ( clk ), .D ( signal_20991 ), .Q ( signal_20992 ) ) ;
    buf_clk cell_6305 ( .C ( clk ), .D ( signal_20997 ), .Q ( signal_20998 ) ) ;
    buf_clk cell_6311 ( .C ( clk ), .D ( signal_21003 ), .Q ( signal_21004 ) ) ;
    buf_clk cell_6317 ( .C ( clk ), .D ( signal_21009 ), .Q ( signal_21010 ) ) ;
    buf_clk cell_6323 ( .C ( clk ), .D ( signal_21015 ), .Q ( signal_21016 ) ) ;
    buf_clk cell_6325 ( .C ( clk ), .D ( signal_2069 ), .Q ( signal_21018 ) ) ;
    buf_clk cell_6327 ( .C ( clk ), .D ( signal_6932 ), .Q ( signal_21020 ) ) ;
    buf_clk cell_6329 ( .C ( clk ), .D ( signal_6933 ), .Q ( signal_21022 ) ) ;
    buf_clk cell_6331 ( .C ( clk ), .D ( signal_6934 ), .Q ( signal_21024 ) ) ;
    buf_clk cell_6333 ( .C ( clk ), .D ( signal_6935 ), .Q ( signal_21026 ) ) ;
    buf_clk cell_6341 ( .C ( clk ), .D ( signal_21033 ), .Q ( signal_21034 ) ) ;
    buf_clk cell_6349 ( .C ( clk ), .D ( signal_21041 ), .Q ( signal_21042 ) ) ;
    buf_clk cell_6357 ( .C ( clk ), .D ( signal_21049 ), .Q ( signal_21050 ) ) ;
    buf_clk cell_6365 ( .C ( clk ), .D ( signal_21057 ), .Q ( signal_21058 ) ) ;
    buf_clk cell_6373 ( .C ( clk ), .D ( signal_21065 ), .Q ( signal_21066 ) ) ;
    buf_clk cell_6377 ( .C ( clk ), .D ( signal_21069 ), .Q ( signal_21070 ) ) ;
    buf_clk cell_6381 ( .C ( clk ), .D ( signal_21073 ), .Q ( signal_21074 ) ) ;
    buf_clk cell_6385 ( .C ( clk ), .D ( signal_21077 ), .Q ( signal_21078 ) ) ;
    buf_clk cell_6389 ( .C ( clk ), .D ( signal_21081 ), .Q ( signal_21082 ) ) ;
    buf_clk cell_6393 ( .C ( clk ), .D ( signal_21085 ), .Q ( signal_21086 ) ) ;
    buf_clk cell_6397 ( .C ( clk ), .D ( signal_21089 ), .Q ( signal_21090 ) ) ;
    buf_clk cell_6401 ( .C ( clk ), .D ( signal_21093 ), .Q ( signal_21094 ) ) ;
    buf_clk cell_6405 ( .C ( clk ), .D ( signal_21097 ), .Q ( signal_21098 ) ) ;
    buf_clk cell_6409 ( .C ( clk ), .D ( signal_21101 ), .Q ( signal_21102 ) ) ;
    buf_clk cell_6413 ( .C ( clk ), .D ( signal_21105 ), .Q ( signal_21106 ) ) ;
    buf_clk cell_6419 ( .C ( clk ), .D ( signal_21111 ), .Q ( signal_21112 ) ) ;
    buf_clk cell_6425 ( .C ( clk ), .D ( signal_21117 ), .Q ( signal_21118 ) ) ;
    buf_clk cell_6431 ( .C ( clk ), .D ( signal_21123 ), .Q ( signal_21124 ) ) ;
    buf_clk cell_6437 ( .C ( clk ), .D ( signal_21129 ), .Q ( signal_21130 ) ) ;
    buf_clk cell_6443 ( .C ( clk ), .D ( signal_21135 ), .Q ( signal_21136 ) ) ;
    buf_clk cell_6449 ( .C ( clk ), .D ( signal_21141 ), .Q ( signal_21142 ) ) ;
    buf_clk cell_6455 ( .C ( clk ), .D ( signal_21147 ), .Q ( signal_21148 ) ) ;
    buf_clk cell_6461 ( .C ( clk ), .D ( signal_21153 ), .Q ( signal_21154 ) ) ;
    buf_clk cell_6467 ( .C ( clk ), .D ( signal_21159 ), .Q ( signal_21160 ) ) ;
    buf_clk cell_6473 ( .C ( clk ), .D ( signal_21165 ), .Q ( signal_21166 ) ) ;
    buf_clk cell_6477 ( .C ( clk ), .D ( signal_21169 ), .Q ( signal_21170 ) ) ;
    buf_clk cell_6481 ( .C ( clk ), .D ( signal_21173 ), .Q ( signal_21174 ) ) ;
    buf_clk cell_6485 ( .C ( clk ), .D ( signal_21177 ), .Q ( signal_21178 ) ) ;
    buf_clk cell_6489 ( .C ( clk ), .D ( signal_21181 ), .Q ( signal_21182 ) ) ;
    buf_clk cell_6493 ( .C ( clk ), .D ( signal_21185 ), .Q ( signal_21186 ) ) ;
    buf_clk cell_6501 ( .C ( clk ), .D ( signal_21193 ), .Q ( signal_21194 ) ) ;
    buf_clk cell_6509 ( .C ( clk ), .D ( signal_21201 ), .Q ( signal_21202 ) ) ;
    buf_clk cell_6517 ( .C ( clk ), .D ( signal_21209 ), .Q ( signal_21210 ) ) ;
    buf_clk cell_6525 ( .C ( clk ), .D ( signal_21217 ), .Q ( signal_21218 ) ) ;
    buf_clk cell_6533 ( .C ( clk ), .D ( signal_21225 ), .Q ( signal_21226 ) ) ;
    buf_clk cell_6539 ( .C ( clk ), .D ( signal_21231 ), .Q ( signal_21232 ) ) ;
    buf_clk cell_6545 ( .C ( clk ), .D ( signal_21237 ), .Q ( signal_21238 ) ) ;
    buf_clk cell_6551 ( .C ( clk ), .D ( signal_21243 ), .Q ( signal_21244 ) ) ;
    buf_clk cell_6557 ( .C ( clk ), .D ( signal_21249 ), .Q ( signal_21250 ) ) ;
    buf_clk cell_6563 ( .C ( clk ), .D ( signal_21255 ), .Q ( signal_21256 ) ) ;
    buf_clk cell_6569 ( .C ( clk ), .D ( signal_21261 ), .Q ( signal_21262 ) ) ;
    buf_clk cell_6575 ( .C ( clk ), .D ( signal_21267 ), .Q ( signal_21268 ) ) ;
    buf_clk cell_6581 ( .C ( clk ), .D ( signal_21273 ), .Q ( signal_21274 ) ) ;
    buf_clk cell_6587 ( .C ( clk ), .D ( signal_21279 ), .Q ( signal_21280 ) ) ;
    buf_clk cell_6593 ( .C ( clk ), .D ( signal_21285 ), .Q ( signal_21286 ) ) ;
    buf_clk cell_6595 ( .C ( clk ), .D ( signal_2201 ), .Q ( signal_21288 ) ) ;
    buf_clk cell_6597 ( .C ( clk ), .D ( signal_7460 ), .Q ( signal_21290 ) ) ;
    buf_clk cell_6599 ( .C ( clk ), .D ( signal_7461 ), .Q ( signal_21292 ) ) ;
    buf_clk cell_6601 ( .C ( clk ), .D ( signal_7462 ), .Q ( signal_21294 ) ) ;
    buf_clk cell_6603 ( .C ( clk ), .D ( signal_7463 ), .Q ( signal_21296 ) ) ;
    buf_clk cell_6605 ( .C ( clk ), .D ( signal_20059 ), .Q ( signal_21298 ) ) ;
    buf_clk cell_6607 ( .C ( clk ), .D ( signal_20061 ), .Q ( signal_21300 ) ) ;
    buf_clk cell_6609 ( .C ( clk ), .D ( signal_20063 ), .Q ( signal_21302 ) ) ;
    buf_clk cell_6611 ( .C ( clk ), .D ( signal_20065 ), .Q ( signal_21304 ) ) ;
    buf_clk cell_6613 ( .C ( clk ), .D ( signal_20067 ), .Q ( signal_21306 ) ) ;
    buf_clk cell_6619 ( .C ( clk ), .D ( signal_21311 ), .Q ( signal_21312 ) ) ;
    buf_clk cell_6625 ( .C ( clk ), .D ( signal_21317 ), .Q ( signal_21318 ) ) ;
    buf_clk cell_6631 ( .C ( clk ), .D ( signal_21323 ), .Q ( signal_21324 ) ) ;
    buf_clk cell_6637 ( .C ( clk ), .D ( signal_21329 ), .Q ( signal_21330 ) ) ;
    buf_clk cell_6643 ( .C ( clk ), .D ( signal_21335 ), .Q ( signal_21336 ) ) ;
    buf_clk cell_6645 ( .C ( clk ), .D ( signal_20049 ), .Q ( signal_21338 ) ) ;
    buf_clk cell_6647 ( .C ( clk ), .D ( signal_20051 ), .Q ( signal_21340 ) ) ;
    buf_clk cell_6649 ( .C ( clk ), .D ( signal_20053 ), .Q ( signal_21342 ) ) ;
    buf_clk cell_6651 ( .C ( clk ), .D ( signal_20055 ), .Q ( signal_21344 ) ) ;
    buf_clk cell_6653 ( .C ( clk ), .D ( signal_20057 ), .Q ( signal_21346 ) ) ;
    buf_clk cell_6655 ( .C ( clk ), .D ( signal_19603 ), .Q ( signal_21348 ) ) ;
    buf_clk cell_6657 ( .C ( clk ), .D ( signal_19609 ), .Q ( signal_21350 ) ) ;
    buf_clk cell_6659 ( .C ( clk ), .D ( signal_19615 ), .Q ( signal_21352 ) ) ;
    buf_clk cell_6661 ( .C ( clk ), .D ( signal_19621 ), .Q ( signal_21354 ) ) ;
    buf_clk cell_6663 ( .C ( clk ), .D ( signal_19627 ), .Q ( signal_21356 ) ) ;
    buf_clk cell_6669 ( .C ( clk ), .D ( signal_21361 ), .Q ( signal_21362 ) ) ;
    buf_clk cell_6675 ( .C ( clk ), .D ( signal_21367 ), .Q ( signal_21368 ) ) ;
    buf_clk cell_6681 ( .C ( clk ), .D ( signal_21373 ), .Q ( signal_21374 ) ) ;
    buf_clk cell_6687 ( .C ( clk ), .D ( signal_21379 ), .Q ( signal_21380 ) ) ;
    buf_clk cell_6693 ( .C ( clk ), .D ( signal_21385 ), .Q ( signal_21386 ) ) ;
    buf_clk cell_6699 ( .C ( clk ), .D ( signal_21391 ), .Q ( signal_21392 ) ) ;
    buf_clk cell_6705 ( .C ( clk ), .D ( signal_21397 ), .Q ( signal_21398 ) ) ;
    buf_clk cell_6711 ( .C ( clk ), .D ( signal_21403 ), .Q ( signal_21404 ) ) ;
    buf_clk cell_6717 ( .C ( clk ), .D ( signal_21409 ), .Q ( signal_21410 ) ) ;
    buf_clk cell_6723 ( .C ( clk ), .D ( signal_21415 ), .Q ( signal_21416 ) ) ;
    buf_clk cell_6727 ( .C ( clk ), .D ( signal_21419 ), .Q ( signal_21420 ) ) ;
    buf_clk cell_6731 ( .C ( clk ), .D ( signal_21423 ), .Q ( signal_21424 ) ) ;
    buf_clk cell_6735 ( .C ( clk ), .D ( signal_21427 ), .Q ( signal_21428 ) ) ;
    buf_clk cell_6739 ( .C ( clk ), .D ( signal_21431 ), .Q ( signal_21432 ) ) ;
    buf_clk cell_6743 ( .C ( clk ), .D ( signal_21435 ), .Q ( signal_21436 ) ) ;
    buf_clk cell_6751 ( .C ( clk ), .D ( signal_21443 ), .Q ( signal_21444 ) ) ;
    buf_clk cell_6761 ( .C ( clk ), .D ( signal_21453 ), .Q ( signal_21454 ) ) ;
    buf_clk cell_6771 ( .C ( clk ), .D ( signal_21463 ), .Q ( signal_21464 ) ) ;
    buf_clk cell_6781 ( .C ( clk ), .D ( signal_21473 ), .Q ( signal_21474 ) ) ;
    buf_clk cell_6791 ( .C ( clk ), .D ( signal_21483 ), .Q ( signal_21484 ) ) ;
    buf_clk cell_6797 ( .C ( clk ), .D ( signal_21489 ), .Q ( signal_21490 ) ) ;
    buf_clk cell_6803 ( .C ( clk ), .D ( signal_21495 ), .Q ( signal_21496 ) ) ;
    buf_clk cell_6809 ( .C ( clk ), .D ( signal_21501 ), .Q ( signal_21502 ) ) ;
    buf_clk cell_6815 ( .C ( clk ), .D ( signal_21507 ), .Q ( signal_21508 ) ) ;
    buf_clk cell_6821 ( .C ( clk ), .D ( signal_21513 ), .Q ( signal_21514 ) ) ;
    buf_clk cell_6829 ( .C ( clk ), .D ( signal_21521 ), .Q ( signal_21522 ) ) ;
    buf_clk cell_6837 ( .C ( clk ), .D ( signal_21529 ), .Q ( signal_21530 ) ) ;
    buf_clk cell_6845 ( .C ( clk ), .D ( signal_21537 ), .Q ( signal_21538 ) ) ;
    buf_clk cell_6853 ( .C ( clk ), .D ( signal_21545 ), .Q ( signal_21546 ) ) ;
    buf_clk cell_6861 ( .C ( clk ), .D ( signal_21553 ), .Q ( signal_21554 ) ) ;
    buf_clk cell_6869 ( .C ( clk ), .D ( signal_21561 ), .Q ( signal_21562 ) ) ;
    buf_clk cell_6877 ( .C ( clk ), .D ( signal_21569 ), .Q ( signal_21570 ) ) ;
    buf_clk cell_6885 ( .C ( clk ), .D ( signal_21577 ), .Q ( signal_21578 ) ) ;
    buf_clk cell_6893 ( .C ( clk ), .D ( signal_21585 ), .Q ( signal_21586 ) ) ;
    buf_clk cell_6901 ( .C ( clk ), .D ( signal_21593 ), .Q ( signal_21594 ) ) ;
    buf_clk cell_6905 ( .C ( clk ), .D ( signal_19979 ), .Q ( signal_21598 ) ) ;
    buf_clk cell_6909 ( .C ( clk ), .D ( signal_19981 ), .Q ( signal_21602 ) ) ;
    buf_clk cell_6913 ( .C ( clk ), .D ( signal_19983 ), .Q ( signal_21606 ) ) ;
    buf_clk cell_6917 ( .C ( clk ), .D ( signal_19985 ), .Q ( signal_21610 ) ) ;
    buf_clk cell_6921 ( .C ( clk ), .D ( signal_19987 ), .Q ( signal_21614 ) ) ;
    buf_clk cell_6925 ( .C ( clk ), .D ( signal_2116 ), .Q ( signal_21618 ) ) ;
    buf_clk cell_6929 ( .C ( clk ), .D ( signal_7120 ), .Q ( signal_21622 ) ) ;
    buf_clk cell_6933 ( .C ( clk ), .D ( signal_7121 ), .Q ( signal_21626 ) ) ;
    buf_clk cell_6937 ( .C ( clk ), .D ( signal_7122 ), .Q ( signal_21630 ) ) ;
    buf_clk cell_6941 ( .C ( clk ), .D ( signal_7123 ), .Q ( signal_21634 ) ) ;
    buf_clk cell_6965 ( .C ( clk ), .D ( signal_2109 ), .Q ( signal_21658 ) ) ;
    buf_clk cell_6969 ( .C ( clk ), .D ( signal_7092 ), .Q ( signal_21662 ) ) ;
    buf_clk cell_6973 ( .C ( clk ), .D ( signal_7093 ), .Q ( signal_21666 ) ) ;
    buf_clk cell_6977 ( .C ( clk ), .D ( signal_7094 ), .Q ( signal_21670 ) ) ;
    buf_clk cell_6981 ( .C ( clk ), .D ( signal_7095 ), .Q ( signal_21674 ) ) ;
    buf_clk cell_6991 ( .C ( clk ), .D ( signal_21683 ), .Q ( signal_21684 ) ) ;
    buf_clk cell_7001 ( .C ( clk ), .D ( signal_21693 ), .Q ( signal_21694 ) ) ;
    buf_clk cell_7011 ( .C ( clk ), .D ( signal_21703 ), .Q ( signal_21704 ) ) ;
    buf_clk cell_7021 ( .C ( clk ), .D ( signal_21713 ), .Q ( signal_21714 ) ) ;
    buf_clk cell_7031 ( .C ( clk ), .D ( signal_21723 ), .Q ( signal_21724 ) ) ;
    buf_clk cell_7037 ( .C ( clk ), .D ( signal_21729 ), .Q ( signal_21730 ) ) ;
    buf_clk cell_7043 ( .C ( clk ), .D ( signal_21735 ), .Q ( signal_21736 ) ) ;
    buf_clk cell_7049 ( .C ( clk ), .D ( signal_21741 ), .Q ( signal_21742 ) ) ;
    buf_clk cell_7055 ( .C ( clk ), .D ( signal_21747 ), .Q ( signal_21748 ) ) ;
    buf_clk cell_7061 ( .C ( clk ), .D ( signal_21753 ), .Q ( signal_21754 ) ) ;
    buf_clk cell_7079 ( .C ( clk ), .D ( signal_21771 ), .Q ( signal_21772 ) ) ;
    buf_clk cell_7087 ( .C ( clk ), .D ( signal_21779 ), .Q ( signal_21780 ) ) ;
    buf_clk cell_7095 ( .C ( clk ), .D ( signal_21787 ), .Q ( signal_21788 ) ) ;
    buf_clk cell_7103 ( .C ( clk ), .D ( signal_21795 ), .Q ( signal_21796 ) ) ;
    buf_clk cell_7111 ( .C ( clk ), .D ( signal_21803 ), .Q ( signal_21804 ) ) ;
    buf_clk cell_7117 ( .C ( clk ), .D ( signal_21809 ), .Q ( signal_21810 ) ) ;
    buf_clk cell_7123 ( .C ( clk ), .D ( signal_21815 ), .Q ( signal_21816 ) ) ;
    buf_clk cell_7129 ( .C ( clk ), .D ( signal_21821 ), .Q ( signal_21822 ) ) ;
    buf_clk cell_7135 ( .C ( clk ), .D ( signal_21827 ), .Q ( signal_21828 ) ) ;
    buf_clk cell_7141 ( .C ( clk ), .D ( signal_21833 ), .Q ( signal_21834 ) ) ;
    buf_clk cell_7149 ( .C ( clk ), .D ( signal_21841 ), .Q ( signal_21842 ) ) ;
    buf_clk cell_7157 ( .C ( clk ), .D ( signal_21849 ), .Q ( signal_21850 ) ) ;
    buf_clk cell_7165 ( .C ( clk ), .D ( signal_21857 ), .Q ( signal_21858 ) ) ;
    buf_clk cell_7173 ( .C ( clk ), .D ( signal_21865 ), .Q ( signal_21866 ) ) ;
    buf_clk cell_7181 ( .C ( clk ), .D ( signal_21873 ), .Q ( signal_21874 ) ) ;
    buf_clk cell_7189 ( .C ( clk ), .D ( signal_21881 ), .Q ( signal_21882 ) ) ;
    buf_clk cell_7197 ( .C ( clk ), .D ( signal_21889 ), .Q ( signal_21890 ) ) ;
    buf_clk cell_7205 ( .C ( clk ), .D ( signal_21897 ), .Q ( signal_21898 ) ) ;
    buf_clk cell_7213 ( .C ( clk ), .D ( signal_21905 ), .Q ( signal_21906 ) ) ;
    buf_clk cell_7221 ( .C ( clk ), .D ( signal_21913 ), .Q ( signal_21914 ) ) ;
    buf_clk cell_7229 ( .C ( clk ), .D ( signal_21921 ), .Q ( signal_21922 ) ) ;
    buf_clk cell_7237 ( .C ( clk ), .D ( signal_21929 ), .Q ( signal_21930 ) ) ;
    buf_clk cell_7245 ( .C ( clk ), .D ( signal_21937 ), .Q ( signal_21938 ) ) ;
    buf_clk cell_7253 ( .C ( clk ), .D ( signal_21945 ), .Q ( signal_21946 ) ) ;
    buf_clk cell_7261 ( .C ( clk ), .D ( signal_21953 ), .Q ( signal_21954 ) ) ;
    buf_clk cell_7271 ( .C ( clk ), .D ( signal_21963 ), .Q ( signal_21964 ) ) ;
    buf_clk cell_7281 ( .C ( clk ), .D ( signal_21973 ), .Q ( signal_21974 ) ) ;
    buf_clk cell_7291 ( .C ( clk ), .D ( signal_21983 ), .Q ( signal_21984 ) ) ;
    buf_clk cell_7301 ( .C ( clk ), .D ( signal_21993 ), .Q ( signal_21994 ) ) ;
    buf_clk cell_7311 ( .C ( clk ), .D ( signal_22003 ), .Q ( signal_22004 ) ) ;
    buf_clk cell_7319 ( .C ( clk ), .D ( signal_22011 ), .Q ( signal_22012 ) ) ;
    buf_clk cell_7327 ( .C ( clk ), .D ( signal_22019 ), .Q ( signal_22020 ) ) ;
    buf_clk cell_7335 ( .C ( clk ), .D ( signal_22027 ), .Q ( signal_22028 ) ) ;
    buf_clk cell_7343 ( .C ( clk ), .D ( signal_22035 ), .Q ( signal_22036 ) ) ;
    buf_clk cell_7351 ( .C ( clk ), .D ( signal_22043 ), .Q ( signal_22044 ) ) ;
    buf_clk cell_7359 ( .C ( clk ), .D ( signal_22051 ), .Q ( signal_22052 ) ) ;
    buf_clk cell_7367 ( .C ( clk ), .D ( signal_22059 ), .Q ( signal_22060 ) ) ;
    buf_clk cell_7375 ( .C ( clk ), .D ( signal_22067 ), .Q ( signal_22068 ) ) ;
    buf_clk cell_7383 ( .C ( clk ), .D ( signal_22075 ), .Q ( signal_22076 ) ) ;
    buf_clk cell_7391 ( .C ( clk ), .D ( signal_22083 ), .Q ( signal_22084 ) ) ;
    buf_clk cell_7409 ( .C ( clk ), .D ( signal_22101 ), .Q ( signal_22102 ) ) ;
    buf_clk cell_7417 ( .C ( clk ), .D ( signal_22109 ), .Q ( signal_22110 ) ) ;
    buf_clk cell_7425 ( .C ( clk ), .D ( signal_22117 ), .Q ( signal_22118 ) ) ;
    buf_clk cell_7433 ( .C ( clk ), .D ( signal_22125 ), .Q ( signal_22126 ) ) ;
    buf_clk cell_7441 ( .C ( clk ), .D ( signal_22133 ), .Q ( signal_22134 ) ) ;
    buf_clk cell_7449 ( .C ( clk ), .D ( signal_22141 ), .Q ( signal_22142 ) ) ;
    buf_clk cell_7457 ( .C ( clk ), .D ( signal_22149 ), .Q ( signal_22150 ) ) ;
    buf_clk cell_7465 ( .C ( clk ), .D ( signal_22157 ), .Q ( signal_22158 ) ) ;
    buf_clk cell_7473 ( .C ( clk ), .D ( signal_22165 ), .Q ( signal_22166 ) ) ;
    buf_clk cell_7481 ( .C ( clk ), .D ( signal_22173 ), .Q ( signal_22174 ) ) ;
    buf_clk cell_7489 ( .C ( clk ), .D ( signal_22181 ), .Q ( signal_22182 ) ) ;
    buf_clk cell_7497 ( .C ( clk ), .D ( signal_22189 ), .Q ( signal_22190 ) ) ;
    buf_clk cell_7505 ( .C ( clk ), .D ( signal_22197 ), .Q ( signal_22198 ) ) ;
    buf_clk cell_7513 ( .C ( clk ), .D ( signal_22205 ), .Q ( signal_22206 ) ) ;
    buf_clk cell_7521 ( .C ( clk ), .D ( signal_22213 ), .Q ( signal_22214 ) ) ;
    buf_clk cell_7525 ( .C ( clk ), .D ( signal_1945 ), .Q ( signal_22218 ) ) ;
    buf_clk cell_7531 ( .C ( clk ), .D ( signal_6436 ), .Q ( signal_22224 ) ) ;
    buf_clk cell_7537 ( .C ( clk ), .D ( signal_6437 ), .Q ( signal_22230 ) ) ;
    buf_clk cell_7543 ( .C ( clk ), .D ( signal_6438 ), .Q ( signal_22236 ) ) ;
    buf_clk cell_7549 ( .C ( clk ), .D ( signal_6439 ), .Q ( signal_22242 ) ) ;
    buf_clk cell_7557 ( .C ( clk ), .D ( signal_22249 ), .Q ( signal_22250 ) ) ;
    buf_clk cell_7565 ( .C ( clk ), .D ( signal_22257 ), .Q ( signal_22258 ) ) ;
    buf_clk cell_7573 ( .C ( clk ), .D ( signal_22265 ), .Q ( signal_22266 ) ) ;
    buf_clk cell_7581 ( .C ( clk ), .D ( signal_22273 ), .Q ( signal_22274 ) ) ;
    buf_clk cell_7589 ( .C ( clk ), .D ( signal_22281 ), .Q ( signal_22282 ) ) ;
    buf_clk cell_7595 ( .C ( clk ), .D ( signal_2111 ), .Q ( signal_22288 ) ) ;
    buf_clk cell_7601 ( .C ( clk ), .D ( signal_7100 ), .Q ( signal_22294 ) ) ;
    buf_clk cell_7607 ( .C ( clk ), .D ( signal_7101 ), .Q ( signal_22300 ) ) ;
    buf_clk cell_7613 ( .C ( clk ), .D ( signal_7102 ), .Q ( signal_22306 ) ) ;
    buf_clk cell_7619 ( .C ( clk ), .D ( signal_7103 ), .Q ( signal_22312 ) ) ;
    buf_clk cell_7625 ( .C ( clk ), .D ( signal_1976 ), .Q ( signal_22318 ) ) ;
    buf_clk cell_7631 ( .C ( clk ), .D ( signal_6560 ), .Q ( signal_22324 ) ) ;
    buf_clk cell_7637 ( .C ( clk ), .D ( signal_6561 ), .Q ( signal_22330 ) ) ;
    buf_clk cell_7643 ( .C ( clk ), .D ( signal_6562 ), .Q ( signal_22336 ) ) ;
    buf_clk cell_7649 ( .C ( clk ), .D ( signal_6563 ), .Q ( signal_22342 ) ) ;
    buf_clk cell_7657 ( .C ( clk ), .D ( signal_22349 ), .Q ( signal_22350 ) ) ;
    buf_clk cell_7665 ( .C ( clk ), .D ( signal_22357 ), .Q ( signal_22358 ) ) ;
    buf_clk cell_7673 ( .C ( clk ), .D ( signal_22365 ), .Q ( signal_22366 ) ) ;
    buf_clk cell_7681 ( .C ( clk ), .D ( signal_22373 ), .Q ( signal_22374 ) ) ;
    buf_clk cell_7689 ( .C ( clk ), .D ( signal_22381 ), .Q ( signal_22382 ) ) ;
    buf_clk cell_7699 ( .C ( clk ), .D ( signal_22391 ), .Q ( signal_22392 ) ) ;
    buf_clk cell_7709 ( .C ( clk ), .D ( signal_22401 ), .Q ( signal_22402 ) ) ;
    buf_clk cell_7719 ( .C ( clk ), .D ( signal_22411 ), .Q ( signal_22412 ) ) ;
    buf_clk cell_7729 ( .C ( clk ), .D ( signal_22421 ), .Q ( signal_22422 ) ) ;
    buf_clk cell_7739 ( .C ( clk ), .D ( signal_22431 ), .Q ( signal_22432 ) ) ;
    buf_clk cell_7755 ( .C ( clk ), .D ( signal_2070 ), .Q ( signal_22448 ) ) ;
    buf_clk cell_7761 ( .C ( clk ), .D ( signal_6936 ), .Q ( signal_22454 ) ) ;
    buf_clk cell_7767 ( .C ( clk ), .D ( signal_6937 ), .Q ( signal_22460 ) ) ;
    buf_clk cell_7773 ( .C ( clk ), .D ( signal_6938 ), .Q ( signal_22466 ) ) ;
    buf_clk cell_7779 ( .C ( clk ), .D ( signal_6939 ), .Q ( signal_22472 ) ) ;
    buf_clk cell_7787 ( .C ( clk ), .D ( signal_22479 ), .Q ( signal_22480 ) ) ;
    buf_clk cell_7795 ( .C ( clk ), .D ( signal_22487 ), .Q ( signal_22488 ) ) ;
    buf_clk cell_7803 ( .C ( clk ), .D ( signal_22495 ), .Q ( signal_22496 ) ) ;
    buf_clk cell_7811 ( .C ( clk ), .D ( signal_22503 ), .Q ( signal_22504 ) ) ;
    buf_clk cell_7819 ( .C ( clk ), .D ( signal_22511 ), .Q ( signal_22512 ) ) ;
    buf_clk cell_7829 ( .C ( clk ), .D ( signal_22521 ), .Q ( signal_22522 ) ) ;
    buf_clk cell_7839 ( .C ( clk ), .D ( signal_22531 ), .Q ( signal_22532 ) ) ;
    buf_clk cell_7849 ( .C ( clk ), .D ( signal_22541 ), .Q ( signal_22542 ) ) ;
    buf_clk cell_7859 ( .C ( clk ), .D ( signal_22551 ), .Q ( signal_22552 ) ) ;
    buf_clk cell_7869 ( .C ( clk ), .D ( signal_22561 ), .Q ( signal_22562 ) ) ;
    buf_clk cell_7877 ( .C ( clk ), .D ( signal_22569 ), .Q ( signal_22570 ) ) ;
    buf_clk cell_7885 ( .C ( clk ), .D ( signal_22577 ), .Q ( signal_22578 ) ) ;
    buf_clk cell_7893 ( .C ( clk ), .D ( signal_22585 ), .Q ( signal_22586 ) ) ;
    buf_clk cell_7901 ( .C ( clk ), .D ( signal_22593 ), .Q ( signal_22594 ) ) ;
    buf_clk cell_7909 ( .C ( clk ), .D ( signal_22601 ), .Q ( signal_22602 ) ) ;
    buf_clk cell_7915 ( .C ( clk ), .D ( signal_1890 ), .Q ( signal_22608 ) ) ;
    buf_clk cell_7921 ( .C ( clk ), .D ( signal_6216 ), .Q ( signal_22614 ) ) ;
    buf_clk cell_7927 ( .C ( clk ), .D ( signal_6217 ), .Q ( signal_22620 ) ) ;
    buf_clk cell_7933 ( .C ( clk ), .D ( signal_6218 ), .Q ( signal_22626 ) ) ;
    buf_clk cell_7939 ( .C ( clk ), .D ( signal_6219 ), .Q ( signal_22632 ) ) ;
    buf_clk cell_7945 ( .C ( clk ), .D ( signal_2002 ), .Q ( signal_22638 ) ) ;
    buf_clk cell_7951 ( .C ( clk ), .D ( signal_6664 ), .Q ( signal_22644 ) ) ;
    buf_clk cell_7957 ( .C ( clk ), .D ( signal_6665 ), .Q ( signal_22650 ) ) ;
    buf_clk cell_7963 ( .C ( clk ), .D ( signal_6666 ), .Q ( signal_22656 ) ) ;
    buf_clk cell_7969 ( .C ( clk ), .D ( signal_6667 ), .Q ( signal_22662 ) ) ;
    buf_clk cell_8025 ( .C ( clk ), .D ( signal_2106 ), .Q ( signal_22718 ) ) ;
    buf_clk cell_8031 ( .C ( clk ), .D ( signal_7080 ), .Q ( signal_22724 ) ) ;
    buf_clk cell_8037 ( .C ( clk ), .D ( signal_7081 ), .Q ( signal_22730 ) ) ;
    buf_clk cell_8043 ( .C ( clk ), .D ( signal_7082 ), .Q ( signal_22736 ) ) ;
    buf_clk cell_8049 ( .C ( clk ), .D ( signal_7083 ), .Q ( signal_22742 ) ) ;
    buf_clk cell_8065 ( .C ( clk ), .D ( signal_2068 ), .Q ( signal_22758 ) ) ;
    buf_clk cell_8071 ( .C ( clk ), .D ( signal_6928 ), .Q ( signal_22764 ) ) ;
    buf_clk cell_8077 ( .C ( clk ), .D ( signal_6929 ), .Q ( signal_22770 ) ) ;
    buf_clk cell_8083 ( .C ( clk ), .D ( signal_6930 ), .Q ( signal_22776 ) ) ;
    buf_clk cell_8089 ( .C ( clk ), .D ( signal_6931 ), .Q ( signal_22782 ) ) ;
    buf_clk cell_8115 ( .C ( clk ), .D ( signal_2073 ), .Q ( signal_22808 ) ) ;
    buf_clk cell_8121 ( .C ( clk ), .D ( signal_6948 ), .Q ( signal_22814 ) ) ;
    buf_clk cell_8127 ( .C ( clk ), .D ( signal_6949 ), .Q ( signal_22820 ) ) ;
    buf_clk cell_8133 ( .C ( clk ), .D ( signal_6950 ), .Q ( signal_22826 ) ) ;
    buf_clk cell_8139 ( .C ( clk ), .D ( signal_6951 ), .Q ( signal_22832 ) ) ;
    buf_clk cell_8205 ( .C ( clk ), .D ( signal_2110 ), .Q ( signal_22898 ) ) ;
    buf_clk cell_8213 ( .C ( clk ), .D ( signal_7096 ), .Q ( signal_22906 ) ) ;
    buf_clk cell_8221 ( .C ( clk ), .D ( signal_7097 ), .Q ( signal_22914 ) ) ;
    buf_clk cell_8229 ( .C ( clk ), .D ( signal_7098 ), .Q ( signal_22922 ) ) ;
    buf_clk cell_8237 ( .C ( clk ), .D ( signal_7099 ), .Q ( signal_22930 ) ) ;
    buf_clk cell_8277 ( .C ( clk ), .D ( signal_22969 ), .Q ( signal_22970 ) ) ;
    buf_clk cell_8287 ( .C ( clk ), .D ( signal_22979 ), .Q ( signal_22980 ) ) ;
    buf_clk cell_8297 ( .C ( clk ), .D ( signal_22989 ), .Q ( signal_22990 ) ) ;
    buf_clk cell_8307 ( .C ( clk ), .D ( signal_22999 ), .Q ( signal_23000 ) ) ;
    buf_clk cell_8317 ( .C ( clk ), .D ( signal_23009 ), .Q ( signal_23010 ) ) ;
    buf_clk cell_8375 ( .C ( clk ), .D ( signal_20101 ), .Q ( signal_23068 ) ) ;
    buf_clk cell_8383 ( .C ( clk ), .D ( signal_20105 ), .Q ( signal_23076 ) ) ;
    buf_clk cell_8391 ( .C ( clk ), .D ( signal_20109 ), .Q ( signal_23084 ) ) ;
    buf_clk cell_8399 ( .C ( clk ), .D ( signal_20113 ), .Q ( signal_23092 ) ) ;
    buf_clk cell_8407 ( .C ( clk ), .D ( signal_20117 ), .Q ( signal_23100 ) ) ;
    buf_clk cell_8445 ( .C ( clk ), .D ( signal_1986 ), .Q ( signal_23138 ) ) ;
    buf_clk cell_8453 ( .C ( clk ), .D ( signal_6600 ), .Q ( signal_23146 ) ) ;
    buf_clk cell_8461 ( .C ( clk ), .D ( signal_6601 ), .Q ( signal_23154 ) ) ;
    buf_clk cell_8469 ( .C ( clk ), .D ( signal_6602 ), .Q ( signal_23162 ) ) ;
    buf_clk cell_8477 ( .C ( clk ), .D ( signal_6603 ), .Q ( signal_23170 ) ) ;
    buf_clk cell_8515 ( .C ( clk ), .D ( signal_2082 ), .Q ( signal_23208 ) ) ;
    buf_clk cell_8523 ( .C ( clk ), .D ( signal_6984 ), .Q ( signal_23216 ) ) ;
    buf_clk cell_8531 ( .C ( clk ), .D ( signal_6985 ), .Q ( signal_23224 ) ) ;
    buf_clk cell_8539 ( .C ( clk ), .D ( signal_6986 ), .Q ( signal_23232 ) ) ;
    buf_clk cell_8547 ( .C ( clk ), .D ( signal_6987 ), .Q ( signal_23240 ) ) ;
    buf_clk cell_8717 ( .C ( clk ), .D ( signal_23409 ), .Q ( signal_23410 ) ) ;
    buf_clk cell_8729 ( .C ( clk ), .D ( signal_23421 ), .Q ( signal_23422 ) ) ;
    buf_clk cell_8741 ( .C ( clk ), .D ( signal_23433 ), .Q ( signal_23434 ) ) ;
    buf_clk cell_8753 ( .C ( clk ), .D ( signal_23445 ), .Q ( signal_23446 ) ) ;
    buf_clk cell_8765 ( .C ( clk ), .D ( signal_23457 ), .Q ( signal_23458 ) ) ;
    buf_clk cell_8839 ( .C ( clk ), .D ( signal_23531 ), .Q ( signal_23532 ) ) ;
    buf_clk cell_8853 ( .C ( clk ), .D ( signal_23545 ), .Q ( signal_23546 ) ) ;
    buf_clk cell_8867 ( .C ( clk ), .D ( signal_23559 ), .Q ( signal_23560 ) ) ;
    buf_clk cell_8881 ( .C ( clk ), .D ( signal_23573 ), .Q ( signal_23574 ) ) ;
    buf_clk cell_8895 ( .C ( clk ), .D ( signal_23587 ), .Q ( signal_23588 ) ) ;
    buf_clk cell_8949 ( .C ( clk ), .D ( signal_23641 ), .Q ( signal_23642 ) ) ;
    buf_clk cell_8963 ( .C ( clk ), .D ( signal_23655 ), .Q ( signal_23656 ) ) ;
    buf_clk cell_8977 ( .C ( clk ), .D ( signal_23669 ), .Q ( signal_23670 ) ) ;
    buf_clk cell_8991 ( .C ( clk ), .D ( signal_23683 ), .Q ( signal_23684 ) ) ;
    buf_clk cell_9005 ( .C ( clk ), .D ( signal_23697 ), .Q ( signal_23698 ) ) ;
    buf_clk cell_9149 ( .C ( clk ), .D ( signal_23841 ), .Q ( signal_23842 ) ) ;
    buf_clk cell_9165 ( .C ( clk ), .D ( signal_23857 ), .Q ( signal_23858 ) ) ;
    buf_clk cell_9181 ( .C ( clk ), .D ( signal_23873 ), .Q ( signal_23874 ) ) ;
    buf_clk cell_9197 ( .C ( clk ), .D ( signal_23889 ), .Q ( signal_23890 ) ) ;
    buf_clk cell_9213 ( .C ( clk ), .D ( signal_23905 ), .Q ( signal_23906 ) ) ;
    buf_clk cell_9249 ( .C ( clk ), .D ( signal_23941 ), .Q ( signal_23942 ) ) ;
    buf_clk cell_9265 ( .C ( clk ), .D ( signal_23957 ), .Q ( signal_23958 ) ) ;
    buf_clk cell_9281 ( .C ( clk ), .D ( signal_23973 ), .Q ( signal_23974 ) ) ;
    buf_clk cell_9297 ( .C ( clk ), .D ( signal_23989 ), .Q ( signal_23990 ) ) ;
    buf_clk cell_9313 ( .C ( clk ), .D ( signal_24005 ), .Q ( signal_24006 ) ) ;
    buf_clk cell_9557 ( .C ( clk ), .D ( signal_24249 ), .Q ( signal_24250 ) ) ;
    buf_clk cell_9573 ( .C ( clk ), .D ( signal_24265 ), .Q ( signal_24266 ) ) ;
    buf_clk cell_9589 ( .C ( clk ), .D ( signal_24281 ), .Q ( signal_24282 ) ) ;
    buf_clk cell_9605 ( .C ( clk ), .D ( signal_24297 ), .Q ( signal_24298 ) ) ;
    buf_clk cell_9621 ( .C ( clk ), .D ( signal_24313 ), .Q ( signal_24314 ) ) ;
    buf_clk cell_9639 ( .C ( clk ), .D ( signal_24331 ), .Q ( signal_24332 ) ) ;
    buf_clk cell_9657 ( .C ( clk ), .D ( signal_24349 ), .Q ( signal_24350 ) ) ;
    buf_clk cell_9675 ( .C ( clk ), .D ( signal_24367 ), .Q ( signal_24368 ) ) ;
    buf_clk cell_9693 ( .C ( clk ), .D ( signal_24385 ), .Q ( signal_24386 ) ) ;
    buf_clk cell_9711 ( .C ( clk ), .D ( signal_24403 ), .Q ( signal_24404 ) ) ;
    buf_clk cell_9889 ( .C ( clk ), .D ( signal_24581 ), .Q ( signal_24582 ) ) ;
    buf_clk cell_9909 ( .C ( clk ), .D ( signal_24601 ), .Q ( signal_24602 ) ) ;
    buf_clk cell_9929 ( .C ( clk ), .D ( signal_24621 ), .Q ( signal_24622 ) ) ;
    buf_clk cell_9949 ( .C ( clk ), .D ( signal_24641 ), .Q ( signal_24642 ) ) ;
    buf_clk cell_9969 ( .C ( clk ), .D ( signal_24661 ), .Q ( signal_24662 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2027 ( .a ({signal_19597, signal_19595, signal_19593, signal_19591, signal_19589}), .b ({signal_6363, signal_6362, signal_6361, signal_6360, signal_1926}), .clk ( clk ), .r ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650]}), .c ({signal_6827, signal_6826, signal_6825, signal_6824, signal_2042}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2032 ( .a ({signal_19627, signal_19621, signal_19615, signal_19609, signal_19603}), .b ({signal_6207, signal_6206, signal_6205, signal_6204, signal_1887}), .clk ( clk ), .r ({Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .c ({signal_6847, signal_6846, signal_6845, signal_6844, signal_2047}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2037 ( .a ({signal_19657, signal_19651, signal_19645, signal_19639, signal_19633}), .b ({signal_6419, signal_6418, signal_6417, signal_6416, signal_1940}), .clk ( clk ), .r ({Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670]}), .c ({signal_6867, signal_6866, signal_6865, signal_6864, signal_2052}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2038 ( .a ({signal_19687, signal_19681, signal_19675, signal_19669, signal_19663}), .b ({signal_6431, signal_6430, signal_6429, signal_6428, signal_1943}), .clk ( clk ), .r ({Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680]}), .c ({signal_6871, signal_6870, signal_6869, signal_6868, signal_2053}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2039 ( .a ({signal_19707, signal_19703, signal_19699, signal_19695, signal_19691}), .b ({signal_6443, signal_6442, signal_6441, signal_6440, signal_1946}), .clk ( clk ), .r ({Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690]}), .c ({signal_6875, signal_6874, signal_6873, signal_6872, signal_2054}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2040 ( .a ({signal_19737, signal_19731, signal_19725, signal_19719, signal_19713}), .b ({signal_6451, signal_6450, signal_6449, signal_6448, signal_1948}), .clk ( clk ), .r ({Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700]}), .c ({signal_6879, signal_6878, signal_6877, signal_6876, signal_2055}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2041 ( .a ({signal_19757, signal_19753, signal_19749, signal_19745, signal_19741}), .b ({signal_6459, signal_6458, signal_6457, signal_6456, signal_1950}), .clk ( clk ), .r ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710]}), .c ({signal_6883, signal_6882, signal_6881, signal_6880, signal_2056}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2042 ( .a ({signal_19777, signal_19773, signal_19769, signal_19765, signal_19761}), .b ({signal_6475, signal_6474, signal_6473, signal_6472, signal_1954}), .clk ( clk ), .r ({Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720]}), .c ({signal_6887, signal_6886, signal_6885, signal_6884, signal_2057}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2043 ( .a ({signal_19797, signal_19793, signal_19789, signal_19785, signal_19781}), .b ({signal_6479, signal_6478, signal_6477, signal_6476, signal_1955}), .clk ( clk ), .r ({Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730]}), .c ({signal_6891, signal_6890, signal_6889, signal_6888, signal_2058}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2044 ( .a ({signal_19817, signal_19813, signal_19809, signal_19805, signal_19801}), .b ({signal_6483, signal_6482, signal_6481, signal_6480, signal_1956}), .clk ( clk ), .r ({Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740]}), .c ({signal_6895, signal_6894, signal_6893, signal_6892, signal_2059}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2045 ( .a ({signal_19837, signal_19833, signal_19829, signal_19825, signal_19821}), .b ({signal_6503, signal_6502, signal_6501, signal_6500, signal_1961}), .clk ( clk ), .r ({Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750]}), .c ({signal_6899, signal_6898, signal_6897, signal_6896, signal_2060}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2064 ( .a ({signal_6827, signal_6826, signal_6825, signal_6824, signal_2042}), .b ({signal_6975, signal_6974, signal_6973, signal_6972, signal_2079}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2068 ( .a ({signal_6847, signal_6846, signal_6845, signal_6844, signal_2047}), .b ({signal_6991, signal_6990, signal_6989, signal_6988, signal_2083}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2072 ( .a ({signal_6867, signal_6866, signal_6865, signal_6864, signal_2052}), .b ({signal_7007, signal_7006, signal_7005, signal_7004, signal_2087}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2073 ( .a ({signal_6891, signal_6890, signal_6889, signal_6888, signal_2058}), .b ({signal_7011, signal_7010, signal_7009, signal_7008, signal_2088}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2084 ( .a ({signal_19867, signal_19861, signal_19855, signal_19849, signal_19843}), .b ({signal_6595, signal_6594, signal_6593, signal_6592, signal_1984}), .clk ( clk ), .r ({Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760]}), .c ({signal_7055, signal_7054, signal_7053, signal_7052, signal_2099}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2090 ( .a ({signal_19887, signal_19883, signal_19879, signal_19875, signal_19871}), .b ({signal_6631, signal_6630, signal_6629, signal_6628, signal_1993}), .clk ( clk ), .r ({Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770]}), .c ({signal_7079, signal_7078, signal_7077, signal_7076, signal_2105}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2098 ( .a ({signal_6391, signal_6390, signal_6389, signal_6388, signal_1933}), .b ({signal_19897, signal_19895, signal_19893, signal_19891, signal_19889}), .clk ( clk ), .r ({Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780]}), .c ({signal_7111, signal_7110, signal_7109, signal_7108, signal_2113}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2100 ( .a ({signal_19907, signal_19905, signal_19903, signal_19901, signal_19899}), .b ({signal_6663, signal_6662, signal_6661, signal_6660, signal_2001}), .clk ( clk ), .r ({Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790]}), .c ({signal_7119, signal_7118, signal_7117, signal_7116, signal_2115}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2102 ( .a ({signal_19917, signal_19915, signal_19913, signal_19911, signal_19909}), .b ({signal_6675, signal_6674, signal_6673, signal_6672, signal_2004}), .clk ( clk ), .r ({Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800]}), .c ({signal_7127, signal_7126, signal_7125, signal_7124, signal_2117}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2103 ( .a ({signal_19927, signal_19925, signal_19923, signal_19921, signal_19919}), .b ({signal_6423, signal_6422, signal_6421, signal_6420, signal_1941}), .clk ( clk ), .r ({Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810]}), .c ({signal_7131, signal_7130, signal_7129, signal_7128, signal_2118}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2105 ( .a ({signal_19937, signal_19935, signal_19933, signal_19931, signal_19929}), .b ({signal_6423, signal_6422, signal_6421, signal_6420, signal_1941}), .clk ( clk ), .r ({Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820]}), .c ({signal_7139, signal_7138, signal_7137, signal_7136, signal_2120}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2106 ( .a ({signal_19957, signal_19953, signal_19949, signal_19945, signal_19941}), .b ({signal_6819, signal_6818, signal_6817, signal_6816, signal_2040}), .clk ( clk ), .r ({Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830]}), .c ({signal_7143, signal_7142, signal_7141, signal_7140, signal_2121}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2107 ( .a ({signal_19967, signal_19965, signal_19963, signal_19961, signal_19959}), .b ({signal_6435, signal_6434, signal_6433, signal_6432, signal_1944}), .clk ( clk ), .r ({Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840]}), .c ({signal_7147, signal_7146, signal_7145, signal_7144, signal_2122}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2108 ( .a ({signal_19977, signal_19975, signal_19973, signal_19971, signal_19969}), .b ({signal_6839, signal_6838, signal_6837, signal_6836, signal_2045}), .clk ( clk ), .r ({Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850]}), .c ({signal_7151, signal_7150, signal_7149, signal_7148, signal_2123}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2109 ( .a ({signal_19987, signal_19985, signal_19983, signal_19981, signal_19979}), .b ({signal_6687, signal_6686, signal_6685, signal_6684, signal_2007}), .clk ( clk ), .r ({Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860]}), .c ({signal_7155, signal_7154, signal_7153, signal_7152, signal_2124}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2111 ( .a ({signal_20017, signal_20011, signal_20005, signal_19999, signal_19993}), .b ({signal_6691, signal_6690, signal_6689, signal_6688, signal_2008}), .clk ( clk ), .r ({Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870]}), .c ({signal_7163, signal_7162, signal_7161, signal_7160, signal_2126}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2112 ( .a ({signal_20027, signal_20025, signal_20023, signal_20021, signal_20019}), .b ({signal_6467, signal_6466, signal_6465, signal_6464, signal_1952}), .clk ( clk ), .r ({Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880]}), .c ({signal_7167, signal_7166, signal_7165, signal_7164, signal_2127}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2113 ( .a ({signal_20047, signal_20043, signal_20039, signal_20035, signal_20031}), .b ({signal_6855, signal_6854, signal_6853, signal_6852, signal_2049}), .clk ( clk ), .r ({Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890]}), .c ({signal_7171, signal_7170, signal_7169, signal_7168, signal_2128}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2114 ( .a ({signal_20057, signal_20055, signal_20053, signal_20051, signal_20049}), .b ({signal_6695, signal_6694, signal_6693, signal_6692, signal_2009}), .clk ( clk ), .r ({Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900]}), .c ({signal_7175, signal_7174, signal_7173, signal_7172, signal_2129}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2115 ( .a ({signal_19867, signal_19861, signal_19855, signal_19849, signal_19843}), .b ({signal_6699, signal_6698, signal_6697, signal_6696, signal_2010}), .clk ( clk ), .r ({Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910]}), .c ({signal_7179, signal_7178, signal_7177, signal_7176, signal_2130}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2117 ( .a ({signal_20067, signal_20065, signal_20063, signal_20061, signal_20059}), .b ({signal_6707, signal_6706, signal_6705, signal_6704, signal_2012}), .clk ( clk ), .r ({Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920]}), .c ({signal_7187, signal_7186, signal_7185, signal_7184, signal_2132}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2120 ( .a ({signal_19887, signal_19883, signal_19879, signal_19875, signal_19871}), .b ({signal_6711, signal_6710, signal_6709, signal_6708, signal_2013}), .clk ( clk ), .r ({Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930]}), .c ({signal_7199, signal_7198, signal_7197, signal_7196, signal_2135}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2129 ( .a ({signal_7055, signal_7054, signal_7053, signal_7052, signal_2099}), .b ({signal_7235, signal_7234, signal_7233, signal_7232, signal_2144}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2131 ( .a ({signal_7079, signal_7078, signal_7077, signal_7076, signal_2105}), .b ({signal_7243, signal_7242, signal_7241, signal_7240, signal_2146}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2132 ( .a ({signal_7119, signal_7118, signal_7117, signal_7116, signal_2115}), .b ({signal_7247, signal_7246, signal_7245, signal_7244, signal_2147}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2134 ( .a ({signal_7155, signal_7154, signal_7153, signal_7152, signal_2124}), .b ({signal_7255, signal_7254, signal_7253, signal_7252, signal_2149}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2136 ( .a ({signal_7163, signal_7162, signal_7161, signal_7160, signal_2126}), .b ({signal_7263, signal_7262, signal_7261, signal_7260, signal_2151}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2137 ( .a ({signal_7175, signal_7174, signal_7173, signal_7172, signal_2129}), .b ({signal_7267, signal_7266, signal_7265, signal_7264, signal_2152}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2138 ( .a ({signal_7179, signal_7178, signal_7177, signal_7176, signal_2130}), .b ({signal_7271, signal_7270, signal_7269, signal_7268, signal_2153}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2139 ( .a ({signal_7187, signal_7186, signal_7185, signal_7184, signal_2132}), .b ({signal_7275, signal_7274, signal_7273, signal_7272, signal_2154}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2141 ( .a ({signal_7199, signal_7198, signal_7197, signal_7196, signal_2135}), .b ({signal_7283, signal_7282, signal_7281, signal_7280, signal_2156}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2142 ( .a ({signal_20097, signal_20091, signal_20085, signal_20079, signal_20073}), .b ({signal_6903, signal_6902, signal_6901, signal_6900, signal_2061}), .clk ( clk ), .r ({Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940]}), .c ({signal_7287, signal_7286, signal_7285, signal_7284, signal_2157}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2143 ( .a ({signal_20117, signal_20113, signal_20109, signal_20105, signal_20101}), .b ({signal_6907, signal_6906, signal_6905, signal_6904, signal_2062}), .clk ( clk ), .r ({Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950]}), .c ({signal_7291, signal_7290, signal_7289, signal_7288, signal_2158}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2145 ( .a ({signal_20127, signal_20125, signal_20123, signal_20121, signal_20119}), .b ({signal_7019, signal_7018, signal_7017, signal_7016, signal_2090}), .clk ( clk ), .r ({Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960]}), .c ({signal_7299, signal_7298, signal_7297, signal_7296, signal_2160}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2146 ( .a ({signal_6919, signal_6918, signal_6917, signal_6916, signal_2065}), .b ({signal_20137, signal_20135, signal_20133, signal_20131, signal_20129}), .clk ( clk ), .r ({Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970]}), .c ({signal_7303, signal_7302, signal_7301, signal_7300, signal_2161}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2147 ( .a ({signal_20157, signal_20153, signal_20149, signal_20145, signal_20141}), .b ({signal_6923, signal_6922, signal_6921, signal_6920, signal_2066}), .clk ( clk ), .r ({Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980]}), .c ({signal_7307, signal_7306, signal_7305, signal_7304, signal_2162}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2149 ( .a ({signal_20177, signal_20173, signal_20169, signal_20165, signal_20161}), .b ({signal_7031, signal_7030, signal_7029, signal_7028, signal_2093}), .clk ( clk ), .r ({Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990]}), .c ({signal_7315, signal_7314, signal_7313, signal_7312, signal_2164}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2150 ( .a ({signal_20197, signal_20193, signal_20189, signal_20185, signal_20181}), .b ({signal_7035, signal_7034, signal_7033, signal_7032, signal_2094}), .clk ( clk ), .r ({Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000]}), .c ({signal_7319, signal_7318, signal_7317, signal_7316, signal_2165}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2151 ( .a ({signal_20207, signal_20205, signal_20203, signal_20201, signal_20199}), .b ({signal_6947, signal_6946, signal_6945, signal_6944, signal_2072}), .clk ( clk ), .r ({Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010]}), .c ({signal_7323, signal_7322, signal_7321, signal_7320, signal_2166}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2152 ( .a ({signal_20237, signal_20231, signal_20225, signal_20219, signal_20213}), .b ({signal_7039, signal_7038, signal_7037, signal_7036, signal_2095}), .clk ( clk ), .r ({Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020]}), .c ({signal_7327, signal_7326, signal_7325, signal_7324, signal_2167}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2153 ( .a ({signal_20257, signal_20253, signal_20249, signal_20245, signal_20241}), .b ({signal_7051, signal_7050, signal_7049, signal_7048, signal_2098}), .clk ( clk ), .r ({Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030]}), .c ({signal_7331, signal_7330, signal_7329, signal_7328, signal_2168}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2154 ( .a ({signal_20287, signal_20281, signal_20275, signal_20269, signal_20263}), .b ({signal_6959, signal_6958, signal_6957, signal_6956, signal_2075}), .clk ( clk ), .r ({Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040]}), .c ({signal_7335, signal_7334, signal_7333, signal_7332, signal_2169}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2155 ( .a ({signal_6915, signal_6914, signal_6913, signal_6912, signal_2064}), .b ({signal_6963, signal_6962, signal_6961, signal_6960, signal_2076}), .clk ( clk ), .r ({Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050]}), .c ({signal_7339, signal_7338, signal_7337, signal_7336, signal_2170}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2156 ( .a ({signal_20307, signal_20303, signal_20299, signal_20295, signal_20291}), .b ({signal_6967, signal_6966, signal_6965, signal_6964, signal_2077}), .clk ( clk ), .r ({Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060]}), .c ({signal_7343, signal_7342, signal_7341, signal_7340, signal_2171}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2157 ( .a ({signal_19627, signal_19621, signal_19615, signal_19609, signal_19603}), .b ({signal_6971, signal_6970, signal_6969, signal_6968, signal_2078}), .clk ( clk ), .r ({Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070]}), .c ({signal_7347, signal_7346, signal_7345, signal_7344, signal_2172}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2158 ( .a ({signal_20327, signal_20323, signal_20319, signal_20315, signal_20311}), .b ({signal_7059, signal_7058, signal_7057, signal_7056, signal_2100}), .clk ( clk ), .r ({Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080]}), .c ({signal_7351, signal_7350, signal_7349, signal_7348, signal_2173}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2159 ( .a ({signal_20347, signal_20343, signal_20339, signal_20335, signal_20331}), .b ({signal_7067, signal_7066, signal_7065, signal_7064, signal_2102}), .clk ( clk ), .r ({Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090]}), .c ({signal_7355, signal_7354, signal_7353, signal_7352, signal_2174}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2160 ( .a ({signal_20357, signal_20355, signal_20353, signal_20351, signal_20349}), .b ({signal_7071, signal_7070, signal_7069, signal_7068, signal_2103}), .clk ( clk ), .r ({Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100]}), .c ({signal_7359, signal_7358, signal_7357, signal_7356, signal_2175}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2161 ( .a ({signal_20377, signal_20373, signal_20369, signal_20365, signal_20361}), .b ({signal_7075, signal_7074, signal_7073, signal_7072, signal_2104}), .clk ( clk ), .r ({Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110]}), .c ({signal_7363, signal_7362, signal_7361, signal_7360, signal_2176}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2163 ( .a ({signal_20397, signal_20393, signal_20389, signal_20385, signal_20381}), .b ({signal_6979, signal_6978, signal_6977, signal_6976, signal_2080}), .clk ( clk ), .r ({Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120]}), .c ({signal_7371, signal_7370, signal_7369, signal_7368, signal_2178}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2164 ( .a ({signal_20427, signal_20421, signal_20415, signal_20409, signal_20403}), .b ({signal_7087, signal_7086, signal_7085, signal_7084, signal_2107}), .clk ( clk ), .r ({Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130]}), .c ({signal_7375, signal_7374, signal_7373, signal_7372, signal_2179}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2165 ( .a ({signal_7091, signal_7090, signal_7089, signal_7088, signal_2108}), .b ({signal_6471, signal_6470, signal_6469, signal_6468, signal_1953}), .clk ( clk ), .r ({Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140]}), .c ({signal_7379, signal_7378, signal_7377, signal_7376, signal_2180}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2166 ( .a ({signal_19627, signal_19621, signal_19615, signal_19609, signal_19603}), .b ({signal_6995, signal_6994, signal_6993, signal_6992, signal_2084}), .clk ( clk ), .r ({Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150]}), .c ({signal_7383, signal_7382, signal_7381, signal_7380, signal_2181}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2167 ( .a ({signal_6999, signal_6998, signal_6997, signal_6996, signal_2085}), .b ({signal_20437, signal_20435, signal_20433, signal_20431, signal_20429}), .clk ( clk ), .r ({Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160]}), .c ({signal_7387, signal_7386, signal_7385, signal_7384, signal_2182}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2168 ( .a ({signal_20447, signal_20445, signal_20443, signal_20441, signal_20439}), .b ({signal_7107, signal_7106, signal_7105, signal_7104, signal_2112}), .clk ( clk ), .r ({Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170]}), .c ({signal_7391, signal_7390, signal_7389, signal_7388, signal_2183}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2169 ( .a ({signal_20467, signal_20463, signal_20459, signal_20455, signal_20451}), .b ({signal_7003, signal_7002, signal_7001, signal_7000, signal_2086}), .clk ( clk ), .r ({Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180]}), .c ({signal_7395, signal_7394, signal_7393, signal_7392, signal_2184}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2171 ( .a ({signal_20497, signal_20491, signal_20485, signal_20479, signal_20473}), .b ({signal_7115, signal_7114, signal_7113, signal_7112, signal_2114}), .clk ( clk ), .r ({Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190]}), .c ({signal_7403, signal_7402, signal_7401, signal_7400, signal_2186}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2184 ( .a ({signal_7291, signal_7290, signal_7289, signal_7288, signal_2158}), .b ({signal_7455, signal_7454, signal_7453, signal_7452, signal_2199}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2187 ( .a ({signal_7323, signal_7322, signal_7321, signal_7320, signal_2166}), .b ({signal_7467, signal_7466, signal_7465, signal_7464, signal_2202}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2188 ( .a ({signal_7347, signal_7346, signal_7345, signal_7344, signal_2172}), .b ({signal_7471, signal_7470, signal_7469, signal_7468, signal_2203}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2189 ( .a ({signal_7355, signal_7354, signal_7353, signal_7352, signal_2174}), .b ({signal_7475, signal_7474, signal_7473, signal_7472, signal_2204}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2191 ( .a ({signal_7375, signal_7374, signal_7373, signal_7372, signal_2179}), .b ({signal_7483, signal_7482, signal_7481, signal_7480, signal_2206}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2192 ( .a ({signal_7379, signal_7378, signal_7377, signal_7376, signal_2180}), .b ({signal_7487, signal_7486, signal_7485, signal_7484, signal_2207}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2193 ( .a ({signal_7383, signal_7382, signal_7381, signal_7380, signal_2181}), .b ({signal_7491, signal_7490, signal_7489, signal_7488, signal_2208}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2194 ( .a ({signal_7403, signal_7402, signal_7401, signal_7400, signal_2186}), .b ({signal_7495, signal_7494, signal_7493, signal_7492, signal_2209}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2201 ( .a ({signal_20527, signal_20521, signal_20515, signal_20509, signal_20503}), .b ({signal_7215, signal_7214, signal_7213, signal_7212, signal_2139}), .clk ( clk ), .r ({Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200]}), .c ({signal_7523, signal_7522, signal_7521, signal_7520, signal_2216}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2202 ( .a ({signal_20557, signal_20551, signal_20545, signal_20539, signal_20533}), .b ({signal_7219, signal_7218, signal_7217, signal_7216, signal_2140}), .clk ( clk ), .r ({Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210]}), .c ({signal_7527, signal_7526, signal_7525, signal_7524, signal_2217}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2203 ( .a ({signal_20577, signal_20573, signal_20569, signal_20565, signal_20561}), .b ({signal_7223, signal_7222, signal_7221, signal_7220, signal_2141}), .clk ( clk ), .r ({Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220]}), .c ({signal_7531, signal_7530, signal_7529, signal_7528, signal_2218}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2204 ( .a ({signal_19627, signal_19621, signal_19615, signal_19609, signal_19603}), .b ({signal_7227, signal_7226, signal_7225, signal_7224, signal_2142}), .clk ( clk ), .r ({Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230]}), .c ({signal_7535, signal_7534, signal_7533, signal_7532, signal_2219}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2205 ( .a ({signal_20587, signal_20585, signal_20583, signal_20581, signal_20579}), .b ({signal_7231, signal_7230, signal_7229, signal_7228, signal_2143}), .clk ( clk ), .r ({Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240]}), .c ({signal_7539, signal_7538, signal_7537, signal_7536, signal_2220}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2206 ( .a ({signal_20057, signal_20055, signal_20053, signal_20051, signal_20049}), .b ({signal_7239, signal_7238, signal_7237, signal_7236, signal_2145}), .clk ( clk ), .r ({Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250]}), .c ({signal_7543, signal_7542, signal_7541, signal_7540, signal_2221}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2213 ( .a ({signal_20597, signal_20595, signal_20593, signal_20591, signal_20589}), .b ({signal_7251, signal_7250, signal_7249, signal_7248, signal_2148}), .clk ( clk ), .r ({Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260]}), .c ({signal_7571, signal_7570, signal_7569, signal_7568, signal_2228}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2221 ( .a ({signal_20557, signal_20551, signal_20545, signal_20539, signal_20533}), .b ({signal_7259, signal_7258, signal_7257, signal_7256, signal_2150}), .clk ( clk ), .r ({Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270]}), .c ({signal_7603, signal_7602, signal_7601, signal_7600, signal_2236}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2233 ( .a ({signal_7523, signal_7522, signal_7521, signal_7520, signal_2216}), .b ({signal_7651, signal_7650, signal_7649, signal_7648, signal_2248}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2234 ( .a ({signal_7527, signal_7526, signal_7525, signal_7524, signal_2217}), .b ({signal_7655, signal_7654, signal_7653, signal_7652, signal_2249}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2235 ( .a ({signal_7531, signal_7530, signal_7529, signal_7528, signal_2218}), .b ({signal_7659, signal_7658, signal_7657, signal_7656, signal_2250}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2236 ( .a ({signal_7535, signal_7534, signal_7533, signal_7532, signal_2219}), .b ({signal_7663, signal_7662, signal_7661, signal_7660, signal_2251}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2237 ( .a ({signal_7539, signal_7538, signal_7537, signal_7536, signal_2220}), .b ({signal_7667, signal_7666, signal_7665, signal_7664, signal_2252}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2238 ( .a ({signal_7543, signal_7542, signal_7541, signal_7540, signal_2221}), .b ({signal_7671, signal_7670, signal_7669, signal_7668, signal_2253}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2240 ( .a ({signal_7571, signal_7570, signal_7569, signal_7568, signal_2228}), .b ({signal_7679, signal_7678, signal_7677, signal_7676, signal_2255}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2242 ( .a ({signal_7603, signal_7602, signal_7601, signal_7600, signal_2236}), .b ({signal_7687, signal_7686, signal_7685, signal_7684, signal_2257}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2248 ( .a ({signal_6955, signal_6954, signal_6953, signal_6952, signal_2074}), .b ({signal_7459, signal_7458, signal_7457, signal_7456, signal_2200}), .clk ( clk ), .r ({Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280]}), .c ({signal_7711, signal_7710, signal_7709, signal_7708, signal_2263}) ) ;
    buf_clk cell_5912 ( .C ( clk ), .D ( signal_20604 ), .Q ( signal_20605 ) ) ;
    buf_clk cell_5920 ( .C ( clk ), .D ( signal_20612 ), .Q ( signal_20613 ) ) ;
    buf_clk cell_5928 ( .C ( clk ), .D ( signal_20620 ), .Q ( signal_20621 ) ) ;
    buf_clk cell_5936 ( .C ( clk ), .D ( signal_20628 ), .Q ( signal_20629 ) ) ;
    buf_clk cell_5944 ( .C ( clk ), .D ( signal_20636 ), .Q ( signal_20637 ) ) ;
    buf_clk cell_5948 ( .C ( clk ), .D ( signal_20640 ), .Q ( signal_20641 ) ) ;
    buf_clk cell_5952 ( .C ( clk ), .D ( signal_20644 ), .Q ( signal_20645 ) ) ;
    buf_clk cell_5956 ( .C ( clk ), .D ( signal_20648 ), .Q ( signal_20649 ) ) ;
    buf_clk cell_5960 ( .C ( clk ), .D ( signal_20652 ), .Q ( signal_20653 ) ) ;
    buf_clk cell_5964 ( .C ( clk ), .D ( signal_20656 ), .Q ( signal_20657 ) ) ;
    buf_clk cell_5970 ( .C ( clk ), .D ( signal_20662 ), .Q ( signal_20663 ) ) ;
    buf_clk cell_5976 ( .C ( clk ), .D ( signal_20668 ), .Q ( signal_20669 ) ) ;
    buf_clk cell_5982 ( .C ( clk ), .D ( signal_20674 ), .Q ( signal_20675 ) ) ;
    buf_clk cell_5988 ( .C ( clk ), .D ( signal_20680 ), .Q ( signal_20681 ) ) ;
    buf_clk cell_5994 ( .C ( clk ), .D ( signal_20686 ), .Q ( signal_20687 ) ) ;
    buf_clk cell_6000 ( .C ( clk ), .D ( signal_20692 ), .Q ( signal_20693 ) ) ;
    buf_clk cell_6006 ( .C ( clk ), .D ( signal_20698 ), .Q ( signal_20699 ) ) ;
    buf_clk cell_6012 ( .C ( clk ), .D ( signal_20704 ), .Q ( signal_20705 ) ) ;
    buf_clk cell_6018 ( .C ( clk ), .D ( signal_20710 ), .Q ( signal_20711 ) ) ;
    buf_clk cell_6024 ( .C ( clk ), .D ( signal_20716 ), .Q ( signal_20717 ) ) ;
    buf_clk cell_6028 ( .C ( clk ), .D ( signal_20720 ), .Q ( signal_20721 ) ) ;
    buf_clk cell_6032 ( .C ( clk ), .D ( signal_20724 ), .Q ( signal_20725 ) ) ;
    buf_clk cell_6036 ( .C ( clk ), .D ( signal_20728 ), .Q ( signal_20729 ) ) ;
    buf_clk cell_6040 ( .C ( clk ), .D ( signal_20732 ), .Q ( signal_20733 ) ) ;
    buf_clk cell_6044 ( .C ( clk ), .D ( signal_20736 ), .Q ( signal_20737 ) ) ;
    buf_clk cell_6050 ( .C ( clk ), .D ( signal_20742 ), .Q ( signal_20743 ) ) ;
    buf_clk cell_6056 ( .C ( clk ), .D ( signal_20748 ), .Q ( signal_20749 ) ) ;
    buf_clk cell_6062 ( .C ( clk ), .D ( signal_20754 ), .Q ( signal_20755 ) ) ;
    buf_clk cell_6068 ( .C ( clk ), .D ( signal_20760 ), .Q ( signal_20761 ) ) ;
    buf_clk cell_6074 ( .C ( clk ), .D ( signal_20766 ), .Q ( signal_20767 ) ) ;
    buf_clk cell_6078 ( .C ( clk ), .D ( signal_20770 ), .Q ( signal_20771 ) ) ;
    buf_clk cell_6082 ( .C ( clk ), .D ( signal_20774 ), .Q ( signal_20775 ) ) ;
    buf_clk cell_6086 ( .C ( clk ), .D ( signal_20778 ), .Q ( signal_20779 ) ) ;
    buf_clk cell_6090 ( .C ( clk ), .D ( signal_20782 ), .Q ( signal_20783 ) ) ;
    buf_clk cell_6094 ( .C ( clk ), .D ( signal_20786 ), .Q ( signal_20787 ) ) ;
    buf_clk cell_6098 ( .C ( clk ), .D ( signal_20790 ), .Q ( signal_20791 ) ) ;
    buf_clk cell_6102 ( .C ( clk ), .D ( signal_20794 ), .Q ( signal_20795 ) ) ;
    buf_clk cell_6106 ( .C ( clk ), .D ( signal_20798 ), .Q ( signal_20799 ) ) ;
    buf_clk cell_6110 ( .C ( clk ), .D ( signal_20802 ), .Q ( signal_20803 ) ) ;
    buf_clk cell_6114 ( .C ( clk ), .D ( signal_20806 ), .Q ( signal_20807 ) ) ;
    buf_clk cell_6116 ( .C ( clk ), .D ( signal_20808 ), .Q ( signal_20809 ) ) ;
    buf_clk cell_6118 ( .C ( clk ), .D ( signal_20810 ), .Q ( signal_20811 ) ) ;
    buf_clk cell_6120 ( .C ( clk ), .D ( signal_20812 ), .Q ( signal_20813 ) ) ;
    buf_clk cell_6122 ( .C ( clk ), .D ( signal_20814 ), .Q ( signal_20815 ) ) ;
    buf_clk cell_6124 ( .C ( clk ), .D ( signal_20816 ), .Q ( signal_20817 ) ) ;
    buf_clk cell_6126 ( .C ( clk ), .D ( signal_20818 ), .Q ( signal_20819 ) ) ;
    buf_clk cell_6128 ( .C ( clk ), .D ( signal_20820 ), .Q ( signal_20821 ) ) ;
    buf_clk cell_6130 ( .C ( clk ), .D ( signal_20822 ), .Q ( signal_20823 ) ) ;
    buf_clk cell_6132 ( .C ( clk ), .D ( signal_20824 ), .Q ( signal_20825 ) ) ;
    buf_clk cell_6134 ( .C ( clk ), .D ( signal_20826 ), .Q ( signal_20827 ) ) ;
    buf_clk cell_6140 ( .C ( clk ), .D ( signal_20832 ), .Q ( signal_20833 ) ) ;
    buf_clk cell_6146 ( .C ( clk ), .D ( signal_20838 ), .Q ( signal_20839 ) ) ;
    buf_clk cell_6152 ( .C ( clk ), .D ( signal_20844 ), .Q ( signal_20845 ) ) ;
    buf_clk cell_6158 ( .C ( clk ), .D ( signal_20850 ), .Q ( signal_20851 ) ) ;
    buf_clk cell_6164 ( .C ( clk ), .D ( signal_20856 ), .Q ( signal_20857 ) ) ;
    buf_clk cell_6170 ( .C ( clk ), .D ( signal_20862 ), .Q ( signal_20863 ) ) ;
    buf_clk cell_6176 ( .C ( clk ), .D ( signal_20868 ), .Q ( signal_20869 ) ) ;
    buf_clk cell_6182 ( .C ( clk ), .D ( signal_20874 ), .Q ( signal_20875 ) ) ;
    buf_clk cell_6188 ( .C ( clk ), .D ( signal_20880 ), .Q ( signal_20881 ) ) ;
    buf_clk cell_6194 ( .C ( clk ), .D ( signal_20886 ), .Q ( signal_20887 ) ) ;
    buf_clk cell_6200 ( .C ( clk ), .D ( signal_20892 ), .Q ( signal_20893 ) ) ;
    buf_clk cell_6206 ( .C ( clk ), .D ( signal_20898 ), .Q ( signal_20899 ) ) ;
    buf_clk cell_6212 ( .C ( clk ), .D ( signal_20904 ), .Q ( signal_20905 ) ) ;
    buf_clk cell_6218 ( .C ( clk ), .D ( signal_20910 ), .Q ( signal_20911 ) ) ;
    buf_clk cell_6224 ( .C ( clk ), .D ( signal_20916 ), .Q ( signal_20917 ) ) ;
    buf_clk cell_6226 ( .C ( clk ), .D ( signal_20918 ), .Q ( signal_20919 ) ) ;
    buf_clk cell_6228 ( .C ( clk ), .D ( signal_20920 ), .Q ( signal_20921 ) ) ;
    buf_clk cell_6230 ( .C ( clk ), .D ( signal_20922 ), .Q ( signal_20923 ) ) ;
    buf_clk cell_6232 ( .C ( clk ), .D ( signal_20924 ), .Q ( signal_20925 ) ) ;
    buf_clk cell_6234 ( .C ( clk ), .D ( signal_20926 ), .Q ( signal_20927 ) ) ;
    buf_clk cell_6238 ( .C ( clk ), .D ( signal_20930 ), .Q ( signal_20931 ) ) ;
    buf_clk cell_6242 ( .C ( clk ), .D ( signal_20934 ), .Q ( signal_20935 ) ) ;
    buf_clk cell_6246 ( .C ( clk ), .D ( signal_20938 ), .Q ( signal_20939 ) ) ;
    buf_clk cell_6250 ( .C ( clk ), .D ( signal_20942 ), .Q ( signal_20943 ) ) ;
    buf_clk cell_6254 ( .C ( clk ), .D ( signal_20946 ), .Q ( signal_20947 ) ) ;
    buf_clk cell_6260 ( .C ( clk ), .D ( signal_20952 ), .Q ( signal_20953 ) ) ;
    buf_clk cell_6266 ( .C ( clk ), .D ( signal_20958 ), .Q ( signal_20959 ) ) ;
    buf_clk cell_6272 ( .C ( clk ), .D ( signal_20964 ), .Q ( signal_20965 ) ) ;
    buf_clk cell_6278 ( .C ( clk ), .D ( signal_20970 ), .Q ( signal_20971 ) ) ;
    buf_clk cell_6284 ( .C ( clk ), .D ( signal_20976 ), .Q ( signal_20977 ) ) ;
    buf_clk cell_6286 ( .C ( clk ), .D ( signal_20978 ), .Q ( signal_20979 ) ) ;
    buf_clk cell_6288 ( .C ( clk ), .D ( signal_20980 ), .Q ( signal_20981 ) ) ;
    buf_clk cell_6290 ( .C ( clk ), .D ( signal_20982 ), .Q ( signal_20983 ) ) ;
    buf_clk cell_6292 ( .C ( clk ), .D ( signal_20984 ), .Q ( signal_20985 ) ) ;
    buf_clk cell_6294 ( .C ( clk ), .D ( signal_20986 ), .Q ( signal_20987 ) ) ;
    buf_clk cell_6300 ( .C ( clk ), .D ( signal_20992 ), .Q ( signal_20993 ) ) ;
    buf_clk cell_6306 ( .C ( clk ), .D ( signal_20998 ), .Q ( signal_20999 ) ) ;
    buf_clk cell_6312 ( .C ( clk ), .D ( signal_21004 ), .Q ( signal_21005 ) ) ;
    buf_clk cell_6318 ( .C ( clk ), .D ( signal_21010 ), .Q ( signal_21011 ) ) ;
    buf_clk cell_6324 ( .C ( clk ), .D ( signal_21016 ), .Q ( signal_21017 ) ) ;
    buf_clk cell_6326 ( .C ( clk ), .D ( signal_21018 ), .Q ( signal_21019 ) ) ;
    buf_clk cell_6328 ( .C ( clk ), .D ( signal_21020 ), .Q ( signal_21021 ) ) ;
    buf_clk cell_6330 ( .C ( clk ), .D ( signal_21022 ), .Q ( signal_21023 ) ) ;
    buf_clk cell_6332 ( .C ( clk ), .D ( signal_21024 ), .Q ( signal_21025 ) ) ;
    buf_clk cell_6334 ( .C ( clk ), .D ( signal_21026 ), .Q ( signal_21027 ) ) ;
    buf_clk cell_6342 ( .C ( clk ), .D ( signal_21034 ), .Q ( signal_21035 ) ) ;
    buf_clk cell_6350 ( .C ( clk ), .D ( signal_21042 ), .Q ( signal_21043 ) ) ;
    buf_clk cell_6358 ( .C ( clk ), .D ( signal_21050 ), .Q ( signal_21051 ) ) ;
    buf_clk cell_6366 ( .C ( clk ), .D ( signal_21058 ), .Q ( signal_21059 ) ) ;
    buf_clk cell_6374 ( .C ( clk ), .D ( signal_21066 ), .Q ( signal_21067 ) ) ;
    buf_clk cell_6378 ( .C ( clk ), .D ( signal_21070 ), .Q ( signal_21071 ) ) ;
    buf_clk cell_6382 ( .C ( clk ), .D ( signal_21074 ), .Q ( signal_21075 ) ) ;
    buf_clk cell_6386 ( .C ( clk ), .D ( signal_21078 ), .Q ( signal_21079 ) ) ;
    buf_clk cell_6390 ( .C ( clk ), .D ( signal_21082 ), .Q ( signal_21083 ) ) ;
    buf_clk cell_6394 ( .C ( clk ), .D ( signal_21086 ), .Q ( signal_21087 ) ) ;
    buf_clk cell_6398 ( .C ( clk ), .D ( signal_21090 ), .Q ( signal_21091 ) ) ;
    buf_clk cell_6402 ( .C ( clk ), .D ( signal_21094 ), .Q ( signal_21095 ) ) ;
    buf_clk cell_6406 ( .C ( clk ), .D ( signal_21098 ), .Q ( signal_21099 ) ) ;
    buf_clk cell_6410 ( .C ( clk ), .D ( signal_21102 ), .Q ( signal_21103 ) ) ;
    buf_clk cell_6414 ( .C ( clk ), .D ( signal_21106 ), .Q ( signal_21107 ) ) ;
    buf_clk cell_6420 ( .C ( clk ), .D ( signal_21112 ), .Q ( signal_21113 ) ) ;
    buf_clk cell_6426 ( .C ( clk ), .D ( signal_21118 ), .Q ( signal_21119 ) ) ;
    buf_clk cell_6432 ( .C ( clk ), .D ( signal_21124 ), .Q ( signal_21125 ) ) ;
    buf_clk cell_6438 ( .C ( clk ), .D ( signal_21130 ), .Q ( signal_21131 ) ) ;
    buf_clk cell_6444 ( .C ( clk ), .D ( signal_21136 ), .Q ( signal_21137 ) ) ;
    buf_clk cell_6450 ( .C ( clk ), .D ( signal_21142 ), .Q ( signal_21143 ) ) ;
    buf_clk cell_6456 ( .C ( clk ), .D ( signal_21148 ), .Q ( signal_21149 ) ) ;
    buf_clk cell_6462 ( .C ( clk ), .D ( signal_21154 ), .Q ( signal_21155 ) ) ;
    buf_clk cell_6468 ( .C ( clk ), .D ( signal_21160 ), .Q ( signal_21161 ) ) ;
    buf_clk cell_6474 ( .C ( clk ), .D ( signal_21166 ), .Q ( signal_21167 ) ) ;
    buf_clk cell_6478 ( .C ( clk ), .D ( signal_21170 ), .Q ( signal_21171 ) ) ;
    buf_clk cell_6482 ( .C ( clk ), .D ( signal_21174 ), .Q ( signal_21175 ) ) ;
    buf_clk cell_6486 ( .C ( clk ), .D ( signal_21178 ), .Q ( signal_21179 ) ) ;
    buf_clk cell_6490 ( .C ( clk ), .D ( signal_21182 ), .Q ( signal_21183 ) ) ;
    buf_clk cell_6494 ( .C ( clk ), .D ( signal_21186 ), .Q ( signal_21187 ) ) ;
    buf_clk cell_6502 ( .C ( clk ), .D ( signal_21194 ), .Q ( signal_21195 ) ) ;
    buf_clk cell_6510 ( .C ( clk ), .D ( signal_21202 ), .Q ( signal_21203 ) ) ;
    buf_clk cell_6518 ( .C ( clk ), .D ( signal_21210 ), .Q ( signal_21211 ) ) ;
    buf_clk cell_6526 ( .C ( clk ), .D ( signal_21218 ), .Q ( signal_21219 ) ) ;
    buf_clk cell_6534 ( .C ( clk ), .D ( signal_21226 ), .Q ( signal_21227 ) ) ;
    buf_clk cell_6540 ( .C ( clk ), .D ( signal_21232 ), .Q ( signal_21233 ) ) ;
    buf_clk cell_6546 ( .C ( clk ), .D ( signal_21238 ), .Q ( signal_21239 ) ) ;
    buf_clk cell_6552 ( .C ( clk ), .D ( signal_21244 ), .Q ( signal_21245 ) ) ;
    buf_clk cell_6558 ( .C ( clk ), .D ( signal_21250 ), .Q ( signal_21251 ) ) ;
    buf_clk cell_6564 ( .C ( clk ), .D ( signal_21256 ), .Q ( signal_21257 ) ) ;
    buf_clk cell_6570 ( .C ( clk ), .D ( signal_21262 ), .Q ( signal_21263 ) ) ;
    buf_clk cell_6576 ( .C ( clk ), .D ( signal_21268 ), .Q ( signal_21269 ) ) ;
    buf_clk cell_6582 ( .C ( clk ), .D ( signal_21274 ), .Q ( signal_21275 ) ) ;
    buf_clk cell_6588 ( .C ( clk ), .D ( signal_21280 ), .Q ( signal_21281 ) ) ;
    buf_clk cell_6594 ( .C ( clk ), .D ( signal_21286 ), .Q ( signal_21287 ) ) ;
    buf_clk cell_6596 ( .C ( clk ), .D ( signal_21288 ), .Q ( signal_21289 ) ) ;
    buf_clk cell_6598 ( .C ( clk ), .D ( signal_21290 ), .Q ( signal_21291 ) ) ;
    buf_clk cell_6600 ( .C ( clk ), .D ( signal_21292 ), .Q ( signal_21293 ) ) ;
    buf_clk cell_6602 ( .C ( clk ), .D ( signal_21294 ), .Q ( signal_21295 ) ) ;
    buf_clk cell_6604 ( .C ( clk ), .D ( signal_21296 ), .Q ( signal_21297 ) ) ;
    buf_clk cell_6606 ( .C ( clk ), .D ( signal_21298 ), .Q ( signal_21299 ) ) ;
    buf_clk cell_6608 ( .C ( clk ), .D ( signal_21300 ), .Q ( signal_21301 ) ) ;
    buf_clk cell_6610 ( .C ( clk ), .D ( signal_21302 ), .Q ( signal_21303 ) ) ;
    buf_clk cell_6612 ( .C ( clk ), .D ( signal_21304 ), .Q ( signal_21305 ) ) ;
    buf_clk cell_6614 ( .C ( clk ), .D ( signal_21306 ), .Q ( signal_21307 ) ) ;
    buf_clk cell_6620 ( .C ( clk ), .D ( signal_21312 ), .Q ( signal_21313 ) ) ;
    buf_clk cell_6626 ( .C ( clk ), .D ( signal_21318 ), .Q ( signal_21319 ) ) ;
    buf_clk cell_6632 ( .C ( clk ), .D ( signal_21324 ), .Q ( signal_21325 ) ) ;
    buf_clk cell_6638 ( .C ( clk ), .D ( signal_21330 ), .Q ( signal_21331 ) ) ;
    buf_clk cell_6644 ( .C ( clk ), .D ( signal_21336 ), .Q ( signal_21337 ) ) ;
    buf_clk cell_6646 ( .C ( clk ), .D ( signal_21338 ), .Q ( signal_21339 ) ) ;
    buf_clk cell_6648 ( .C ( clk ), .D ( signal_21340 ), .Q ( signal_21341 ) ) ;
    buf_clk cell_6650 ( .C ( clk ), .D ( signal_21342 ), .Q ( signal_21343 ) ) ;
    buf_clk cell_6652 ( .C ( clk ), .D ( signal_21344 ), .Q ( signal_21345 ) ) ;
    buf_clk cell_6654 ( .C ( clk ), .D ( signal_21346 ), .Q ( signal_21347 ) ) ;
    buf_clk cell_6656 ( .C ( clk ), .D ( signal_21348 ), .Q ( signal_21349 ) ) ;
    buf_clk cell_6658 ( .C ( clk ), .D ( signal_21350 ), .Q ( signal_21351 ) ) ;
    buf_clk cell_6660 ( .C ( clk ), .D ( signal_21352 ), .Q ( signal_21353 ) ) ;
    buf_clk cell_6662 ( .C ( clk ), .D ( signal_21354 ), .Q ( signal_21355 ) ) ;
    buf_clk cell_6664 ( .C ( clk ), .D ( signal_21356 ), .Q ( signal_21357 ) ) ;
    buf_clk cell_6670 ( .C ( clk ), .D ( signal_21362 ), .Q ( signal_21363 ) ) ;
    buf_clk cell_6676 ( .C ( clk ), .D ( signal_21368 ), .Q ( signal_21369 ) ) ;
    buf_clk cell_6682 ( .C ( clk ), .D ( signal_21374 ), .Q ( signal_21375 ) ) ;
    buf_clk cell_6688 ( .C ( clk ), .D ( signal_21380 ), .Q ( signal_21381 ) ) ;
    buf_clk cell_6694 ( .C ( clk ), .D ( signal_21386 ), .Q ( signal_21387 ) ) ;
    buf_clk cell_6700 ( .C ( clk ), .D ( signal_21392 ), .Q ( signal_21393 ) ) ;
    buf_clk cell_6706 ( .C ( clk ), .D ( signal_21398 ), .Q ( signal_21399 ) ) ;
    buf_clk cell_6712 ( .C ( clk ), .D ( signal_21404 ), .Q ( signal_21405 ) ) ;
    buf_clk cell_6718 ( .C ( clk ), .D ( signal_21410 ), .Q ( signal_21411 ) ) ;
    buf_clk cell_6724 ( .C ( clk ), .D ( signal_21416 ), .Q ( signal_21417 ) ) ;
    buf_clk cell_6728 ( .C ( clk ), .D ( signal_21420 ), .Q ( signal_21421 ) ) ;
    buf_clk cell_6732 ( .C ( clk ), .D ( signal_21424 ), .Q ( signal_21425 ) ) ;
    buf_clk cell_6736 ( .C ( clk ), .D ( signal_21428 ), .Q ( signal_21429 ) ) ;
    buf_clk cell_6740 ( .C ( clk ), .D ( signal_21432 ), .Q ( signal_21433 ) ) ;
    buf_clk cell_6744 ( .C ( clk ), .D ( signal_21436 ), .Q ( signal_21437 ) ) ;
    buf_clk cell_6752 ( .C ( clk ), .D ( signal_21444 ), .Q ( signal_21445 ) ) ;
    buf_clk cell_6762 ( .C ( clk ), .D ( signal_21454 ), .Q ( signal_21455 ) ) ;
    buf_clk cell_6772 ( .C ( clk ), .D ( signal_21464 ), .Q ( signal_21465 ) ) ;
    buf_clk cell_6782 ( .C ( clk ), .D ( signal_21474 ), .Q ( signal_21475 ) ) ;
    buf_clk cell_6792 ( .C ( clk ), .D ( signal_21484 ), .Q ( signal_21485 ) ) ;
    buf_clk cell_6798 ( .C ( clk ), .D ( signal_21490 ), .Q ( signal_21491 ) ) ;
    buf_clk cell_6804 ( .C ( clk ), .D ( signal_21496 ), .Q ( signal_21497 ) ) ;
    buf_clk cell_6810 ( .C ( clk ), .D ( signal_21502 ), .Q ( signal_21503 ) ) ;
    buf_clk cell_6816 ( .C ( clk ), .D ( signal_21508 ), .Q ( signal_21509 ) ) ;
    buf_clk cell_6822 ( .C ( clk ), .D ( signal_21514 ), .Q ( signal_21515 ) ) ;
    buf_clk cell_6830 ( .C ( clk ), .D ( signal_21522 ), .Q ( signal_21523 ) ) ;
    buf_clk cell_6838 ( .C ( clk ), .D ( signal_21530 ), .Q ( signal_21531 ) ) ;
    buf_clk cell_6846 ( .C ( clk ), .D ( signal_21538 ), .Q ( signal_21539 ) ) ;
    buf_clk cell_6854 ( .C ( clk ), .D ( signal_21546 ), .Q ( signal_21547 ) ) ;
    buf_clk cell_6862 ( .C ( clk ), .D ( signal_21554 ), .Q ( signal_21555 ) ) ;
    buf_clk cell_6870 ( .C ( clk ), .D ( signal_21562 ), .Q ( signal_21563 ) ) ;
    buf_clk cell_6878 ( .C ( clk ), .D ( signal_21570 ), .Q ( signal_21571 ) ) ;
    buf_clk cell_6886 ( .C ( clk ), .D ( signal_21578 ), .Q ( signal_21579 ) ) ;
    buf_clk cell_6894 ( .C ( clk ), .D ( signal_21586 ), .Q ( signal_21587 ) ) ;
    buf_clk cell_6902 ( .C ( clk ), .D ( signal_21594 ), .Q ( signal_21595 ) ) ;
    buf_clk cell_6906 ( .C ( clk ), .D ( signal_21598 ), .Q ( signal_21599 ) ) ;
    buf_clk cell_6910 ( .C ( clk ), .D ( signal_21602 ), .Q ( signal_21603 ) ) ;
    buf_clk cell_6914 ( .C ( clk ), .D ( signal_21606 ), .Q ( signal_21607 ) ) ;
    buf_clk cell_6918 ( .C ( clk ), .D ( signal_21610 ), .Q ( signal_21611 ) ) ;
    buf_clk cell_6922 ( .C ( clk ), .D ( signal_21614 ), .Q ( signal_21615 ) ) ;
    buf_clk cell_6926 ( .C ( clk ), .D ( signal_21618 ), .Q ( signal_21619 ) ) ;
    buf_clk cell_6930 ( .C ( clk ), .D ( signal_21622 ), .Q ( signal_21623 ) ) ;
    buf_clk cell_6934 ( .C ( clk ), .D ( signal_21626 ), .Q ( signal_21627 ) ) ;
    buf_clk cell_6938 ( .C ( clk ), .D ( signal_21630 ), .Q ( signal_21631 ) ) ;
    buf_clk cell_6942 ( .C ( clk ), .D ( signal_21634 ), .Q ( signal_21635 ) ) ;
    buf_clk cell_6966 ( .C ( clk ), .D ( signal_21658 ), .Q ( signal_21659 ) ) ;
    buf_clk cell_6970 ( .C ( clk ), .D ( signal_21662 ), .Q ( signal_21663 ) ) ;
    buf_clk cell_6974 ( .C ( clk ), .D ( signal_21666 ), .Q ( signal_21667 ) ) ;
    buf_clk cell_6978 ( .C ( clk ), .D ( signal_21670 ), .Q ( signal_21671 ) ) ;
    buf_clk cell_6982 ( .C ( clk ), .D ( signal_21674 ), .Q ( signal_21675 ) ) ;
    buf_clk cell_6992 ( .C ( clk ), .D ( signal_21684 ), .Q ( signal_21685 ) ) ;
    buf_clk cell_7002 ( .C ( clk ), .D ( signal_21694 ), .Q ( signal_21695 ) ) ;
    buf_clk cell_7012 ( .C ( clk ), .D ( signal_21704 ), .Q ( signal_21705 ) ) ;
    buf_clk cell_7022 ( .C ( clk ), .D ( signal_21714 ), .Q ( signal_21715 ) ) ;
    buf_clk cell_7032 ( .C ( clk ), .D ( signal_21724 ), .Q ( signal_21725 ) ) ;
    buf_clk cell_7038 ( .C ( clk ), .D ( signal_21730 ), .Q ( signal_21731 ) ) ;
    buf_clk cell_7044 ( .C ( clk ), .D ( signal_21736 ), .Q ( signal_21737 ) ) ;
    buf_clk cell_7050 ( .C ( clk ), .D ( signal_21742 ), .Q ( signal_21743 ) ) ;
    buf_clk cell_7056 ( .C ( clk ), .D ( signal_21748 ), .Q ( signal_21749 ) ) ;
    buf_clk cell_7062 ( .C ( clk ), .D ( signal_21754 ), .Q ( signal_21755 ) ) ;
    buf_clk cell_7080 ( .C ( clk ), .D ( signal_21772 ), .Q ( signal_21773 ) ) ;
    buf_clk cell_7088 ( .C ( clk ), .D ( signal_21780 ), .Q ( signal_21781 ) ) ;
    buf_clk cell_7096 ( .C ( clk ), .D ( signal_21788 ), .Q ( signal_21789 ) ) ;
    buf_clk cell_7104 ( .C ( clk ), .D ( signal_21796 ), .Q ( signal_21797 ) ) ;
    buf_clk cell_7112 ( .C ( clk ), .D ( signal_21804 ), .Q ( signal_21805 ) ) ;
    buf_clk cell_7118 ( .C ( clk ), .D ( signal_21810 ), .Q ( signal_21811 ) ) ;
    buf_clk cell_7124 ( .C ( clk ), .D ( signal_21816 ), .Q ( signal_21817 ) ) ;
    buf_clk cell_7130 ( .C ( clk ), .D ( signal_21822 ), .Q ( signal_21823 ) ) ;
    buf_clk cell_7136 ( .C ( clk ), .D ( signal_21828 ), .Q ( signal_21829 ) ) ;
    buf_clk cell_7142 ( .C ( clk ), .D ( signal_21834 ), .Q ( signal_21835 ) ) ;
    buf_clk cell_7150 ( .C ( clk ), .D ( signal_21842 ), .Q ( signal_21843 ) ) ;
    buf_clk cell_7158 ( .C ( clk ), .D ( signal_21850 ), .Q ( signal_21851 ) ) ;
    buf_clk cell_7166 ( .C ( clk ), .D ( signal_21858 ), .Q ( signal_21859 ) ) ;
    buf_clk cell_7174 ( .C ( clk ), .D ( signal_21866 ), .Q ( signal_21867 ) ) ;
    buf_clk cell_7182 ( .C ( clk ), .D ( signal_21874 ), .Q ( signal_21875 ) ) ;
    buf_clk cell_7190 ( .C ( clk ), .D ( signal_21882 ), .Q ( signal_21883 ) ) ;
    buf_clk cell_7198 ( .C ( clk ), .D ( signal_21890 ), .Q ( signal_21891 ) ) ;
    buf_clk cell_7206 ( .C ( clk ), .D ( signal_21898 ), .Q ( signal_21899 ) ) ;
    buf_clk cell_7214 ( .C ( clk ), .D ( signal_21906 ), .Q ( signal_21907 ) ) ;
    buf_clk cell_7222 ( .C ( clk ), .D ( signal_21914 ), .Q ( signal_21915 ) ) ;
    buf_clk cell_7230 ( .C ( clk ), .D ( signal_21922 ), .Q ( signal_21923 ) ) ;
    buf_clk cell_7238 ( .C ( clk ), .D ( signal_21930 ), .Q ( signal_21931 ) ) ;
    buf_clk cell_7246 ( .C ( clk ), .D ( signal_21938 ), .Q ( signal_21939 ) ) ;
    buf_clk cell_7254 ( .C ( clk ), .D ( signal_21946 ), .Q ( signal_21947 ) ) ;
    buf_clk cell_7262 ( .C ( clk ), .D ( signal_21954 ), .Q ( signal_21955 ) ) ;
    buf_clk cell_7272 ( .C ( clk ), .D ( signal_21964 ), .Q ( signal_21965 ) ) ;
    buf_clk cell_7282 ( .C ( clk ), .D ( signal_21974 ), .Q ( signal_21975 ) ) ;
    buf_clk cell_7292 ( .C ( clk ), .D ( signal_21984 ), .Q ( signal_21985 ) ) ;
    buf_clk cell_7302 ( .C ( clk ), .D ( signal_21994 ), .Q ( signal_21995 ) ) ;
    buf_clk cell_7312 ( .C ( clk ), .D ( signal_22004 ), .Q ( signal_22005 ) ) ;
    buf_clk cell_7320 ( .C ( clk ), .D ( signal_22012 ), .Q ( signal_22013 ) ) ;
    buf_clk cell_7328 ( .C ( clk ), .D ( signal_22020 ), .Q ( signal_22021 ) ) ;
    buf_clk cell_7336 ( .C ( clk ), .D ( signal_22028 ), .Q ( signal_22029 ) ) ;
    buf_clk cell_7344 ( .C ( clk ), .D ( signal_22036 ), .Q ( signal_22037 ) ) ;
    buf_clk cell_7352 ( .C ( clk ), .D ( signal_22044 ), .Q ( signal_22045 ) ) ;
    buf_clk cell_7360 ( .C ( clk ), .D ( signal_22052 ), .Q ( signal_22053 ) ) ;
    buf_clk cell_7368 ( .C ( clk ), .D ( signal_22060 ), .Q ( signal_22061 ) ) ;
    buf_clk cell_7376 ( .C ( clk ), .D ( signal_22068 ), .Q ( signal_22069 ) ) ;
    buf_clk cell_7384 ( .C ( clk ), .D ( signal_22076 ), .Q ( signal_22077 ) ) ;
    buf_clk cell_7392 ( .C ( clk ), .D ( signal_22084 ), .Q ( signal_22085 ) ) ;
    buf_clk cell_7410 ( .C ( clk ), .D ( signal_22102 ), .Q ( signal_22103 ) ) ;
    buf_clk cell_7418 ( .C ( clk ), .D ( signal_22110 ), .Q ( signal_22111 ) ) ;
    buf_clk cell_7426 ( .C ( clk ), .D ( signal_22118 ), .Q ( signal_22119 ) ) ;
    buf_clk cell_7434 ( .C ( clk ), .D ( signal_22126 ), .Q ( signal_22127 ) ) ;
    buf_clk cell_7442 ( .C ( clk ), .D ( signal_22134 ), .Q ( signal_22135 ) ) ;
    buf_clk cell_7450 ( .C ( clk ), .D ( signal_22142 ), .Q ( signal_22143 ) ) ;
    buf_clk cell_7458 ( .C ( clk ), .D ( signal_22150 ), .Q ( signal_22151 ) ) ;
    buf_clk cell_7466 ( .C ( clk ), .D ( signal_22158 ), .Q ( signal_22159 ) ) ;
    buf_clk cell_7474 ( .C ( clk ), .D ( signal_22166 ), .Q ( signal_22167 ) ) ;
    buf_clk cell_7482 ( .C ( clk ), .D ( signal_22174 ), .Q ( signal_22175 ) ) ;
    buf_clk cell_7490 ( .C ( clk ), .D ( signal_22182 ), .Q ( signal_22183 ) ) ;
    buf_clk cell_7498 ( .C ( clk ), .D ( signal_22190 ), .Q ( signal_22191 ) ) ;
    buf_clk cell_7506 ( .C ( clk ), .D ( signal_22198 ), .Q ( signal_22199 ) ) ;
    buf_clk cell_7514 ( .C ( clk ), .D ( signal_22206 ), .Q ( signal_22207 ) ) ;
    buf_clk cell_7522 ( .C ( clk ), .D ( signal_22214 ), .Q ( signal_22215 ) ) ;
    buf_clk cell_7526 ( .C ( clk ), .D ( signal_22218 ), .Q ( signal_22219 ) ) ;
    buf_clk cell_7532 ( .C ( clk ), .D ( signal_22224 ), .Q ( signal_22225 ) ) ;
    buf_clk cell_7538 ( .C ( clk ), .D ( signal_22230 ), .Q ( signal_22231 ) ) ;
    buf_clk cell_7544 ( .C ( clk ), .D ( signal_22236 ), .Q ( signal_22237 ) ) ;
    buf_clk cell_7550 ( .C ( clk ), .D ( signal_22242 ), .Q ( signal_22243 ) ) ;
    buf_clk cell_7558 ( .C ( clk ), .D ( signal_22250 ), .Q ( signal_22251 ) ) ;
    buf_clk cell_7566 ( .C ( clk ), .D ( signal_22258 ), .Q ( signal_22259 ) ) ;
    buf_clk cell_7574 ( .C ( clk ), .D ( signal_22266 ), .Q ( signal_22267 ) ) ;
    buf_clk cell_7582 ( .C ( clk ), .D ( signal_22274 ), .Q ( signal_22275 ) ) ;
    buf_clk cell_7590 ( .C ( clk ), .D ( signal_22282 ), .Q ( signal_22283 ) ) ;
    buf_clk cell_7596 ( .C ( clk ), .D ( signal_22288 ), .Q ( signal_22289 ) ) ;
    buf_clk cell_7602 ( .C ( clk ), .D ( signal_22294 ), .Q ( signal_22295 ) ) ;
    buf_clk cell_7608 ( .C ( clk ), .D ( signal_22300 ), .Q ( signal_22301 ) ) ;
    buf_clk cell_7614 ( .C ( clk ), .D ( signal_22306 ), .Q ( signal_22307 ) ) ;
    buf_clk cell_7620 ( .C ( clk ), .D ( signal_22312 ), .Q ( signal_22313 ) ) ;
    buf_clk cell_7626 ( .C ( clk ), .D ( signal_22318 ), .Q ( signal_22319 ) ) ;
    buf_clk cell_7632 ( .C ( clk ), .D ( signal_22324 ), .Q ( signal_22325 ) ) ;
    buf_clk cell_7638 ( .C ( clk ), .D ( signal_22330 ), .Q ( signal_22331 ) ) ;
    buf_clk cell_7644 ( .C ( clk ), .D ( signal_22336 ), .Q ( signal_22337 ) ) ;
    buf_clk cell_7650 ( .C ( clk ), .D ( signal_22342 ), .Q ( signal_22343 ) ) ;
    buf_clk cell_7658 ( .C ( clk ), .D ( signal_22350 ), .Q ( signal_22351 ) ) ;
    buf_clk cell_7666 ( .C ( clk ), .D ( signal_22358 ), .Q ( signal_22359 ) ) ;
    buf_clk cell_7674 ( .C ( clk ), .D ( signal_22366 ), .Q ( signal_22367 ) ) ;
    buf_clk cell_7682 ( .C ( clk ), .D ( signal_22374 ), .Q ( signal_22375 ) ) ;
    buf_clk cell_7690 ( .C ( clk ), .D ( signal_22382 ), .Q ( signal_22383 ) ) ;
    buf_clk cell_7700 ( .C ( clk ), .D ( signal_22392 ), .Q ( signal_22393 ) ) ;
    buf_clk cell_7710 ( .C ( clk ), .D ( signal_22402 ), .Q ( signal_22403 ) ) ;
    buf_clk cell_7720 ( .C ( clk ), .D ( signal_22412 ), .Q ( signal_22413 ) ) ;
    buf_clk cell_7730 ( .C ( clk ), .D ( signal_22422 ), .Q ( signal_22423 ) ) ;
    buf_clk cell_7740 ( .C ( clk ), .D ( signal_22432 ), .Q ( signal_22433 ) ) ;
    buf_clk cell_7756 ( .C ( clk ), .D ( signal_22448 ), .Q ( signal_22449 ) ) ;
    buf_clk cell_7762 ( .C ( clk ), .D ( signal_22454 ), .Q ( signal_22455 ) ) ;
    buf_clk cell_7768 ( .C ( clk ), .D ( signal_22460 ), .Q ( signal_22461 ) ) ;
    buf_clk cell_7774 ( .C ( clk ), .D ( signal_22466 ), .Q ( signal_22467 ) ) ;
    buf_clk cell_7780 ( .C ( clk ), .D ( signal_22472 ), .Q ( signal_22473 ) ) ;
    buf_clk cell_7788 ( .C ( clk ), .D ( signal_22480 ), .Q ( signal_22481 ) ) ;
    buf_clk cell_7796 ( .C ( clk ), .D ( signal_22488 ), .Q ( signal_22489 ) ) ;
    buf_clk cell_7804 ( .C ( clk ), .D ( signal_22496 ), .Q ( signal_22497 ) ) ;
    buf_clk cell_7812 ( .C ( clk ), .D ( signal_22504 ), .Q ( signal_22505 ) ) ;
    buf_clk cell_7820 ( .C ( clk ), .D ( signal_22512 ), .Q ( signal_22513 ) ) ;
    buf_clk cell_7830 ( .C ( clk ), .D ( signal_22522 ), .Q ( signal_22523 ) ) ;
    buf_clk cell_7840 ( .C ( clk ), .D ( signal_22532 ), .Q ( signal_22533 ) ) ;
    buf_clk cell_7850 ( .C ( clk ), .D ( signal_22542 ), .Q ( signal_22543 ) ) ;
    buf_clk cell_7860 ( .C ( clk ), .D ( signal_22552 ), .Q ( signal_22553 ) ) ;
    buf_clk cell_7870 ( .C ( clk ), .D ( signal_22562 ), .Q ( signal_22563 ) ) ;
    buf_clk cell_7878 ( .C ( clk ), .D ( signal_22570 ), .Q ( signal_22571 ) ) ;
    buf_clk cell_7886 ( .C ( clk ), .D ( signal_22578 ), .Q ( signal_22579 ) ) ;
    buf_clk cell_7894 ( .C ( clk ), .D ( signal_22586 ), .Q ( signal_22587 ) ) ;
    buf_clk cell_7902 ( .C ( clk ), .D ( signal_22594 ), .Q ( signal_22595 ) ) ;
    buf_clk cell_7910 ( .C ( clk ), .D ( signal_22602 ), .Q ( signal_22603 ) ) ;
    buf_clk cell_7916 ( .C ( clk ), .D ( signal_22608 ), .Q ( signal_22609 ) ) ;
    buf_clk cell_7922 ( .C ( clk ), .D ( signal_22614 ), .Q ( signal_22615 ) ) ;
    buf_clk cell_7928 ( .C ( clk ), .D ( signal_22620 ), .Q ( signal_22621 ) ) ;
    buf_clk cell_7934 ( .C ( clk ), .D ( signal_22626 ), .Q ( signal_22627 ) ) ;
    buf_clk cell_7940 ( .C ( clk ), .D ( signal_22632 ), .Q ( signal_22633 ) ) ;
    buf_clk cell_7946 ( .C ( clk ), .D ( signal_22638 ), .Q ( signal_22639 ) ) ;
    buf_clk cell_7952 ( .C ( clk ), .D ( signal_22644 ), .Q ( signal_22645 ) ) ;
    buf_clk cell_7958 ( .C ( clk ), .D ( signal_22650 ), .Q ( signal_22651 ) ) ;
    buf_clk cell_7964 ( .C ( clk ), .D ( signal_22656 ), .Q ( signal_22657 ) ) ;
    buf_clk cell_7970 ( .C ( clk ), .D ( signal_22662 ), .Q ( signal_22663 ) ) ;
    buf_clk cell_8026 ( .C ( clk ), .D ( signal_22718 ), .Q ( signal_22719 ) ) ;
    buf_clk cell_8032 ( .C ( clk ), .D ( signal_22724 ), .Q ( signal_22725 ) ) ;
    buf_clk cell_8038 ( .C ( clk ), .D ( signal_22730 ), .Q ( signal_22731 ) ) ;
    buf_clk cell_8044 ( .C ( clk ), .D ( signal_22736 ), .Q ( signal_22737 ) ) ;
    buf_clk cell_8050 ( .C ( clk ), .D ( signal_22742 ), .Q ( signal_22743 ) ) ;
    buf_clk cell_8066 ( .C ( clk ), .D ( signal_22758 ), .Q ( signal_22759 ) ) ;
    buf_clk cell_8072 ( .C ( clk ), .D ( signal_22764 ), .Q ( signal_22765 ) ) ;
    buf_clk cell_8078 ( .C ( clk ), .D ( signal_22770 ), .Q ( signal_22771 ) ) ;
    buf_clk cell_8084 ( .C ( clk ), .D ( signal_22776 ), .Q ( signal_22777 ) ) ;
    buf_clk cell_8090 ( .C ( clk ), .D ( signal_22782 ), .Q ( signal_22783 ) ) ;
    buf_clk cell_8116 ( .C ( clk ), .D ( signal_22808 ), .Q ( signal_22809 ) ) ;
    buf_clk cell_8122 ( .C ( clk ), .D ( signal_22814 ), .Q ( signal_22815 ) ) ;
    buf_clk cell_8128 ( .C ( clk ), .D ( signal_22820 ), .Q ( signal_22821 ) ) ;
    buf_clk cell_8134 ( .C ( clk ), .D ( signal_22826 ), .Q ( signal_22827 ) ) ;
    buf_clk cell_8140 ( .C ( clk ), .D ( signal_22832 ), .Q ( signal_22833 ) ) ;
    buf_clk cell_8206 ( .C ( clk ), .D ( signal_22898 ), .Q ( signal_22899 ) ) ;
    buf_clk cell_8214 ( .C ( clk ), .D ( signal_22906 ), .Q ( signal_22907 ) ) ;
    buf_clk cell_8222 ( .C ( clk ), .D ( signal_22914 ), .Q ( signal_22915 ) ) ;
    buf_clk cell_8230 ( .C ( clk ), .D ( signal_22922 ), .Q ( signal_22923 ) ) ;
    buf_clk cell_8238 ( .C ( clk ), .D ( signal_22930 ), .Q ( signal_22931 ) ) ;
    buf_clk cell_8278 ( .C ( clk ), .D ( signal_22970 ), .Q ( signal_22971 ) ) ;
    buf_clk cell_8288 ( .C ( clk ), .D ( signal_22980 ), .Q ( signal_22981 ) ) ;
    buf_clk cell_8298 ( .C ( clk ), .D ( signal_22990 ), .Q ( signal_22991 ) ) ;
    buf_clk cell_8308 ( .C ( clk ), .D ( signal_23000 ), .Q ( signal_23001 ) ) ;
    buf_clk cell_8318 ( .C ( clk ), .D ( signal_23010 ), .Q ( signal_23011 ) ) ;
    buf_clk cell_8376 ( .C ( clk ), .D ( signal_23068 ), .Q ( signal_23069 ) ) ;
    buf_clk cell_8384 ( .C ( clk ), .D ( signal_23076 ), .Q ( signal_23077 ) ) ;
    buf_clk cell_8392 ( .C ( clk ), .D ( signal_23084 ), .Q ( signal_23085 ) ) ;
    buf_clk cell_8400 ( .C ( clk ), .D ( signal_23092 ), .Q ( signal_23093 ) ) ;
    buf_clk cell_8408 ( .C ( clk ), .D ( signal_23100 ), .Q ( signal_23101 ) ) ;
    buf_clk cell_8446 ( .C ( clk ), .D ( signal_23138 ), .Q ( signal_23139 ) ) ;
    buf_clk cell_8454 ( .C ( clk ), .D ( signal_23146 ), .Q ( signal_23147 ) ) ;
    buf_clk cell_8462 ( .C ( clk ), .D ( signal_23154 ), .Q ( signal_23155 ) ) ;
    buf_clk cell_8470 ( .C ( clk ), .D ( signal_23162 ), .Q ( signal_23163 ) ) ;
    buf_clk cell_8478 ( .C ( clk ), .D ( signal_23170 ), .Q ( signal_23171 ) ) ;
    buf_clk cell_8516 ( .C ( clk ), .D ( signal_23208 ), .Q ( signal_23209 ) ) ;
    buf_clk cell_8524 ( .C ( clk ), .D ( signal_23216 ), .Q ( signal_23217 ) ) ;
    buf_clk cell_8532 ( .C ( clk ), .D ( signal_23224 ), .Q ( signal_23225 ) ) ;
    buf_clk cell_8540 ( .C ( clk ), .D ( signal_23232 ), .Q ( signal_23233 ) ) ;
    buf_clk cell_8548 ( .C ( clk ), .D ( signal_23240 ), .Q ( signal_23241 ) ) ;
    buf_clk cell_8718 ( .C ( clk ), .D ( signal_23410 ), .Q ( signal_23411 ) ) ;
    buf_clk cell_8730 ( .C ( clk ), .D ( signal_23422 ), .Q ( signal_23423 ) ) ;
    buf_clk cell_8742 ( .C ( clk ), .D ( signal_23434 ), .Q ( signal_23435 ) ) ;
    buf_clk cell_8754 ( .C ( clk ), .D ( signal_23446 ), .Q ( signal_23447 ) ) ;
    buf_clk cell_8766 ( .C ( clk ), .D ( signal_23458 ), .Q ( signal_23459 ) ) ;
    buf_clk cell_8840 ( .C ( clk ), .D ( signal_23532 ), .Q ( signal_23533 ) ) ;
    buf_clk cell_8854 ( .C ( clk ), .D ( signal_23546 ), .Q ( signal_23547 ) ) ;
    buf_clk cell_8868 ( .C ( clk ), .D ( signal_23560 ), .Q ( signal_23561 ) ) ;
    buf_clk cell_8882 ( .C ( clk ), .D ( signal_23574 ), .Q ( signal_23575 ) ) ;
    buf_clk cell_8896 ( .C ( clk ), .D ( signal_23588 ), .Q ( signal_23589 ) ) ;
    buf_clk cell_8950 ( .C ( clk ), .D ( signal_23642 ), .Q ( signal_23643 ) ) ;
    buf_clk cell_8964 ( .C ( clk ), .D ( signal_23656 ), .Q ( signal_23657 ) ) ;
    buf_clk cell_8978 ( .C ( clk ), .D ( signal_23670 ), .Q ( signal_23671 ) ) ;
    buf_clk cell_8992 ( .C ( clk ), .D ( signal_23684 ), .Q ( signal_23685 ) ) ;
    buf_clk cell_9006 ( .C ( clk ), .D ( signal_23698 ), .Q ( signal_23699 ) ) ;
    buf_clk cell_9150 ( .C ( clk ), .D ( signal_23842 ), .Q ( signal_23843 ) ) ;
    buf_clk cell_9166 ( .C ( clk ), .D ( signal_23858 ), .Q ( signal_23859 ) ) ;
    buf_clk cell_9182 ( .C ( clk ), .D ( signal_23874 ), .Q ( signal_23875 ) ) ;
    buf_clk cell_9198 ( .C ( clk ), .D ( signal_23890 ), .Q ( signal_23891 ) ) ;
    buf_clk cell_9214 ( .C ( clk ), .D ( signal_23906 ), .Q ( signal_23907 ) ) ;
    buf_clk cell_9250 ( .C ( clk ), .D ( signal_23942 ), .Q ( signal_23943 ) ) ;
    buf_clk cell_9266 ( .C ( clk ), .D ( signal_23958 ), .Q ( signal_23959 ) ) ;
    buf_clk cell_9282 ( .C ( clk ), .D ( signal_23974 ), .Q ( signal_23975 ) ) ;
    buf_clk cell_9298 ( .C ( clk ), .D ( signal_23990 ), .Q ( signal_23991 ) ) ;
    buf_clk cell_9314 ( .C ( clk ), .D ( signal_24006 ), .Q ( signal_24007 ) ) ;
    buf_clk cell_9558 ( .C ( clk ), .D ( signal_24250 ), .Q ( signal_24251 ) ) ;
    buf_clk cell_9574 ( .C ( clk ), .D ( signal_24266 ), .Q ( signal_24267 ) ) ;
    buf_clk cell_9590 ( .C ( clk ), .D ( signal_24282 ), .Q ( signal_24283 ) ) ;
    buf_clk cell_9606 ( .C ( clk ), .D ( signal_24298 ), .Q ( signal_24299 ) ) ;
    buf_clk cell_9622 ( .C ( clk ), .D ( signal_24314 ), .Q ( signal_24315 ) ) ;
    buf_clk cell_9640 ( .C ( clk ), .D ( signal_24332 ), .Q ( signal_24333 ) ) ;
    buf_clk cell_9658 ( .C ( clk ), .D ( signal_24350 ), .Q ( signal_24351 ) ) ;
    buf_clk cell_9676 ( .C ( clk ), .D ( signal_24368 ), .Q ( signal_24369 ) ) ;
    buf_clk cell_9694 ( .C ( clk ), .D ( signal_24386 ), .Q ( signal_24387 ) ) ;
    buf_clk cell_9712 ( .C ( clk ), .D ( signal_24404 ), .Q ( signal_24405 ) ) ;
    buf_clk cell_9890 ( .C ( clk ), .D ( signal_24582 ), .Q ( signal_24583 ) ) ;
    buf_clk cell_9910 ( .C ( clk ), .D ( signal_24602 ), .Q ( signal_24603 ) ) ;
    buf_clk cell_9930 ( .C ( clk ), .D ( signal_24622 ), .Q ( signal_24623 ) ) ;
    buf_clk cell_9950 ( .C ( clk ), .D ( signal_24642 ), .Q ( signal_24643 ) ) ;
    buf_clk cell_9970 ( .C ( clk ), .D ( signal_24662 ), .Q ( signal_24663 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_6753 ( .C ( clk ), .D ( signal_21445 ), .Q ( signal_21446 ) ) ;
    buf_clk cell_6763 ( .C ( clk ), .D ( signal_21455 ), .Q ( signal_21456 ) ) ;
    buf_clk cell_6773 ( .C ( clk ), .D ( signal_21465 ), .Q ( signal_21466 ) ) ;
    buf_clk cell_6783 ( .C ( clk ), .D ( signal_21475 ), .Q ( signal_21476 ) ) ;
    buf_clk cell_6793 ( .C ( clk ), .D ( signal_21485 ), .Q ( signal_21486 ) ) ;
    buf_clk cell_6799 ( .C ( clk ), .D ( signal_21491 ), .Q ( signal_21492 ) ) ;
    buf_clk cell_6805 ( .C ( clk ), .D ( signal_21497 ), .Q ( signal_21498 ) ) ;
    buf_clk cell_6811 ( .C ( clk ), .D ( signal_21503 ), .Q ( signal_21504 ) ) ;
    buf_clk cell_6817 ( .C ( clk ), .D ( signal_21509 ), .Q ( signal_21510 ) ) ;
    buf_clk cell_6823 ( .C ( clk ), .D ( signal_21515 ), .Q ( signal_21516 ) ) ;
    buf_clk cell_6831 ( .C ( clk ), .D ( signal_21523 ), .Q ( signal_21524 ) ) ;
    buf_clk cell_6839 ( .C ( clk ), .D ( signal_21531 ), .Q ( signal_21532 ) ) ;
    buf_clk cell_6847 ( .C ( clk ), .D ( signal_21539 ), .Q ( signal_21540 ) ) ;
    buf_clk cell_6855 ( .C ( clk ), .D ( signal_21547 ), .Q ( signal_21548 ) ) ;
    buf_clk cell_6863 ( .C ( clk ), .D ( signal_21555 ), .Q ( signal_21556 ) ) ;
    buf_clk cell_6871 ( .C ( clk ), .D ( signal_21563 ), .Q ( signal_21564 ) ) ;
    buf_clk cell_6879 ( .C ( clk ), .D ( signal_21571 ), .Q ( signal_21572 ) ) ;
    buf_clk cell_6887 ( .C ( clk ), .D ( signal_21579 ), .Q ( signal_21580 ) ) ;
    buf_clk cell_6895 ( .C ( clk ), .D ( signal_21587 ), .Q ( signal_21588 ) ) ;
    buf_clk cell_6903 ( .C ( clk ), .D ( signal_21595 ), .Q ( signal_21596 ) ) ;
    buf_clk cell_6907 ( .C ( clk ), .D ( signal_21599 ), .Q ( signal_21600 ) ) ;
    buf_clk cell_6911 ( .C ( clk ), .D ( signal_21603 ), .Q ( signal_21604 ) ) ;
    buf_clk cell_6915 ( .C ( clk ), .D ( signal_21607 ), .Q ( signal_21608 ) ) ;
    buf_clk cell_6919 ( .C ( clk ), .D ( signal_21611 ), .Q ( signal_21612 ) ) ;
    buf_clk cell_6923 ( .C ( clk ), .D ( signal_21615 ), .Q ( signal_21616 ) ) ;
    buf_clk cell_6927 ( .C ( clk ), .D ( signal_21619 ), .Q ( signal_21620 ) ) ;
    buf_clk cell_6931 ( .C ( clk ), .D ( signal_21623 ), .Q ( signal_21624 ) ) ;
    buf_clk cell_6935 ( .C ( clk ), .D ( signal_21627 ), .Q ( signal_21628 ) ) ;
    buf_clk cell_6939 ( .C ( clk ), .D ( signal_21631 ), .Q ( signal_21632 ) ) ;
    buf_clk cell_6943 ( .C ( clk ), .D ( signal_21635 ), .Q ( signal_21636 ) ) ;
    buf_clk cell_6945 ( .C ( clk ), .D ( signal_21349 ), .Q ( signal_21638 ) ) ;
    buf_clk cell_6947 ( .C ( clk ), .D ( signal_21351 ), .Q ( signal_21640 ) ) ;
    buf_clk cell_6949 ( .C ( clk ), .D ( signal_21353 ), .Q ( signal_21642 ) ) ;
    buf_clk cell_6951 ( .C ( clk ), .D ( signal_21355 ), .Q ( signal_21644 ) ) ;
    buf_clk cell_6953 ( .C ( clk ), .D ( signal_21357 ), .Q ( signal_21646 ) ) ;
    buf_clk cell_6955 ( .C ( clk ), .D ( signal_2156 ), .Q ( signal_21648 ) ) ;
    buf_clk cell_6957 ( .C ( clk ), .D ( signal_7280 ), .Q ( signal_21650 ) ) ;
    buf_clk cell_6959 ( .C ( clk ), .D ( signal_7281 ), .Q ( signal_21652 ) ) ;
    buf_clk cell_6961 ( .C ( clk ), .D ( signal_7282 ), .Q ( signal_21654 ) ) ;
    buf_clk cell_6963 ( .C ( clk ), .D ( signal_7283 ), .Q ( signal_21656 ) ) ;
    buf_clk cell_6967 ( .C ( clk ), .D ( signal_21659 ), .Q ( signal_21660 ) ) ;
    buf_clk cell_6971 ( .C ( clk ), .D ( signal_21663 ), .Q ( signal_21664 ) ) ;
    buf_clk cell_6975 ( .C ( clk ), .D ( signal_21667 ), .Q ( signal_21668 ) ) ;
    buf_clk cell_6979 ( .C ( clk ), .D ( signal_21671 ), .Q ( signal_21672 ) ) ;
    buf_clk cell_6983 ( .C ( clk ), .D ( signal_21675 ), .Q ( signal_21676 ) ) ;
    buf_clk cell_6993 ( .C ( clk ), .D ( signal_21685 ), .Q ( signal_21686 ) ) ;
    buf_clk cell_7003 ( .C ( clk ), .D ( signal_21695 ), .Q ( signal_21696 ) ) ;
    buf_clk cell_7013 ( .C ( clk ), .D ( signal_21705 ), .Q ( signal_21706 ) ) ;
    buf_clk cell_7023 ( .C ( clk ), .D ( signal_21715 ), .Q ( signal_21716 ) ) ;
    buf_clk cell_7033 ( .C ( clk ), .D ( signal_21725 ), .Q ( signal_21726 ) ) ;
    buf_clk cell_7039 ( .C ( clk ), .D ( signal_21731 ), .Q ( signal_21732 ) ) ;
    buf_clk cell_7045 ( .C ( clk ), .D ( signal_21737 ), .Q ( signal_21738 ) ) ;
    buf_clk cell_7051 ( .C ( clk ), .D ( signal_21743 ), .Q ( signal_21744 ) ) ;
    buf_clk cell_7057 ( .C ( clk ), .D ( signal_21749 ), .Q ( signal_21750 ) ) ;
    buf_clk cell_7063 ( .C ( clk ), .D ( signal_21755 ), .Q ( signal_21756 ) ) ;
    buf_clk cell_7065 ( .C ( clk ), .D ( signal_20931 ), .Q ( signal_21758 ) ) ;
    buf_clk cell_7067 ( .C ( clk ), .D ( signal_20935 ), .Q ( signal_21760 ) ) ;
    buf_clk cell_7069 ( .C ( clk ), .D ( signal_20939 ), .Q ( signal_21762 ) ) ;
    buf_clk cell_7071 ( .C ( clk ), .D ( signal_20943 ), .Q ( signal_21764 ) ) ;
    buf_clk cell_7073 ( .C ( clk ), .D ( signal_20947 ), .Q ( signal_21766 ) ) ;
    buf_clk cell_7081 ( .C ( clk ), .D ( signal_21773 ), .Q ( signal_21774 ) ) ;
    buf_clk cell_7089 ( .C ( clk ), .D ( signal_21781 ), .Q ( signal_21782 ) ) ;
    buf_clk cell_7097 ( .C ( clk ), .D ( signal_21789 ), .Q ( signal_21790 ) ) ;
    buf_clk cell_7105 ( .C ( clk ), .D ( signal_21797 ), .Q ( signal_21798 ) ) ;
    buf_clk cell_7113 ( .C ( clk ), .D ( signal_21805 ), .Q ( signal_21806 ) ) ;
    buf_clk cell_7119 ( .C ( clk ), .D ( signal_21811 ), .Q ( signal_21812 ) ) ;
    buf_clk cell_7125 ( .C ( clk ), .D ( signal_21817 ), .Q ( signal_21818 ) ) ;
    buf_clk cell_7131 ( .C ( clk ), .D ( signal_21823 ), .Q ( signal_21824 ) ) ;
    buf_clk cell_7137 ( .C ( clk ), .D ( signal_21829 ), .Q ( signal_21830 ) ) ;
    buf_clk cell_7143 ( .C ( clk ), .D ( signal_21835 ), .Q ( signal_21836 ) ) ;
    buf_clk cell_7151 ( .C ( clk ), .D ( signal_21843 ), .Q ( signal_21844 ) ) ;
    buf_clk cell_7159 ( .C ( clk ), .D ( signal_21851 ), .Q ( signal_21852 ) ) ;
    buf_clk cell_7167 ( .C ( clk ), .D ( signal_21859 ), .Q ( signal_21860 ) ) ;
    buf_clk cell_7175 ( .C ( clk ), .D ( signal_21867 ), .Q ( signal_21868 ) ) ;
    buf_clk cell_7183 ( .C ( clk ), .D ( signal_21875 ), .Q ( signal_21876 ) ) ;
    buf_clk cell_7191 ( .C ( clk ), .D ( signal_21883 ), .Q ( signal_21884 ) ) ;
    buf_clk cell_7199 ( .C ( clk ), .D ( signal_21891 ), .Q ( signal_21892 ) ) ;
    buf_clk cell_7207 ( .C ( clk ), .D ( signal_21899 ), .Q ( signal_21900 ) ) ;
    buf_clk cell_7215 ( .C ( clk ), .D ( signal_21907 ), .Q ( signal_21908 ) ) ;
    buf_clk cell_7223 ( .C ( clk ), .D ( signal_21915 ), .Q ( signal_21916 ) ) ;
    buf_clk cell_7231 ( .C ( clk ), .D ( signal_21923 ), .Q ( signal_21924 ) ) ;
    buf_clk cell_7239 ( .C ( clk ), .D ( signal_21931 ), .Q ( signal_21932 ) ) ;
    buf_clk cell_7247 ( .C ( clk ), .D ( signal_21939 ), .Q ( signal_21940 ) ) ;
    buf_clk cell_7255 ( .C ( clk ), .D ( signal_21947 ), .Q ( signal_21948 ) ) ;
    buf_clk cell_7263 ( .C ( clk ), .D ( signal_21955 ), .Q ( signal_21956 ) ) ;
    buf_clk cell_7273 ( .C ( clk ), .D ( signal_21965 ), .Q ( signal_21966 ) ) ;
    buf_clk cell_7283 ( .C ( clk ), .D ( signal_21975 ), .Q ( signal_21976 ) ) ;
    buf_clk cell_7293 ( .C ( clk ), .D ( signal_21985 ), .Q ( signal_21986 ) ) ;
    buf_clk cell_7303 ( .C ( clk ), .D ( signal_21995 ), .Q ( signal_21996 ) ) ;
    buf_clk cell_7313 ( .C ( clk ), .D ( signal_22005 ), .Q ( signal_22006 ) ) ;
    buf_clk cell_7321 ( .C ( clk ), .D ( signal_22013 ), .Q ( signal_22014 ) ) ;
    buf_clk cell_7329 ( .C ( clk ), .D ( signal_22021 ), .Q ( signal_22022 ) ) ;
    buf_clk cell_7337 ( .C ( clk ), .D ( signal_22029 ), .Q ( signal_22030 ) ) ;
    buf_clk cell_7345 ( .C ( clk ), .D ( signal_22037 ), .Q ( signal_22038 ) ) ;
    buf_clk cell_7353 ( .C ( clk ), .D ( signal_22045 ), .Q ( signal_22046 ) ) ;
    buf_clk cell_7361 ( .C ( clk ), .D ( signal_22053 ), .Q ( signal_22054 ) ) ;
    buf_clk cell_7369 ( .C ( clk ), .D ( signal_22061 ), .Q ( signal_22062 ) ) ;
    buf_clk cell_7377 ( .C ( clk ), .D ( signal_22069 ), .Q ( signal_22070 ) ) ;
    buf_clk cell_7385 ( .C ( clk ), .D ( signal_22077 ), .Q ( signal_22078 ) ) ;
    buf_clk cell_7393 ( .C ( clk ), .D ( signal_22085 ), .Q ( signal_22086 ) ) ;
    buf_clk cell_7395 ( .C ( clk ), .D ( signal_20819 ), .Q ( signal_22088 ) ) ;
    buf_clk cell_7397 ( .C ( clk ), .D ( signal_20821 ), .Q ( signal_22090 ) ) ;
    buf_clk cell_7399 ( .C ( clk ), .D ( signal_20823 ), .Q ( signal_22092 ) ) ;
    buf_clk cell_7401 ( .C ( clk ), .D ( signal_20825 ), .Q ( signal_22094 ) ) ;
    buf_clk cell_7403 ( .C ( clk ), .D ( signal_20827 ), .Q ( signal_22096 ) ) ;
    buf_clk cell_7411 ( .C ( clk ), .D ( signal_22103 ), .Q ( signal_22104 ) ) ;
    buf_clk cell_7419 ( .C ( clk ), .D ( signal_22111 ), .Q ( signal_22112 ) ) ;
    buf_clk cell_7427 ( .C ( clk ), .D ( signal_22119 ), .Q ( signal_22120 ) ) ;
    buf_clk cell_7435 ( .C ( clk ), .D ( signal_22127 ), .Q ( signal_22128 ) ) ;
    buf_clk cell_7443 ( .C ( clk ), .D ( signal_22135 ), .Q ( signal_22136 ) ) ;
    buf_clk cell_7451 ( .C ( clk ), .D ( signal_22143 ), .Q ( signal_22144 ) ) ;
    buf_clk cell_7459 ( .C ( clk ), .D ( signal_22151 ), .Q ( signal_22152 ) ) ;
    buf_clk cell_7467 ( .C ( clk ), .D ( signal_22159 ), .Q ( signal_22160 ) ) ;
    buf_clk cell_7475 ( .C ( clk ), .D ( signal_22167 ), .Q ( signal_22168 ) ) ;
    buf_clk cell_7483 ( .C ( clk ), .D ( signal_22175 ), .Q ( signal_22176 ) ) ;
    buf_clk cell_7491 ( .C ( clk ), .D ( signal_22183 ), .Q ( signal_22184 ) ) ;
    buf_clk cell_7499 ( .C ( clk ), .D ( signal_22191 ), .Q ( signal_22192 ) ) ;
    buf_clk cell_7507 ( .C ( clk ), .D ( signal_22199 ), .Q ( signal_22200 ) ) ;
    buf_clk cell_7515 ( .C ( clk ), .D ( signal_22207 ), .Q ( signal_22208 ) ) ;
    buf_clk cell_7523 ( .C ( clk ), .D ( signal_22215 ), .Q ( signal_22216 ) ) ;
    buf_clk cell_7527 ( .C ( clk ), .D ( signal_22219 ), .Q ( signal_22220 ) ) ;
    buf_clk cell_7533 ( .C ( clk ), .D ( signal_22225 ), .Q ( signal_22226 ) ) ;
    buf_clk cell_7539 ( .C ( clk ), .D ( signal_22231 ), .Q ( signal_22232 ) ) ;
    buf_clk cell_7545 ( .C ( clk ), .D ( signal_22237 ), .Q ( signal_22238 ) ) ;
    buf_clk cell_7551 ( .C ( clk ), .D ( signal_22243 ), .Q ( signal_22244 ) ) ;
    buf_clk cell_7559 ( .C ( clk ), .D ( signal_22251 ), .Q ( signal_22252 ) ) ;
    buf_clk cell_7567 ( .C ( clk ), .D ( signal_22259 ), .Q ( signal_22260 ) ) ;
    buf_clk cell_7575 ( .C ( clk ), .D ( signal_22267 ), .Q ( signal_22268 ) ) ;
    buf_clk cell_7583 ( .C ( clk ), .D ( signal_22275 ), .Q ( signal_22276 ) ) ;
    buf_clk cell_7591 ( .C ( clk ), .D ( signal_22283 ), .Q ( signal_22284 ) ) ;
    buf_clk cell_7597 ( .C ( clk ), .D ( signal_22289 ), .Q ( signal_22290 ) ) ;
    buf_clk cell_7603 ( .C ( clk ), .D ( signal_22295 ), .Q ( signal_22296 ) ) ;
    buf_clk cell_7609 ( .C ( clk ), .D ( signal_22301 ), .Q ( signal_22302 ) ) ;
    buf_clk cell_7615 ( .C ( clk ), .D ( signal_22307 ), .Q ( signal_22308 ) ) ;
    buf_clk cell_7621 ( .C ( clk ), .D ( signal_22313 ), .Q ( signal_22314 ) ) ;
    buf_clk cell_7627 ( .C ( clk ), .D ( signal_22319 ), .Q ( signal_22320 ) ) ;
    buf_clk cell_7633 ( .C ( clk ), .D ( signal_22325 ), .Q ( signal_22326 ) ) ;
    buf_clk cell_7639 ( .C ( clk ), .D ( signal_22331 ), .Q ( signal_22332 ) ) ;
    buf_clk cell_7645 ( .C ( clk ), .D ( signal_22337 ), .Q ( signal_22338 ) ) ;
    buf_clk cell_7651 ( .C ( clk ), .D ( signal_22343 ), .Q ( signal_22344 ) ) ;
    buf_clk cell_7659 ( .C ( clk ), .D ( signal_22351 ), .Q ( signal_22352 ) ) ;
    buf_clk cell_7667 ( .C ( clk ), .D ( signal_22359 ), .Q ( signal_22360 ) ) ;
    buf_clk cell_7675 ( .C ( clk ), .D ( signal_22367 ), .Q ( signal_22368 ) ) ;
    buf_clk cell_7683 ( .C ( clk ), .D ( signal_22375 ), .Q ( signal_22376 ) ) ;
    buf_clk cell_7691 ( .C ( clk ), .D ( signal_22383 ), .Q ( signal_22384 ) ) ;
    buf_clk cell_7701 ( .C ( clk ), .D ( signal_22393 ), .Q ( signal_22394 ) ) ;
    buf_clk cell_7711 ( .C ( clk ), .D ( signal_22403 ), .Q ( signal_22404 ) ) ;
    buf_clk cell_7721 ( .C ( clk ), .D ( signal_22413 ), .Q ( signal_22414 ) ) ;
    buf_clk cell_7731 ( .C ( clk ), .D ( signal_22423 ), .Q ( signal_22424 ) ) ;
    buf_clk cell_7741 ( .C ( clk ), .D ( signal_22433 ), .Q ( signal_22434 ) ) ;
    buf_clk cell_7757 ( .C ( clk ), .D ( signal_22449 ), .Q ( signal_22450 ) ) ;
    buf_clk cell_7763 ( .C ( clk ), .D ( signal_22455 ), .Q ( signal_22456 ) ) ;
    buf_clk cell_7769 ( .C ( clk ), .D ( signal_22461 ), .Q ( signal_22462 ) ) ;
    buf_clk cell_7775 ( .C ( clk ), .D ( signal_22467 ), .Q ( signal_22468 ) ) ;
    buf_clk cell_7781 ( .C ( clk ), .D ( signal_22473 ), .Q ( signal_22474 ) ) ;
    buf_clk cell_7789 ( .C ( clk ), .D ( signal_22481 ), .Q ( signal_22482 ) ) ;
    buf_clk cell_7797 ( .C ( clk ), .D ( signal_22489 ), .Q ( signal_22490 ) ) ;
    buf_clk cell_7805 ( .C ( clk ), .D ( signal_22497 ), .Q ( signal_22498 ) ) ;
    buf_clk cell_7813 ( .C ( clk ), .D ( signal_22505 ), .Q ( signal_22506 ) ) ;
    buf_clk cell_7821 ( .C ( clk ), .D ( signal_22513 ), .Q ( signal_22514 ) ) ;
    buf_clk cell_7831 ( .C ( clk ), .D ( signal_22523 ), .Q ( signal_22524 ) ) ;
    buf_clk cell_7841 ( .C ( clk ), .D ( signal_22533 ), .Q ( signal_22534 ) ) ;
    buf_clk cell_7851 ( .C ( clk ), .D ( signal_22543 ), .Q ( signal_22544 ) ) ;
    buf_clk cell_7861 ( .C ( clk ), .D ( signal_22553 ), .Q ( signal_22554 ) ) ;
    buf_clk cell_7871 ( .C ( clk ), .D ( signal_22563 ), .Q ( signal_22564 ) ) ;
    buf_clk cell_7879 ( .C ( clk ), .D ( signal_22571 ), .Q ( signal_22572 ) ) ;
    buf_clk cell_7887 ( .C ( clk ), .D ( signal_22579 ), .Q ( signal_22580 ) ) ;
    buf_clk cell_7895 ( .C ( clk ), .D ( signal_22587 ), .Q ( signal_22588 ) ) ;
    buf_clk cell_7903 ( .C ( clk ), .D ( signal_22595 ), .Q ( signal_22596 ) ) ;
    buf_clk cell_7911 ( .C ( clk ), .D ( signal_22603 ), .Q ( signal_22604 ) ) ;
    buf_clk cell_7917 ( .C ( clk ), .D ( signal_22609 ), .Q ( signal_22610 ) ) ;
    buf_clk cell_7923 ( .C ( clk ), .D ( signal_22615 ), .Q ( signal_22616 ) ) ;
    buf_clk cell_7929 ( .C ( clk ), .D ( signal_22621 ), .Q ( signal_22622 ) ) ;
    buf_clk cell_7935 ( .C ( clk ), .D ( signal_22627 ), .Q ( signal_22628 ) ) ;
    buf_clk cell_7941 ( .C ( clk ), .D ( signal_22633 ), .Q ( signal_22634 ) ) ;
    buf_clk cell_7947 ( .C ( clk ), .D ( signal_22639 ), .Q ( signal_22640 ) ) ;
    buf_clk cell_7953 ( .C ( clk ), .D ( signal_22645 ), .Q ( signal_22646 ) ) ;
    buf_clk cell_7959 ( .C ( clk ), .D ( signal_22651 ), .Q ( signal_22652 ) ) ;
    buf_clk cell_7965 ( .C ( clk ), .D ( signal_22657 ), .Q ( signal_22658 ) ) ;
    buf_clk cell_7971 ( .C ( clk ), .D ( signal_22663 ), .Q ( signal_22664 ) ) ;
    buf_clk cell_7985 ( .C ( clk ), .D ( signal_21263 ), .Q ( signal_22678 ) ) ;
    buf_clk cell_7989 ( .C ( clk ), .D ( signal_21269 ), .Q ( signal_22682 ) ) ;
    buf_clk cell_7993 ( .C ( clk ), .D ( signal_21275 ), .Q ( signal_22686 ) ) ;
    buf_clk cell_7997 ( .C ( clk ), .D ( signal_21281 ), .Q ( signal_22690 ) ) ;
    buf_clk cell_8001 ( .C ( clk ), .D ( signal_21287 ), .Q ( signal_22694 ) ) ;
    buf_clk cell_8005 ( .C ( clk ), .D ( signal_2253 ), .Q ( signal_22698 ) ) ;
    buf_clk cell_8009 ( .C ( clk ), .D ( signal_7668 ), .Q ( signal_22702 ) ) ;
    buf_clk cell_8013 ( .C ( clk ), .D ( signal_7669 ), .Q ( signal_22706 ) ) ;
    buf_clk cell_8017 ( .C ( clk ), .D ( signal_7670 ), .Q ( signal_22710 ) ) ;
    buf_clk cell_8021 ( .C ( clk ), .D ( signal_7671 ), .Q ( signal_22714 ) ) ;
    buf_clk cell_8027 ( .C ( clk ), .D ( signal_22719 ), .Q ( signal_22720 ) ) ;
    buf_clk cell_8033 ( .C ( clk ), .D ( signal_22725 ), .Q ( signal_22726 ) ) ;
    buf_clk cell_8039 ( .C ( clk ), .D ( signal_22731 ), .Q ( signal_22732 ) ) ;
    buf_clk cell_8045 ( .C ( clk ), .D ( signal_22737 ), .Q ( signal_22738 ) ) ;
    buf_clk cell_8051 ( .C ( clk ), .D ( signal_22743 ), .Q ( signal_22744 ) ) ;
    buf_clk cell_8067 ( .C ( clk ), .D ( signal_22759 ), .Q ( signal_22760 ) ) ;
    buf_clk cell_8073 ( .C ( clk ), .D ( signal_22765 ), .Q ( signal_22766 ) ) ;
    buf_clk cell_8079 ( .C ( clk ), .D ( signal_22771 ), .Q ( signal_22772 ) ) ;
    buf_clk cell_8085 ( .C ( clk ), .D ( signal_22777 ), .Q ( signal_22778 ) ) ;
    buf_clk cell_8091 ( .C ( clk ), .D ( signal_22783 ), .Q ( signal_22784 ) ) ;
    buf_clk cell_8095 ( .C ( clk ), .D ( signal_2208 ), .Q ( signal_22788 ) ) ;
    buf_clk cell_8099 ( .C ( clk ), .D ( signal_7488 ), .Q ( signal_22792 ) ) ;
    buf_clk cell_8103 ( .C ( clk ), .D ( signal_7489 ), .Q ( signal_22796 ) ) ;
    buf_clk cell_8107 ( .C ( clk ), .D ( signal_7490 ), .Q ( signal_22800 ) ) ;
    buf_clk cell_8111 ( .C ( clk ), .D ( signal_7491 ), .Q ( signal_22804 ) ) ;
    buf_clk cell_8117 ( .C ( clk ), .D ( signal_22809 ), .Q ( signal_22810 ) ) ;
    buf_clk cell_8123 ( .C ( clk ), .D ( signal_22815 ), .Q ( signal_22816 ) ) ;
    buf_clk cell_8129 ( .C ( clk ), .D ( signal_22821 ), .Q ( signal_22822 ) ) ;
    buf_clk cell_8135 ( .C ( clk ), .D ( signal_22827 ), .Q ( signal_22828 ) ) ;
    buf_clk cell_8141 ( .C ( clk ), .D ( signal_22833 ), .Q ( signal_22834 ) ) ;
    buf_clk cell_8155 ( .C ( clk ), .D ( signal_2249 ), .Q ( signal_22848 ) ) ;
    buf_clk cell_8159 ( .C ( clk ), .D ( signal_7652 ), .Q ( signal_22852 ) ) ;
    buf_clk cell_8163 ( .C ( clk ), .D ( signal_7653 ), .Q ( signal_22856 ) ) ;
    buf_clk cell_8167 ( .C ( clk ), .D ( signal_7654 ), .Q ( signal_22860 ) ) ;
    buf_clk cell_8171 ( .C ( clk ), .D ( signal_7655 ), .Q ( signal_22864 ) ) ;
    buf_clk cell_8175 ( .C ( clk ), .D ( signal_2161 ), .Q ( signal_22868 ) ) ;
    buf_clk cell_8181 ( .C ( clk ), .D ( signal_7300 ), .Q ( signal_22874 ) ) ;
    buf_clk cell_8187 ( .C ( clk ), .D ( signal_7301 ), .Q ( signal_22880 ) ) ;
    buf_clk cell_8193 ( .C ( clk ), .D ( signal_7302 ), .Q ( signal_22886 ) ) ;
    buf_clk cell_8199 ( .C ( clk ), .D ( signal_7303 ), .Q ( signal_22892 ) ) ;
    buf_clk cell_8207 ( .C ( clk ), .D ( signal_22899 ), .Q ( signal_22900 ) ) ;
    buf_clk cell_8215 ( .C ( clk ), .D ( signal_22907 ), .Q ( signal_22908 ) ) ;
    buf_clk cell_8223 ( .C ( clk ), .D ( signal_22915 ), .Q ( signal_22916 ) ) ;
    buf_clk cell_8231 ( .C ( clk ), .D ( signal_22923 ), .Q ( signal_22924 ) ) ;
    buf_clk cell_8239 ( .C ( clk ), .D ( signal_22931 ), .Q ( signal_22932 ) ) ;
    buf_clk cell_8245 ( .C ( clk ), .D ( signal_2199 ), .Q ( signal_22938 ) ) ;
    buf_clk cell_8251 ( .C ( clk ), .D ( signal_7452 ), .Q ( signal_22944 ) ) ;
    buf_clk cell_8257 ( .C ( clk ), .D ( signal_7453 ), .Q ( signal_22950 ) ) ;
    buf_clk cell_8263 ( .C ( clk ), .D ( signal_7454 ), .Q ( signal_22956 ) ) ;
    buf_clk cell_8269 ( .C ( clk ), .D ( signal_7455 ), .Q ( signal_22962 ) ) ;
    buf_clk cell_8279 ( .C ( clk ), .D ( signal_22971 ), .Q ( signal_22972 ) ) ;
    buf_clk cell_8289 ( .C ( clk ), .D ( signal_22981 ), .Q ( signal_22982 ) ) ;
    buf_clk cell_8299 ( .C ( clk ), .D ( signal_22991 ), .Q ( signal_22992 ) ) ;
    buf_clk cell_8309 ( .C ( clk ), .D ( signal_23001 ), .Q ( signal_23002 ) ) ;
    buf_clk cell_8319 ( .C ( clk ), .D ( signal_23011 ), .Q ( signal_23012 ) ) ;
    buf_clk cell_8325 ( .C ( clk ), .D ( signal_2255 ), .Q ( signal_23018 ) ) ;
    buf_clk cell_8331 ( .C ( clk ), .D ( signal_7676 ), .Q ( signal_23024 ) ) ;
    buf_clk cell_8337 ( .C ( clk ), .D ( signal_7677 ), .Q ( signal_23030 ) ) ;
    buf_clk cell_8343 ( .C ( clk ), .D ( signal_7678 ), .Q ( signal_23036 ) ) ;
    buf_clk cell_8349 ( .C ( clk ), .D ( signal_7679 ), .Q ( signal_23042 ) ) ;
    buf_clk cell_8377 ( .C ( clk ), .D ( signal_23069 ), .Q ( signal_23070 ) ) ;
    buf_clk cell_8385 ( .C ( clk ), .D ( signal_23077 ), .Q ( signal_23078 ) ) ;
    buf_clk cell_8393 ( .C ( clk ), .D ( signal_23085 ), .Q ( signal_23086 ) ) ;
    buf_clk cell_8401 ( .C ( clk ), .D ( signal_23093 ), .Q ( signal_23094 ) ) ;
    buf_clk cell_8409 ( .C ( clk ), .D ( signal_23101 ), .Q ( signal_23102 ) ) ;
    buf_clk cell_8415 ( .C ( clk ), .D ( signal_2183 ), .Q ( signal_23108 ) ) ;
    buf_clk cell_8421 ( .C ( clk ), .D ( signal_7388 ), .Q ( signal_23114 ) ) ;
    buf_clk cell_8427 ( .C ( clk ), .D ( signal_7389 ), .Q ( signal_23120 ) ) ;
    buf_clk cell_8433 ( .C ( clk ), .D ( signal_7390 ), .Q ( signal_23126 ) ) ;
    buf_clk cell_8439 ( .C ( clk ), .D ( signal_7391 ), .Q ( signal_23132 ) ) ;
    buf_clk cell_8447 ( .C ( clk ), .D ( signal_23139 ), .Q ( signal_23140 ) ) ;
    buf_clk cell_8455 ( .C ( clk ), .D ( signal_23147 ), .Q ( signal_23148 ) ) ;
    buf_clk cell_8463 ( .C ( clk ), .D ( signal_23155 ), .Q ( signal_23156 ) ) ;
    buf_clk cell_8471 ( .C ( clk ), .D ( signal_23163 ), .Q ( signal_23164 ) ) ;
    buf_clk cell_8479 ( .C ( clk ), .D ( signal_23171 ), .Q ( signal_23172 ) ) ;
    buf_clk cell_8485 ( .C ( clk ), .D ( signal_21339 ), .Q ( signal_23178 ) ) ;
    buf_clk cell_8491 ( .C ( clk ), .D ( signal_21341 ), .Q ( signal_23184 ) ) ;
    buf_clk cell_8497 ( .C ( clk ), .D ( signal_21343 ), .Q ( signal_23190 ) ) ;
    buf_clk cell_8503 ( .C ( clk ), .D ( signal_21345 ), .Q ( signal_23196 ) ) ;
    buf_clk cell_8509 ( .C ( clk ), .D ( signal_21347 ), .Q ( signal_23202 ) ) ;
    buf_clk cell_8517 ( .C ( clk ), .D ( signal_23209 ), .Q ( signal_23210 ) ) ;
    buf_clk cell_8525 ( .C ( clk ), .D ( signal_23217 ), .Q ( signal_23218 ) ) ;
    buf_clk cell_8533 ( .C ( clk ), .D ( signal_23225 ), .Q ( signal_23226 ) ) ;
    buf_clk cell_8541 ( .C ( clk ), .D ( signal_23233 ), .Q ( signal_23234 ) ) ;
    buf_clk cell_8549 ( .C ( clk ), .D ( signal_23241 ), .Q ( signal_23242 ) ) ;
    buf_clk cell_8575 ( .C ( clk ), .D ( signal_2252 ), .Q ( signal_23268 ) ) ;
    buf_clk cell_8581 ( .C ( clk ), .D ( signal_7664 ), .Q ( signal_23274 ) ) ;
    buf_clk cell_8587 ( .C ( clk ), .D ( signal_7665 ), .Q ( signal_23280 ) ) ;
    buf_clk cell_8593 ( .C ( clk ), .D ( signal_7666 ), .Q ( signal_23286 ) ) ;
    buf_clk cell_8599 ( .C ( clk ), .D ( signal_7667 ), .Q ( signal_23292 ) ) ;
    buf_clk cell_8605 ( .C ( clk ), .D ( signal_2160 ), .Q ( signal_23298 ) ) ;
    buf_clk cell_8611 ( .C ( clk ), .D ( signal_7296 ), .Q ( signal_23304 ) ) ;
    buf_clk cell_8617 ( .C ( clk ), .D ( signal_7297 ), .Q ( signal_23310 ) ) ;
    buf_clk cell_8623 ( .C ( clk ), .D ( signal_7298 ), .Q ( signal_23316 ) ) ;
    buf_clk cell_8629 ( .C ( clk ), .D ( signal_7299 ), .Q ( signal_23322 ) ) ;
    buf_clk cell_8675 ( .C ( clk ), .D ( signal_2202 ), .Q ( signal_23368 ) ) ;
    buf_clk cell_8683 ( .C ( clk ), .D ( signal_7464 ), .Q ( signal_23376 ) ) ;
    buf_clk cell_8691 ( .C ( clk ), .D ( signal_7465 ), .Q ( signal_23384 ) ) ;
    buf_clk cell_8699 ( .C ( clk ), .D ( signal_7466 ), .Q ( signal_23392 ) ) ;
    buf_clk cell_8707 ( .C ( clk ), .D ( signal_7467 ), .Q ( signal_23400 ) ) ;
    buf_clk cell_8719 ( .C ( clk ), .D ( signal_23411 ), .Q ( signal_23412 ) ) ;
    buf_clk cell_8731 ( .C ( clk ), .D ( signal_23423 ), .Q ( signal_23424 ) ) ;
    buf_clk cell_8743 ( .C ( clk ), .D ( signal_23435 ), .Q ( signal_23436 ) ) ;
    buf_clk cell_8755 ( .C ( clk ), .D ( signal_23447 ), .Q ( signal_23448 ) ) ;
    buf_clk cell_8767 ( .C ( clk ), .D ( signal_23459 ), .Q ( signal_23460 ) ) ;
    buf_clk cell_8841 ( .C ( clk ), .D ( signal_23533 ), .Q ( signal_23534 ) ) ;
    buf_clk cell_8855 ( .C ( clk ), .D ( signal_23547 ), .Q ( signal_23548 ) ) ;
    buf_clk cell_8869 ( .C ( clk ), .D ( signal_23561 ), .Q ( signal_23562 ) ) ;
    buf_clk cell_8883 ( .C ( clk ), .D ( signal_23575 ), .Q ( signal_23576 ) ) ;
    buf_clk cell_8897 ( .C ( clk ), .D ( signal_23589 ), .Q ( signal_23590 ) ) ;
    buf_clk cell_8905 ( .C ( clk ), .D ( signal_2154 ), .Q ( signal_23598 ) ) ;
    buf_clk cell_8913 ( .C ( clk ), .D ( signal_7272 ), .Q ( signal_23606 ) ) ;
    buf_clk cell_8921 ( .C ( clk ), .D ( signal_7273 ), .Q ( signal_23614 ) ) ;
    buf_clk cell_8929 ( .C ( clk ), .D ( signal_7274 ), .Q ( signal_23622 ) ) ;
    buf_clk cell_8937 ( .C ( clk ), .D ( signal_7275 ), .Q ( signal_23630 ) ) ;
    buf_clk cell_8951 ( .C ( clk ), .D ( signal_23643 ), .Q ( signal_23644 ) ) ;
    buf_clk cell_8965 ( .C ( clk ), .D ( signal_23657 ), .Q ( signal_23658 ) ) ;
    buf_clk cell_8979 ( .C ( clk ), .D ( signal_23671 ), .Q ( signal_23672 ) ) ;
    buf_clk cell_8993 ( .C ( clk ), .D ( signal_23685 ), .Q ( signal_23686 ) ) ;
    buf_clk cell_9007 ( .C ( clk ), .D ( signal_23699 ), .Q ( signal_23700 ) ) ;
    buf_clk cell_9015 ( .C ( clk ), .D ( signal_2149 ), .Q ( signal_23708 ) ) ;
    buf_clk cell_9023 ( .C ( clk ), .D ( signal_7252 ), .Q ( signal_23716 ) ) ;
    buf_clk cell_9031 ( .C ( clk ), .D ( signal_7253 ), .Q ( signal_23724 ) ) ;
    buf_clk cell_9039 ( .C ( clk ), .D ( signal_7254 ), .Q ( signal_23732 ) ) ;
    buf_clk cell_9047 ( .C ( clk ), .D ( signal_7255 ), .Q ( signal_23740 ) ) ;
    buf_clk cell_9075 ( .C ( clk ), .D ( signal_2152 ), .Q ( signal_23768 ) ) ;
    buf_clk cell_9085 ( .C ( clk ), .D ( signal_7264 ), .Q ( signal_23778 ) ) ;
    buf_clk cell_9095 ( .C ( clk ), .D ( signal_7265 ), .Q ( signal_23788 ) ) ;
    buf_clk cell_9105 ( .C ( clk ), .D ( signal_7266 ), .Q ( signal_23798 ) ) ;
    buf_clk cell_9115 ( .C ( clk ), .D ( signal_7267 ), .Q ( signal_23808 ) ) ;
    buf_clk cell_9151 ( .C ( clk ), .D ( signal_23843 ), .Q ( signal_23844 ) ) ;
    buf_clk cell_9167 ( .C ( clk ), .D ( signal_23859 ), .Q ( signal_23860 ) ) ;
    buf_clk cell_9183 ( .C ( clk ), .D ( signal_23875 ), .Q ( signal_23876 ) ) ;
    buf_clk cell_9199 ( .C ( clk ), .D ( signal_23891 ), .Q ( signal_23892 ) ) ;
    buf_clk cell_9215 ( .C ( clk ), .D ( signal_23907 ), .Q ( signal_23908 ) ) ;
    buf_clk cell_9251 ( .C ( clk ), .D ( signal_23943 ), .Q ( signal_23944 ) ) ;
    buf_clk cell_9267 ( .C ( clk ), .D ( signal_23959 ), .Q ( signal_23960 ) ) ;
    buf_clk cell_9283 ( .C ( clk ), .D ( signal_23975 ), .Q ( signal_23976 ) ) ;
    buf_clk cell_9299 ( .C ( clk ), .D ( signal_23991 ), .Q ( signal_23992 ) ) ;
    buf_clk cell_9315 ( .C ( clk ), .D ( signal_24007 ), .Q ( signal_24008 ) ) ;
    buf_clk cell_9325 ( .C ( clk ), .D ( signal_2257 ), .Q ( signal_24018 ) ) ;
    buf_clk cell_9335 ( .C ( clk ), .D ( signal_7684 ), .Q ( signal_24028 ) ) ;
    buf_clk cell_9345 ( .C ( clk ), .D ( signal_7685 ), .Q ( signal_24038 ) ) ;
    buf_clk cell_9355 ( .C ( clk ), .D ( signal_7686 ), .Q ( signal_24048 ) ) ;
    buf_clk cell_9365 ( .C ( clk ), .D ( signal_7687 ), .Q ( signal_24058 ) ) ;
    buf_clk cell_9559 ( .C ( clk ), .D ( signal_24251 ), .Q ( signal_24252 ) ) ;
    buf_clk cell_9575 ( .C ( clk ), .D ( signal_24267 ), .Q ( signal_24268 ) ) ;
    buf_clk cell_9591 ( .C ( clk ), .D ( signal_24283 ), .Q ( signal_24284 ) ) ;
    buf_clk cell_9607 ( .C ( clk ), .D ( signal_24299 ), .Q ( signal_24300 ) ) ;
    buf_clk cell_9623 ( .C ( clk ), .D ( signal_24315 ), .Q ( signal_24316 ) ) ;
    buf_clk cell_9641 ( .C ( clk ), .D ( signal_24333 ), .Q ( signal_24334 ) ) ;
    buf_clk cell_9659 ( .C ( clk ), .D ( signal_24351 ), .Q ( signal_24352 ) ) ;
    buf_clk cell_9677 ( .C ( clk ), .D ( signal_24369 ), .Q ( signal_24370 ) ) ;
    buf_clk cell_9695 ( .C ( clk ), .D ( signal_24387 ), .Q ( signal_24388 ) ) ;
    buf_clk cell_9713 ( .C ( clk ), .D ( signal_24405 ), .Q ( signal_24406 ) ) ;
    buf_clk cell_9891 ( .C ( clk ), .D ( signal_24583 ), .Q ( signal_24584 ) ) ;
    buf_clk cell_9911 ( .C ( clk ), .D ( signal_24603 ), .Q ( signal_24604 ) ) ;
    buf_clk cell_9931 ( .C ( clk ), .D ( signal_24623 ), .Q ( signal_24624 ) ) ;
    buf_clk cell_9951 ( .C ( clk ), .D ( signal_24643 ), .Q ( signal_24644 ) ) ;
    buf_clk cell_9971 ( .C ( clk ), .D ( signal_24663 ), .Q ( signal_24664 ) ) ;

    /* cells in depth 14 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2116 ( .a ({signal_20637, signal_20629, signal_20621, signal_20613, signal_20605}), .b ({signal_6871, signal_6870, signal_6869, signal_6868, signal_2053}), .clk ( clk ), .r ({Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290]}), .c ({signal_7183, signal_7182, signal_7181, signal_7180, signal_2131}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2118 ( .a ({signal_20657, signal_20653, signal_20649, signal_20645, signal_20641}), .b ({signal_6875, signal_6874, signal_6873, signal_6872, signal_2054}), .clk ( clk ), .r ({Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300]}), .c ({signal_7191, signal_7190, signal_7189, signal_7188, signal_2133}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2119 ( .a ({signal_20687, signal_20681, signal_20675, signal_20669, signal_20663}), .b ({signal_6879, signal_6878, signal_6877, signal_6876, signal_2055}), .clk ( clk ), .r ({Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310]}), .c ({signal_7195, signal_7194, signal_7193, signal_7192, signal_2134}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2121 ( .a ({signal_20717, signal_20711, signal_20705, signal_20699, signal_20693}), .b ({signal_6887, signal_6886, signal_6885, signal_6884, signal_2057}), .clk ( clk ), .r ({Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320]}), .c ({signal_7203, signal_7202, signal_7201, signal_7200, signal_2136}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2122 ( .a ({signal_20737, signal_20733, signal_20729, signal_20725, signal_20721}), .b ({signal_6895, signal_6894, signal_6893, signal_6892, signal_2059}), .clk ( clk ), .r ({Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330]}), .c ({signal_7207, signal_7206, signal_7205, signal_7204, signal_2137}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2123 ( .a ({signal_20767, signal_20761, signal_20755, signal_20749, signal_20743}), .b ({signal_6899, signal_6898, signal_6897, signal_6896, signal_2060}), .clk ( clk ), .r ({Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340]}), .c ({signal_7211, signal_7210, signal_7209, signal_7208, signal_2138}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2140 ( .a ({signal_7195, signal_7194, signal_7193, signal_7192, signal_2134}), .b ({signal_7279, signal_7278, signal_7277, signal_7276, signal_2155}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2162 ( .a ({signal_20787, signal_20783, signal_20779, signal_20775, signal_20771}), .b ({signal_6975, signal_6974, signal_6973, signal_6972, signal_2079}), .clk ( clk ), .r ({Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350]}), .c ({signal_7367, signal_7366, signal_7365, signal_7364, signal_2177}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2170 ( .a ({signal_20807, signal_20803, signal_20799, signal_20795, signal_20791}), .b ({signal_7111, signal_7110, signal_7109, signal_7108, signal_2113}), .clk ( clk ), .r ({Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360]}), .c ({signal_7399, signal_7398, signal_7397, signal_7396, signal_2185}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2172 ( .a ({signal_20817, signal_20815, signal_20813, signal_20811, signal_20809}), .b ({signal_7127, signal_7126, signal_7125, signal_7124, signal_2117}), .clk ( clk ), .r ({Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370]}), .c ({signal_7407, signal_7406, signal_7405, signal_7404, signal_2187}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2173 ( .a ({signal_20827, signal_20825, signal_20823, signal_20821, signal_20819}), .b ({signal_7007, signal_7006, signal_7005, signal_7004, signal_2087}), .clk ( clk ), .r ({Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380]}), .c ({signal_7411, signal_7410, signal_7409, signal_7408, signal_2188}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2174 ( .a ({signal_20857, signal_20851, signal_20845, signal_20839, signal_20833}), .b ({signal_7143, signal_7142, signal_7141, signal_7140, signal_2121}), .clk ( clk ), .r ({Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390]}), .c ({signal_7415, signal_7414, signal_7413, signal_7412, signal_2189}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2175 ( .a ({signal_20887, signal_20881, signal_20875, signal_20869, signal_20863}), .b ({signal_7147, signal_7146, signal_7145, signal_7144, signal_2122}), .clk ( clk ), .r ({Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400]}), .c ({signal_7419, signal_7418, signal_7417, signal_7416, signal_2190}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2176 ( .a ({signal_20917, signal_20911, signal_20905, signal_20899, signal_20893}), .b ({signal_7151, signal_7150, signal_7149, signal_7148, signal_2123}), .clk ( clk ), .r ({Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410]}), .c ({signal_7423, signal_7422, signal_7421, signal_7420, signal_2191}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2177 ( .a ({signal_6991, signal_6990, signal_6989, signal_6988, signal_2083}), .b ({signal_6883, signal_6882, signal_6881, signal_6880, signal_2056}), .clk ( clk ), .r ({Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420]}), .c ({signal_7427, signal_7426, signal_7425, signal_7424, signal_2192}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2178 ( .a ({signal_20927, signal_20925, signal_20923, signal_20921, signal_20919}), .b ({signal_7011, signal_7010, signal_7009, signal_7008, signal_2088}), .clk ( clk ), .r ({Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430]}), .c ({signal_7431, signal_7430, signal_7429, signal_7428, signal_2193}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2179 ( .a ({signal_20947, signal_20943, signal_20939, signal_20935, signal_20931}), .b ({signal_7171, signal_7170, signal_7169, signal_7168, signal_2128}), .clk ( clk ), .r ({Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440]}), .c ({signal_7435, signal_7434, signal_7433, signal_7432, signal_2194}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2190 ( .a ({signal_7367, signal_7366, signal_7365, signal_7364, signal_2177}), .b ({signal_7479, signal_7478, signal_7477, signal_7476, signal_2205}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2195 ( .a ({signal_7411, signal_7410, signal_7409, signal_7408, signal_2188}), .b ({signal_7499, signal_7498, signal_7497, signal_7496, signal_2210}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2196 ( .a ({signal_7419, signal_7418, signal_7417, signal_7416, signal_2190}), .b ({signal_7503, signal_7502, signal_7501, signal_7500, signal_2211}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2197 ( .a ({signal_7423, signal_7422, signal_7421, signal_7420, signal_2191}), .b ({signal_7507, signal_7506, signal_7505, signal_7504, signal_2212}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2198 ( .a ({signal_7431, signal_7430, signal_7429, signal_7428, signal_2193}), .b ({signal_7511, signal_7510, signal_7509, signal_7508, signal_2213}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2200 ( .a ({signal_20977, signal_20971, signal_20965, signal_20959, signal_20953}), .b ({signal_7287, signal_7286, signal_7285, signal_7284, signal_2157}), .clk ( clk ), .r ({Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450]}), .c ({signal_7519, signal_7518, signal_7517, signal_7516, signal_2215}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2207 ( .a ({signal_20987, signal_20985, signal_20983, signal_20981, signal_20979}), .b ({signal_7243, signal_7242, signal_7241, signal_7240, signal_2146}), .clk ( clk ), .r ({Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460]}), .c ({signal_7547, signal_7546, signal_7545, signal_7544, signal_2222}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2208 ( .a ({signal_21017, signal_21011, signal_21005, signal_20999, signal_20993}), .b ({signal_7315, signal_7314, signal_7313, signal_7312, signal_2164}), .clk ( clk ), .r ({Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470]}), .c ({signal_7551, signal_7550, signal_7549, signal_7548, signal_2223}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2209 ( .a ({signal_21027, signal_21025, signal_21023, signal_21021, signal_21019}), .b ({signal_7247, signal_7246, signal_7245, signal_7244, signal_2147}), .clk ( clk ), .r ({Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480]}), .c ({signal_7555, signal_7554, signal_7553, signal_7552, signal_2224}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2210 ( .a ({signal_21067, signal_21059, signal_21051, signal_21043, signal_21035}), .b ({signal_7319, signal_7318, signal_7317, signal_7316, signal_2165}), .clk ( clk ), .r ({Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490]}), .c ({signal_7559, signal_7558, signal_7557, signal_7556, signal_2225}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2211 ( .a ({signal_21087, signal_21083, signal_21079, signal_21075, signal_21071}), .b ({signal_7327, signal_7326, signal_7325, signal_7324, signal_2167}), .clk ( clk ), .r ({Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500]}), .c ({signal_7563, signal_7562, signal_7561, signal_7560, signal_2226}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2212 ( .a ({signal_7131, signal_7130, signal_7129, signal_7128, signal_2118}), .b ({signal_7331, signal_7330, signal_7329, signal_7328, signal_2168}), .clk ( clk ), .r ({Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510]}), .c ({signal_7567, signal_7566, signal_7565, signal_7564, signal_2227}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2214 ( .a ({signal_21107, signal_21103, signal_21099, signal_21095, signal_21091}), .b ({signal_7335, signal_7334, signal_7333, signal_7332, signal_2169}), .clk ( clk ), .r ({Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520]}), .c ({signal_7575, signal_7574, signal_7573, signal_7572, signal_2229}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2215 ( .a ({signal_7139, signal_7138, signal_7137, signal_7136, signal_2120}), .b ({signal_7339, signal_7338, signal_7337, signal_7336, signal_2170}), .clk ( clk ), .r ({Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530]}), .c ({signal_7579, signal_7578, signal_7577, signal_7576, signal_2230}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2216 ( .a ({signal_21137, signal_21131, signal_21125, signal_21119, signal_21113}), .b ({signal_7343, signal_7342, signal_7341, signal_7340, signal_2171}), .clk ( clk ), .r ({Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540]}), .c ({signal_7583, signal_7582, signal_7581, signal_7580, signal_2231}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2217 ( .a ({signal_21167, signal_21161, signal_21155, signal_21149, signal_21143}), .b ({signal_7351, signal_7350, signal_7349, signal_7348, signal_2173}), .clk ( clk ), .r ({Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550]}), .c ({signal_7587, signal_7586, signal_7585, signal_7584, signal_2232}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2218 ( .a ({signal_21187, signal_21183, signal_21179, signal_21175, signal_21171}), .b ({signal_7359, signal_7358, signal_7357, signal_7356, signal_2175}), .clk ( clk ), .r ({Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560]}), .c ({signal_7591, signal_7590, signal_7589, signal_7588, signal_2233}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2219 ( .a ({signal_21227, signal_21219, signal_21211, signal_21203, signal_21195}), .b ({signal_7363, signal_7362, signal_7361, signal_7360, signal_2176}), .clk ( clk ), .r ({Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570]}), .c ({signal_7595, signal_7594, signal_7593, signal_7592, signal_2234}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2220 ( .a ({signal_21257, signal_21251, signal_21245, signal_21239, signal_21233}), .b ({signal_7371, signal_7370, signal_7369, signal_7368, signal_2178}), .clk ( clk ), .r ({Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580]}), .c ({signal_7599, signal_7598, signal_7597, signal_7596, signal_2235}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2222 ( .a ({signal_7263, signal_7262, signal_7261, signal_7260, signal_2151}), .b ({signal_7167, signal_7166, signal_7165, signal_7164, signal_2127}), .clk ( clk ), .r ({Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590]}), .c ({signal_7607, signal_7606, signal_7605, signal_7604, signal_2237}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2223 ( .a ({signal_7271, signal_7270, signal_7269, signal_7268, signal_2153}), .b ({signal_7387, signal_7386, signal_7385, signal_7384, signal_2182}), .clk ( clk ), .r ({Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600]}), .c ({signal_7611, signal_7610, signal_7609, signal_7608, signal_2238}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2224 ( .a ({signal_21287, signal_21281, signal_21275, signal_21269, signal_21263}), .b ({signal_7395, signal_7394, signal_7393, signal_7392, signal_2184}), .clk ( clk ), .r ({Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610]}), .c ({signal_7615, signal_7614, signal_7613, signal_7612, signal_2239}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2239 ( .a ({signal_7551, signal_7550, signal_7549, signal_7548, signal_2223}), .b ({signal_7675, signal_7674, signal_7673, signal_7672, signal_2254}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2241 ( .a ({signal_7587, signal_7586, signal_7585, signal_7584, signal_2232}), .b ({signal_7683, signal_7682, signal_7681, signal_7680, signal_2256}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2243 ( .a ({signal_7615, signal_7614, signal_7613, signal_7612, signal_2239}), .b ({signal_7691, signal_7690, signal_7689, signal_7688, signal_2258}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2249 ( .a ({signal_7307, signal_7306, signal_7305, signal_7304, signal_2162}), .b ({signal_21297, signal_21295, signal_21293, signal_21291, signal_21289}), .clk ( clk ), .r ({Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620]}), .c ({signal_7715, signal_7714, signal_7713, signal_7712, signal_2264}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2250 ( .a ({signal_7235, signal_7234, signal_7233, signal_7232, signal_2144}), .b ({signal_7471, signal_7470, signal_7469, signal_7468, signal_2203}), .clk ( clk ), .r ({Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630]}), .c ({signal_7719, signal_7718, signal_7717, signal_7716, signal_2265}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2251 ( .a ({signal_21307, signal_21305, signal_21303, signal_21301, signal_21299}), .b ({signal_7475, signal_7474, signal_7473, signal_7472, signal_2204}), .clk ( clk ), .r ({Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640]}), .c ({signal_7723, signal_7722, signal_7721, signal_7720, signal_2266}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2252 ( .a ({signal_21337, signal_21331, signal_21325, signal_21319, signal_21313}), .b ({signal_7483, signal_7482, signal_7481, signal_7480, signal_2206}), .clk ( clk ), .r ({Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650]}), .c ({signal_7727, signal_7726, signal_7725, signal_7724, signal_2267}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2253 ( .a ({signal_21347, signal_21345, signal_21343, signal_21341, signal_21339}), .b ({signal_7487, signal_7486, signal_7485, signal_7484, signal_2207}), .clk ( clk ), .r ({Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660]}), .c ({signal_7731, signal_7730, signal_7729, signal_7728, signal_2268}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2254 ( .a ({signal_21357, signal_21355, signal_21353, signal_21351, signal_21349}), .b ({signal_7495, signal_7494, signal_7493, signal_7492, signal_2209}), .clk ( clk ), .r ({Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670]}), .c ({signal_7735, signal_7734, signal_7733, signal_7732, signal_2269}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2271 ( .a ({signal_7723, signal_7722, signal_7721, signal_7720, signal_2266}), .b ({signal_7803, signal_7802, signal_7801, signal_7800, signal_2286}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2272 ( .a ({signal_7727, signal_7726, signal_7725, signal_7724, signal_2267}), .b ({signal_7807, signal_7806, signal_7805, signal_7804, signal_2287}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2273 ( .a ({signal_7731, signal_7730, signal_7729, signal_7728, signal_2268}), .b ({signal_7811, signal_7810, signal_7809, signal_7808, signal_2288}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2274 ( .a ({signal_7735, signal_7734, signal_7733, signal_7732, signal_2269}), .b ({signal_7815, signal_7814, signal_7813, signal_7812, signal_2289}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2282 ( .a ({signal_7659, signal_7658, signal_7657, signal_7656, signal_2250}), .b ({signal_21387, signal_21381, signal_21375, signal_21369, signal_21363}), .clk ( clk ), .r ({Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680]}), .c ({signal_7847, signal_7846, signal_7845, signal_7844, signal_2297}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2283 ( .a ({signal_21347, signal_21345, signal_21343, signal_21341, signal_21339}), .b ({signal_7651, signal_7650, signal_7649, signal_7648, signal_2248}), .clk ( clk ), .r ({Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690]}), .c ({signal_7851, signal_7850, signal_7849, signal_7848, signal_2298}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2285 ( .a ({signal_21417, signal_21411, signal_21405, signal_21399, signal_21393}), .b ({signal_7711, signal_7710, signal_7709, signal_7708, signal_2263}), .clk ( clk ), .r ({Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700]}), .c ({signal_7859, signal_7858, signal_7857, signal_7856, signal_2300}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2286 ( .a ({signal_21437, signal_21433, signal_21429, signal_21425, signal_21421}), .b ({signal_7663, signal_7662, signal_7661, signal_7660, signal_2251}), .clk ( clk ), .r ({Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710]}), .c ({signal_7863, signal_7862, signal_7861, signal_7860, signal_2301}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2297 ( .a ({signal_7851, signal_7850, signal_7849, signal_7848, signal_2298}), .b ({signal_7907, signal_7906, signal_7905, signal_7904, signal_2312}) ) ;
    buf_clk cell_6754 ( .C ( clk ), .D ( signal_21446 ), .Q ( signal_21447 ) ) ;
    buf_clk cell_6764 ( .C ( clk ), .D ( signal_21456 ), .Q ( signal_21457 ) ) ;
    buf_clk cell_6774 ( .C ( clk ), .D ( signal_21466 ), .Q ( signal_21467 ) ) ;
    buf_clk cell_6784 ( .C ( clk ), .D ( signal_21476 ), .Q ( signal_21477 ) ) ;
    buf_clk cell_6794 ( .C ( clk ), .D ( signal_21486 ), .Q ( signal_21487 ) ) ;
    buf_clk cell_6800 ( .C ( clk ), .D ( signal_21492 ), .Q ( signal_21493 ) ) ;
    buf_clk cell_6806 ( .C ( clk ), .D ( signal_21498 ), .Q ( signal_21499 ) ) ;
    buf_clk cell_6812 ( .C ( clk ), .D ( signal_21504 ), .Q ( signal_21505 ) ) ;
    buf_clk cell_6818 ( .C ( clk ), .D ( signal_21510 ), .Q ( signal_21511 ) ) ;
    buf_clk cell_6824 ( .C ( clk ), .D ( signal_21516 ), .Q ( signal_21517 ) ) ;
    buf_clk cell_6832 ( .C ( clk ), .D ( signal_21524 ), .Q ( signal_21525 ) ) ;
    buf_clk cell_6840 ( .C ( clk ), .D ( signal_21532 ), .Q ( signal_21533 ) ) ;
    buf_clk cell_6848 ( .C ( clk ), .D ( signal_21540 ), .Q ( signal_21541 ) ) ;
    buf_clk cell_6856 ( .C ( clk ), .D ( signal_21548 ), .Q ( signal_21549 ) ) ;
    buf_clk cell_6864 ( .C ( clk ), .D ( signal_21556 ), .Q ( signal_21557 ) ) ;
    buf_clk cell_6872 ( .C ( clk ), .D ( signal_21564 ), .Q ( signal_21565 ) ) ;
    buf_clk cell_6880 ( .C ( clk ), .D ( signal_21572 ), .Q ( signal_21573 ) ) ;
    buf_clk cell_6888 ( .C ( clk ), .D ( signal_21580 ), .Q ( signal_21581 ) ) ;
    buf_clk cell_6896 ( .C ( clk ), .D ( signal_21588 ), .Q ( signal_21589 ) ) ;
    buf_clk cell_6904 ( .C ( clk ), .D ( signal_21596 ), .Q ( signal_21597 ) ) ;
    buf_clk cell_6908 ( .C ( clk ), .D ( signal_21600 ), .Q ( signal_21601 ) ) ;
    buf_clk cell_6912 ( .C ( clk ), .D ( signal_21604 ), .Q ( signal_21605 ) ) ;
    buf_clk cell_6916 ( .C ( clk ), .D ( signal_21608 ), .Q ( signal_21609 ) ) ;
    buf_clk cell_6920 ( .C ( clk ), .D ( signal_21612 ), .Q ( signal_21613 ) ) ;
    buf_clk cell_6924 ( .C ( clk ), .D ( signal_21616 ), .Q ( signal_21617 ) ) ;
    buf_clk cell_6928 ( .C ( clk ), .D ( signal_21620 ), .Q ( signal_21621 ) ) ;
    buf_clk cell_6932 ( .C ( clk ), .D ( signal_21624 ), .Q ( signal_21625 ) ) ;
    buf_clk cell_6936 ( .C ( clk ), .D ( signal_21628 ), .Q ( signal_21629 ) ) ;
    buf_clk cell_6940 ( .C ( clk ), .D ( signal_21632 ), .Q ( signal_21633 ) ) ;
    buf_clk cell_6944 ( .C ( clk ), .D ( signal_21636 ), .Q ( signal_21637 ) ) ;
    buf_clk cell_6946 ( .C ( clk ), .D ( signal_21638 ), .Q ( signal_21639 ) ) ;
    buf_clk cell_6948 ( .C ( clk ), .D ( signal_21640 ), .Q ( signal_21641 ) ) ;
    buf_clk cell_6950 ( .C ( clk ), .D ( signal_21642 ), .Q ( signal_21643 ) ) ;
    buf_clk cell_6952 ( .C ( clk ), .D ( signal_21644 ), .Q ( signal_21645 ) ) ;
    buf_clk cell_6954 ( .C ( clk ), .D ( signal_21646 ), .Q ( signal_21647 ) ) ;
    buf_clk cell_6956 ( .C ( clk ), .D ( signal_21648 ), .Q ( signal_21649 ) ) ;
    buf_clk cell_6958 ( .C ( clk ), .D ( signal_21650 ), .Q ( signal_21651 ) ) ;
    buf_clk cell_6960 ( .C ( clk ), .D ( signal_21652 ), .Q ( signal_21653 ) ) ;
    buf_clk cell_6962 ( .C ( clk ), .D ( signal_21654 ), .Q ( signal_21655 ) ) ;
    buf_clk cell_6964 ( .C ( clk ), .D ( signal_21656 ), .Q ( signal_21657 ) ) ;
    buf_clk cell_6968 ( .C ( clk ), .D ( signal_21660 ), .Q ( signal_21661 ) ) ;
    buf_clk cell_6972 ( .C ( clk ), .D ( signal_21664 ), .Q ( signal_21665 ) ) ;
    buf_clk cell_6976 ( .C ( clk ), .D ( signal_21668 ), .Q ( signal_21669 ) ) ;
    buf_clk cell_6980 ( .C ( clk ), .D ( signal_21672 ), .Q ( signal_21673 ) ) ;
    buf_clk cell_6984 ( .C ( clk ), .D ( signal_21676 ), .Q ( signal_21677 ) ) ;
    buf_clk cell_6994 ( .C ( clk ), .D ( signal_21686 ), .Q ( signal_21687 ) ) ;
    buf_clk cell_7004 ( .C ( clk ), .D ( signal_21696 ), .Q ( signal_21697 ) ) ;
    buf_clk cell_7014 ( .C ( clk ), .D ( signal_21706 ), .Q ( signal_21707 ) ) ;
    buf_clk cell_7024 ( .C ( clk ), .D ( signal_21716 ), .Q ( signal_21717 ) ) ;
    buf_clk cell_7034 ( .C ( clk ), .D ( signal_21726 ), .Q ( signal_21727 ) ) ;
    buf_clk cell_7040 ( .C ( clk ), .D ( signal_21732 ), .Q ( signal_21733 ) ) ;
    buf_clk cell_7046 ( .C ( clk ), .D ( signal_21738 ), .Q ( signal_21739 ) ) ;
    buf_clk cell_7052 ( .C ( clk ), .D ( signal_21744 ), .Q ( signal_21745 ) ) ;
    buf_clk cell_7058 ( .C ( clk ), .D ( signal_21750 ), .Q ( signal_21751 ) ) ;
    buf_clk cell_7064 ( .C ( clk ), .D ( signal_21756 ), .Q ( signal_21757 ) ) ;
    buf_clk cell_7066 ( .C ( clk ), .D ( signal_21758 ), .Q ( signal_21759 ) ) ;
    buf_clk cell_7068 ( .C ( clk ), .D ( signal_21760 ), .Q ( signal_21761 ) ) ;
    buf_clk cell_7070 ( .C ( clk ), .D ( signal_21762 ), .Q ( signal_21763 ) ) ;
    buf_clk cell_7072 ( .C ( clk ), .D ( signal_21764 ), .Q ( signal_21765 ) ) ;
    buf_clk cell_7074 ( .C ( clk ), .D ( signal_21766 ), .Q ( signal_21767 ) ) ;
    buf_clk cell_7082 ( .C ( clk ), .D ( signal_21774 ), .Q ( signal_21775 ) ) ;
    buf_clk cell_7090 ( .C ( clk ), .D ( signal_21782 ), .Q ( signal_21783 ) ) ;
    buf_clk cell_7098 ( .C ( clk ), .D ( signal_21790 ), .Q ( signal_21791 ) ) ;
    buf_clk cell_7106 ( .C ( clk ), .D ( signal_21798 ), .Q ( signal_21799 ) ) ;
    buf_clk cell_7114 ( .C ( clk ), .D ( signal_21806 ), .Q ( signal_21807 ) ) ;
    buf_clk cell_7120 ( .C ( clk ), .D ( signal_21812 ), .Q ( signal_21813 ) ) ;
    buf_clk cell_7126 ( .C ( clk ), .D ( signal_21818 ), .Q ( signal_21819 ) ) ;
    buf_clk cell_7132 ( .C ( clk ), .D ( signal_21824 ), .Q ( signal_21825 ) ) ;
    buf_clk cell_7138 ( .C ( clk ), .D ( signal_21830 ), .Q ( signal_21831 ) ) ;
    buf_clk cell_7144 ( .C ( clk ), .D ( signal_21836 ), .Q ( signal_21837 ) ) ;
    buf_clk cell_7152 ( .C ( clk ), .D ( signal_21844 ), .Q ( signal_21845 ) ) ;
    buf_clk cell_7160 ( .C ( clk ), .D ( signal_21852 ), .Q ( signal_21853 ) ) ;
    buf_clk cell_7168 ( .C ( clk ), .D ( signal_21860 ), .Q ( signal_21861 ) ) ;
    buf_clk cell_7176 ( .C ( clk ), .D ( signal_21868 ), .Q ( signal_21869 ) ) ;
    buf_clk cell_7184 ( .C ( clk ), .D ( signal_21876 ), .Q ( signal_21877 ) ) ;
    buf_clk cell_7192 ( .C ( clk ), .D ( signal_21884 ), .Q ( signal_21885 ) ) ;
    buf_clk cell_7200 ( .C ( clk ), .D ( signal_21892 ), .Q ( signal_21893 ) ) ;
    buf_clk cell_7208 ( .C ( clk ), .D ( signal_21900 ), .Q ( signal_21901 ) ) ;
    buf_clk cell_7216 ( .C ( clk ), .D ( signal_21908 ), .Q ( signal_21909 ) ) ;
    buf_clk cell_7224 ( .C ( clk ), .D ( signal_21916 ), .Q ( signal_21917 ) ) ;
    buf_clk cell_7232 ( .C ( clk ), .D ( signal_21924 ), .Q ( signal_21925 ) ) ;
    buf_clk cell_7240 ( .C ( clk ), .D ( signal_21932 ), .Q ( signal_21933 ) ) ;
    buf_clk cell_7248 ( .C ( clk ), .D ( signal_21940 ), .Q ( signal_21941 ) ) ;
    buf_clk cell_7256 ( .C ( clk ), .D ( signal_21948 ), .Q ( signal_21949 ) ) ;
    buf_clk cell_7264 ( .C ( clk ), .D ( signal_21956 ), .Q ( signal_21957 ) ) ;
    buf_clk cell_7274 ( .C ( clk ), .D ( signal_21966 ), .Q ( signal_21967 ) ) ;
    buf_clk cell_7284 ( .C ( clk ), .D ( signal_21976 ), .Q ( signal_21977 ) ) ;
    buf_clk cell_7294 ( .C ( clk ), .D ( signal_21986 ), .Q ( signal_21987 ) ) ;
    buf_clk cell_7304 ( .C ( clk ), .D ( signal_21996 ), .Q ( signal_21997 ) ) ;
    buf_clk cell_7314 ( .C ( clk ), .D ( signal_22006 ), .Q ( signal_22007 ) ) ;
    buf_clk cell_7322 ( .C ( clk ), .D ( signal_22014 ), .Q ( signal_22015 ) ) ;
    buf_clk cell_7330 ( .C ( clk ), .D ( signal_22022 ), .Q ( signal_22023 ) ) ;
    buf_clk cell_7338 ( .C ( clk ), .D ( signal_22030 ), .Q ( signal_22031 ) ) ;
    buf_clk cell_7346 ( .C ( clk ), .D ( signal_22038 ), .Q ( signal_22039 ) ) ;
    buf_clk cell_7354 ( .C ( clk ), .D ( signal_22046 ), .Q ( signal_22047 ) ) ;
    buf_clk cell_7362 ( .C ( clk ), .D ( signal_22054 ), .Q ( signal_22055 ) ) ;
    buf_clk cell_7370 ( .C ( clk ), .D ( signal_22062 ), .Q ( signal_22063 ) ) ;
    buf_clk cell_7378 ( .C ( clk ), .D ( signal_22070 ), .Q ( signal_22071 ) ) ;
    buf_clk cell_7386 ( .C ( clk ), .D ( signal_22078 ), .Q ( signal_22079 ) ) ;
    buf_clk cell_7394 ( .C ( clk ), .D ( signal_22086 ), .Q ( signal_22087 ) ) ;
    buf_clk cell_7396 ( .C ( clk ), .D ( signal_22088 ), .Q ( signal_22089 ) ) ;
    buf_clk cell_7398 ( .C ( clk ), .D ( signal_22090 ), .Q ( signal_22091 ) ) ;
    buf_clk cell_7400 ( .C ( clk ), .D ( signal_22092 ), .Q ( signal_22093 ) ) ;
    buf_clk cell_7402 ( .C ( clk ), .D ( signal_22094 ), .Q ( signal_22095 ) ) ;
    buf_clk cell_7404 ( .C ( clk ), .D ( signal_22096 ), .Q ( signal_22097 ) ) ;
    buf_clk cell_7412 ( .C ( clk ), .D ( signal_22104 ), .Q ( signal_22105 ) ) ;
    buf_clk cell_7420 ( .C ( clk ), .D ( signal_22112 ), .Q ( signal_22113 ) ) ;
    buf_clk cell_7428 ( .C ( clk ), .D ( signal_22120 ), .Q ( signal_22121 ) ) ;
    buf_clk cell_7436 ( .C ( clk ), .D ( signal_22128 ), .Q ( signal_22129 ) ) ;
    buf_clk cell_7444 ( .C ( clk ), .D ( signal_22136 ), .Q ( signal_22137 ) ) ;
    buf_clk cell_7452 ( .C ( clk ), .D ( signal_22144 ), .Q ( signal_22145 ) ) ;
    buf_clk cell_7460 ( .C ( clk ), .D ( signal_22152 ), .Q ( signal_22153 ) ) ;
    buf_clk cell_7468 ( .C ( clk ), .D ( signal_22160 ), .Q ( signal_22161 ) ) ;
    buf_clk cell_7476 ( .C ( clk ), .D ( signal_22168 ), .Q ( signal_22169 ) ) ;
    buf_clk cell_7484 ( .C ( clk ), .D ( signal_22176 ), .Q ( signal_22177 ) ) ;
    buf_clk cell_7492 ( .C ( clk ), .D ( signal_22184 ), .Q ( signal_22185 ) ) ;
    buf_clk cell_7500 ( .C ( clk ), .D ( signal_22192 ), .Q ( signal_22193 ) ) ;
    buf_clk cell_7508 ( .C ( clk ), .D ( signal_22200 ), .Q ( signal_22201 ) ) ;
    buf_clk cell_7516 ( .C ( clk ), .D ( signal_22208 ), .Q ( signal_22209 ) ) ;
    buf_clk cell_7524 ( .C ( clk ), .D ( signal_22216 ), .Q ( signal_22217 ) ) ;
    buf_clk cell_7528 ( .C ( clk ), .D ( signal_22220 ), .Q ( signal_22221 ) ) ;
    buf_clk cell_7534 ( .C ( clk ), .D ( signal_22226 ), .Q ( signal_22227 ) ) ;
    buf_clk cell_7540 ( .C ( clk ), .D ( signal_22232 ), .Q ( signal_22233 ) ) ;
    buf_clk cell_7546 ( .C ( clk ), .D ( signal_22238 ), .Q ( signal_22239 ) ) ;
    buf_clk cell_7552 ( .C ( clk ), .D ( signal_22244 ), .Q ( signal_22245 ) ) ;
    buf_clk cell_7560 ( .C ( clk ), .D ( signal_22252 ), .Q ( signal_22253 ) ) ;
    buf_clk cell_7568 ( .C ( clk ), .D ( signal_22260 ), .Q ( signal_22261 ) ) ;
    buf_clk cell_7576 ( .C ( clk ), .D ( signal_22268 ), .Q ( signal_22269 ) ) ;
    buf_clk cell_7584 ( .C ( clk ), .D ( signal_22276 ), .Q ( signal_22277 ) ) ;
    buf_clk cell_7592 ( .C ( clk ), .D ( signal_22284 ), .Q ( signal_22285 ) ) ;
    buf_clk cell_7598 ( .C ( clk ), .D ( signal_22290 ), .Q ( signal_22291 ) ) ;
    buf_clk cell_7604 ( .C ( clk ), .D ( signal_22296 ), .Q ( signal_22297 ) ) ;
    buf_clk cell_7610 ( .C ( clk ), .D ( signal_22302 ), .Q ( signal_22303 ) ) ;
    buf_clk cell_7616 ( .C ( clk ), .D ( signal_22308 ), .Q ( signal_22309 ) ) ;
    buf_clk cell_7622 ( .C ( clk ), .D ( signal_22314 ), .Q ( signal_22315 ) ) ;
    buf_clk cell_7628 ( .C ( clk ), .D ( signal_22320 ), .Q ( signal_22321 ) ) ;
    buf_clk cell_7634 ( .C ( clk ), .D ( signal_22326 ), .Q ( signal_22327 ) ) ;
    buf_clk cell_7640 ( .C ( clk ), .D ( signal_22332 ), .Q ( signal_22333 ) ) ;
    buf_clk cell_7646 ( .C ( clk ), .D ( signal_22338 ), .Q ( signal_22339 ) ) ;
    buf_clk cell_7652 ( .C ( clk ), .D ( signal_22344 ), .Q ( signal_22345 ) ) ;
    buf_clk cell_7660 ( .C ( clk ), .D ( signal_22352 ), .Q ( signal_22353 ) ) ;
    buf_clk cell_7668 ( .C ( clk ), .D ( signal_22360 ), .Q ( signal_22361 ) ) ;
    buf_clk cell_7676 ( .C ( clk ), .D ( signal_22368 ), .Q ( signal_22369 ) ) ;
    buf_clk cell_7684 ( .C ( clk ), .D ( signal_22376 ), .Q ( signal_22377 ) ) ;
    buf_clk cell_7692 ( .C ( clk ), .D ( signal_22384 ), .Q ( signal_22385 ) ) ;
    buf_clk cell_7702 ( .C ( clk ), .D ( signal_22394 ), .Q ( signal_22395 ) ) ;
    buf_clk cell_7712 ( .C ( clk ), .D ( signal_22404 ), .Q ( signal_22405 ) ) ;
    buf_clk cell_7722 ( .C ( clk ), .D ( signal_22414 ), .Q ( signal_22415 ) ) ;
    buf_clk cell_7732 ( .C ( clk ), .D ( signal_22424 ), .Q ( signal_22425 ) ) ;
    buf_clk cell_7742 ( .C ( clk ), .D ( signal_22434 ), .Q ( signal_22435 ) ) ;
    buf_clk cell_7758 ( .C ( clk ), .D ( signal_22450 ), .Q ( signal_22451 ) ) ;
    buf_clk cell_7764 ( .C ( clk ), .D ( signal_22456 ), .Q ( signal_22457 ) ) ;
    buf_clk cell_7770 ( .C ( clk ), .D ( signal_22462 ), .Q ( signal_22463 ) ) ;
    buf_clk cell_7776 ( .C ( clk ), .D ( signal_22468 ), .Q ( signal_22469 ) ) ;
    buf_clk cell_7782 ( .C ( clk ), .D ( signal_22474 ), .Q ( signal_22475 ) ) ;
    buf_clk cell_7790 ( .C ( clk ), .D ( signal_22482 ), .Q ( signal_22483 ) ) ;
    buf_clk cell_7798 ( .C ( clk ), .D ( signal_22490 ), .Q ( signal_22491 ) ) ;
    buf_clk cell_7806 ( .C ( clk ), .D ( signal_22498 ), .Q ( signal_22499 ) ) ;
    buf_clk cell_7814 ( .C ( clk ), .D ( signal_22506 ), .Q ( signal_22507 ) ) ;
    buf_clk cell_7822 ( .C ( clk ), .D ( signal_22514 ), .Q ( signal_22515 ) ) ;
    buf_clk cell_7832 ( .C ( clk ), .D ( signal_22524 ), .Q ( signal_22525 ) ) ;
    buf_clk cell_7842 ( .C ( clk ), .D ( signal_22534 ), .Q ( signal_22535 ) ) ;
    buf_clk cell_7852 ( .C ( clk ), .D ( signal_22544 ), .Q ( signal_22545 ) ) ;
    buf_clk cell_7862 ( .C ( clk ), .D ( signal_22554 ), .Q ( signal_22555 ) ) ;
    buf_clk cell_7872 ( .C ( clk ), .D ( signal_22564 ), .Q ( signal_22565 ) ) ;
    buf_clk cell_7880 ( .C ( clk ), .D ( signal_22572 ), .Q ( signal_22573 ) ) ;
    buf_clk cell_7888 ( .C ( clk ), .D ( signal_22580 ), .Q ( signal_22581 ) ) ;
    buf_clk cell_7896 ( .C ( clk ), .D ( signal_22588 ), .Q ( signal_22589 ) ) ;
    buf_clk cell_7904 ( .C ( clk ), .D ( signal_22596 ), .Q ( signal_22597 ) ) ;
    buf_clk cell_7912 ( .C ( clk ), .D ( signal_22604 ), .Q ( signal_22605 ) ) ;
    buf_clk cell_7918 ( .C ( clk ), .D ( signal_22610 ), .Q ( signal_22611 ) ) ;
    buf_clk cell_7924 ( .C ( clk ), .D ( signal_22616 ), .Q ( signal_22617 ) ) ;
    buf_clk cell_7930 ( .C ( clk ), .D ( signal_22622 ), .Q ( signal_22623 ) ) ;
    buf_clk cell_7936 ( .C ( clk ), .D ( signal_22628 ), .Q ( signal_22629 ) ) ;
    buf_clk cell_7942 ( .C ( clk ), .D ( signal_22634 ), .Q ( signal_22635 ) ) ;
    buf_clk cell_7948 ( .C ( clk ), .D ( signal_22640 ), .Q ( signal_22641 ) ) ;
    buf_clk cell_7954 ( .C ( clk ), .D ( signal_22646 ), .Q ( signal_22647 ) ) ;
    buf_clk cell_7960 ( .C ( clk ), .D ( signal_22652 ), .Q ( signal_22653 ) ) ;
    buf_clk cell_7966 ( .C ( clk ), .D ( signal_22658 ), .Q ( signal_22659 ) ) ;
    buf_clk cell_7972 ( .C ( clk ), .D ( signal_22664 ), .Q ( signal_22665 ) ) ;
    buf_clk cell_7986 ( .C ( clk ), .D ( signal_22678 ), .Q ( signal_22679 ) ) ;
    buf_clk cell_7990 ( .C ( clk ), .D ( signal_22682 ), .Q ( signal_22683 ) ) ;
    buf_clk cell_7994 ( .C ( clk ), .D ( signal_22686 ), .Q ( signal_22687 ) ) ;
    buf_clk cell_7998 ( .C ( clk ), .D ( signal_22690 ), .Q ( signal_22691 ) ) ;
    buf_clk cell_8002 ( .C ( clk ), .D ( signal_22694 ), .Q ( signal_22695 ) ) ;
    buf_clk cell_8006 ( .C ( clk ), .D ( signal_22698 ), .Q ( signal_22699 ) ) ;
    buf_clk cell_8010 ( .C ( clk ), .D ( signal_22702 ), .Q ( signal_22703 ) ) ;
    buf_clk cell_8014 ( .C ( clk ), .D ( signal_22706 ), .Q ( signal_22707 ) ) ;
    buf_clk cell_8018 ( .C ( clk ), .D ( signal_22710 ), .Q ( signal_22711 ) ) ;
    buf_clk cell_8022 ( .C ( clk ), .D ( signal_22714 ), .Q ( signal_22715 ) ) ;
    buf_clk cell_8028 ( .C ( clk ), .D ( signal_22720 ), .Q ( signal_22721 ) ) ;
    buf_clk cell_8034 ( .C ( clk ), .D ( signal_22726 ), .Q ( signal_22727 ) ) ;
    buf_clk cell_8040 ( .C ( clk ), .D ( signal_22732 ), .Q ( signal_22733 ) ) ;
    buf_clk cell_8046 ( .C ( clk ), .D ( signal_22738 ), .Q ( signal_22739 ) ) ;
    buf_clk cell_8052 ( .C ( clk ), .D ( signal_22744 ), .Q ( signal_22745 ) ) ;
    buf_clk cell_8068 ( .C ( clk ), .D ( signal_22760 ), .Q ( signal_22761 ) ) ;
    buf_clk cell_8074 ( .C ( clk ), .D ( signal_22766 ), .Q ( signal_22767 ) ) ;
    buf_clk cell_8080 ( .C ( clk ), .D ( signal_22772 ), .Q ( signal_22773 ) ) ;
    buf_clk cell_8086 ( .C ( clk ), .D ( signal_22778 ), .Q ( signal_22779 ) ) ;
    buf_clk cell_8092 ( .C ( clk ), .D ( signal_22784 ), .Q ( signal_22785 ) ) ;
    buf_clk cell_8096 ( .C ( clk ), .D ( signal_22788 ), .Q ( signal_22789 ) ) ;
    buf_clk cell_8100 ( .C ( clk ), .D ( signal_22792 ), .Q ( signal_22793 ) ) ;
    buf_clk cell_8104 ( .C ( clk ), .D ( signal_22796 ), .Q ( signal_22797 ) ) ;
    buf_clk cell_8108 ( .C ( clk ), .D ( signal_22800 ), .Q ( signal_22801 ) ) ;
    buf_clk cell_8112 ( .C ( clk ), .D ( signal_22804 ), .Q ( signal_22805 ) ) ;
    buf_clk cell_8118 ( .C ( clk ), .D ( signal_22810 ), .Q ( signal_22811 ) ) ;
    buf_clk cell_8124 ( .C ( clk ), .D ( signal_22816 ), .Q ( signal_22817 ) ) ;
    buf_clk cell_8130 ( .C ( clk ), .D ( signal_22822 ), .Q ( signal_22823 ) ) ;
    buf_clk cell_8136 ( .C ( clk ), .D ( signal_22828 ), .Q ( signal_22829 ) ) ;
    buf_clk cell_8142 ( .C ( clk ), .D ( signal_22834 ), .Q ( signal_22835 ) ) ;
    buf_clk cell_8156 ( .C ( clk ), .D ( signal_22848 ), .Q ( signal_22849 ) ) ;
    buf_clk cell_8160 ( .C ( clk ), .D ( signal_22852 ), .Q ( signal_22853 ) ) ;
    buf_clk cell_8164 ( .C ( clk ), .D ( signal_22856 ), .Q ( signal_22857 ) ) ;
    buf_clk cell_8168 ( .C ( clk ), .D ( signal_22860 ), .Q ( signal_22861 ) ) ;
    buf_clk cell_8172 ( .C ( clk ), .D ( signal_22864 ), .Q ( signal_22865 ) ) ;
    buf_clk cell_8176 ( .C ( clk ), .D ( signal_22868 ), .Q ( signal_22869 ) ) ;
    buf_clk cell_8182 ( .C ( clk ), .D ( signal_22874 ), .Q ( signal_22875 ) ) ;
    buf_clk cell_8188 ( .C ( clk ), .D ( signal_22880 ), .Q ( signal_22881 ) ) ;
    buf_clk cell_8194 ( .C ( clk ), .D ( signal_22886 ), .Q ( signal_22887 ) ) ;
    buf_clk cell_8200 ( .C ( clk ), .D ( signal_22892 ), .Q ( signal_22893 ) ) ;
    buf_clk cell_8208 ( .C ( clk ), .D ( signal_22900 ), .Q ( signal_22901 ) ) ;
    buf_clk cell_8216 ( .C ( clk ), .D ( signal_22908 ), .Q ( signal_22909 ) ) ;
    buf_clk cell_8224 ( .C ( clk ), .D ( signal_22916 ), .Q ( signal_22917 ) ) ;
    buf_clk cell_8232 ( .C ( clk ), .D ( signal_22924 ), .Q ( signal_22925 ) ) ;
    buf_clk cell_8240 ( .C ( clk ), .D ( signal_22932 ), .Q ( signal_22933 ) ) ;
    buf_clk cell_8246 ( .C ( clk ), .D ( signal_22938 ), .Q ( signal_22939 ) ) ;
    buf_clk cell_8252 ( .C ( clk ), .D ( signal_22944 ), .Q ( signal_22945 ) ) ;
    buf_clk cell_8258 ( .C ( clk ), .D ( signal_22950 ), .Q ( signal_22951 ) ) ;
    buf_clk cell_8264 ( .C ( clk ), .D ( signal_22956 ), .Q ( signal_22957 ) ) ;
    buf_clk cell_8270 ( .C ( clk ), .D ( signal_22962 ), .Q ( signal_22963 ) ) ;
    buf_clk cell_8280 ( .C ( clk ), .D ( signal_22972 ), .Q ( signal_22973 ) ) ;
    buf_clk cell_8290 ( .C ( clk ), .D ( signal_22982 ), .Q ( signal_22983 ) ) ;
    buf_clk cell_8300 ( .C ( clk ), .D ( signal_22992 ), .Q ( signal_22993 ) ) ;
    buf_clk cell_8310 ( .C ( clk ), .D ( signal_23002 ), .Q ( signal_23003 ) ) ;
    buf_clk cell_8320 ( .C ( clk ), .D ( signal_23012 ), .Q ( signal_23013 ) ) ;
    buf_clk cell_8326 ( .C ( clk ), .D ( signal_23018 ), .Q ( signal_23019 ) ) ;
    buf_clk cell_8332 ( .C ( clk ), .D ( signal_23024 ), .Q ( signal_23025 ) ) ;
    buf_clk cell_8338 ( .C ( clk ), .D ( signal_23030 ), .Q ( signal_23031 ) ) ;
    buf_clk cell_8344 ( .C ( clk ), .D ( signal_23036 ), .Q ( signal_23037 ) ) ;
    buf_clk cell_8350 ( .C ( clk ), .D ( signal_23042 ), .Q ( signal_23043 ) ) ;
    buf_clk cell_8378 ( .C ( clk ), .D ( signal_23070 ), .Q ( signal_23071 ) ) ;
    buf_clk cell_8386 ( .C ( clk ), .D ( signal_23078 ), .Q ( signal_23079 ) ) ;
    buf_clk cell_8394 ( .C ( clk ), .D ( signal_23086 ), .Q ( signal_23087 ) ) ;
    buf_clk cell_8402 ( .C ( clk ), .D ( signal_23094 ), .Q ( signal_23095 ) ) ;
    buf_clk cell_8410 ( .C ( clk ), .D ( signal_23102 ), .Q ( signal_23103 ) ) ;
    buf_clk cell_8416 ( .C ( clk ), .D ( signal_23108 ), .Q ( signal_23109 ) ) ;
    buf_clk cell_8422 ( .C ( clk ), .D ( signal_23114 ), .Q ( signal_23115 ) ) ;
    buf_clk cell_8428 ( .C ( clk ), .D ( signal_23120 ), .Q ( signal_23121 ) ) ;
    buf_clk cell_8434 ( .C ( clk ), .D ( signal_23126 ), .Q ( signal_23127 ) ) ;
    buf_clk cell_8440 ( .C ( clk ), .D ( signal_23132 ), .Q ( signal_23133 ) ) ;
    buf_clk cell_8448 ( .C ( clk ), .D ( signal_23140 ), .Q ( signal_23141 ) ) ;
    buf_clk cell_8456 ( .C ( clk ), .D ( signal_23148 ), .Q ( signal_23149 ) ) ;
    buf_clk cell_8464 ( .C ( clk ), .D ( signal_23156 ), .Q ( signal_23157 ) ) ;
    buf_clk cell_8472 ( .C ( clk ), .D ( signal_23164 ), .Q ( signal_23165 ) ) ;
    buf_clk cell_8480 ( .C ( clk ), .D ( signal_23172 ), .Q ( signal_23173 ) ) ;
    buf_clk cell_8486 ( .C ( clk ), .D ( signal_23178 ), .Q ( signal_23179 ) ) ;
    buf_clk cell_8492 ( .C ( clk ), .D ( signal_23184 ), .Q ( signal_23185 ) ) ;
    buf_clk cell_8498 ( .C ( clk ), .D ( signal_23190 ), .Q ( signal_23191 ) ) ;
    buf_clk cell_8504 ( .C ( clk ), .D ( signal_23196 ), .Q ( signal_23197 ) ) ;
    buf_clk cell_8510 ( .C ( clk ), .D ( signal_23202 ), .Q ( signal_23203 ) ) ;
    buf_clk cell_8518 ( .C ( clk ), .D ( signal_23210 ), .Q ( signal_23211 ) ) ;
    buf_clk cell_8526 ( .C ( clk ), .D ( signal_23218 ), .Q ( signal_23219 ) ) ;
    buf_clk cell_8534 ( .C ( clk ), .D ( signal_23226 ), .Q ( signal_23227 ) ) ;
    buf_clk cell_8542 ( .C ( clk ), .D ( signal_23234 ), .Q ( signal_23235 ) ) ;
    buf_clk cell_8550 ( .C ( clk ), .D ( signal_23242 ), .Q ( signal_23243 ) ) ;
    buf_clk cell_8576 ( .C ( clk ), .D ( signal_23268 ), .Q ( signal_23269 ) ) ;
    buf_clk cell_8582 ( .C ( clk ), .D ( signal_23274 ), .Q ( signal_23275 ) ) ;
    buf_clk cell_8588 ( .C ( clk ), .D ( signal_23280 ), .Q ( signal_23281 ) ) ;
    buf_clk cell_8594 ( .C ( clk ), .D ( signal_23286 ), .Q ( signal_23287 ) ) ;
    buf_clk cell_8600 ( .C ( clk ), .D ( signal_23292 ), .Q ( signal_23293 ) ) ;
    buf_clk cell_8606 ( .C ( clk ), .D ( signal_23298 ), .Q ( signal_23299 ) ) ;
    buf_clk cell_8612 ( .C ( clk ), .D ( signal_23304 ), .Q ( signal_23305 ) ) ;
    buf_clk cell_8618 ( .C ( clk ), .D ( signal_23310 ), .Q ( signal_23311 ) ) ;
    buf_clk cell_8624 ( .C ( clk ), .D ( signal_23316 ), .Q ( signal_23317 ) ) ;
    buf_clk cell_8630 ( .C ( clk ), .D ( signal_23322 ), .Q ( signal_23323 ) ) ;
    buf_clk cell_8676 ( .C ( clk ), .D ( signal_23368 ), .Q ( signal_23369 ) ) ;
    buf_clk cell_8684 ( .C ( clk ), .D ( signal_23376 ), .Q ( signal_23377 ) ) ;
    buf_clk cell_8692 ( .C ( clk ), .D ( signal_23384 ), .Q ( signal_23385 ) ) ;
    buf_clk cell_8700 ( .C ( clk ), .D ( signal_23392 ), .Q ( signal_23393 ) ) ;
    buf_clk cell_8708 ( .C ( clk ), .D ( signal_23400 ), .Q ( signal_23401 ) ) ;
    buf_clk cell_8720 ( .C ( clk ), .D ( signal_23412 ), .Q ( signal_23413 ) ) ;
    buf_clk cell_8732 ( .C ( clk ), .D ( signal_23424 ), .Q ( signal_23425 ) ) ;
    buf_clk cell_8744 ( .C ( clk ), .D ( signal_23436 ), .Q ( signal_23437 ) ) ;
    buf_clk cell_8756 ( .C ( clk ), .D ( signal_23448 ), .Q ( signal_23449 ) ) ;
    buf_clk cell_8768 ( .C ( clk ), .D ( signal_23460 ), .Q ( signal_23461 ) ) ;
    buf_clk cell_8842 ( .C ( clk ), .D ( signal_23534 ), .Q ( signal_23535 ) ) ;
    buf_clk cell_8856 ( .C ( clk ), .D ( signal_23548 ), .Q ( signal_23549 ) ) ;
    buf_clk cell_8870 ( .C ( clk ), .D ( signal_23562 ), .Q ( signal_23563 ) ) ;
    buf_clk cell_8884 ( .C ( clk ), .D ( signal_23576 ), .Q ( signal_23577 ) ) ;
    buf_clk cell_8898 ( .C ( clk ), .D ( signal_23590 ), .Q ( signal_23591 ) ) ;
    buf_clk cell_8906 ( .C ( clk ), .D ( signal_23598 ), .Q ( signal_23599 ) ) ;
    buf_clk cell_8914 ( .C ( clk ), .D ( signal_23606 ), .Q ( signal_23607 ) ) ;
    buf_clk cell_8922 ( .C ( clk ), .D ( signal_23614 ), .Q ( signal_23615 ) ) ;
    buf_clk cell_8930 ( .C ( clk ), .D ( signal_23622 ), .Q ( signal_23623 ) ) ;
    buf_clk cell_8938 ( .C ( clk ), .D ( signal_23630 ), .Q ( signal_23631 ) ) ;
    buf_clk cell_8952 ( .C ( clk ), .D ( signal_23644 ), .Q ( signal_23645 ) ) ;
    buf_clk cell_8966 ( .C ( clk ), .D ( signal_23658 ), .Q ( signal_23659 ) ) ;
    buf_clk cell_8980 ( .C ( clk ), .D ( signal_23672 ), .Q ( signal_23673 ) ) ;
    buf_clk cell_8994 ( .C ( clk ), .D ( signal_23686 ), .Q ( signal_23687 ) ) ;
    buf_clk cell_9008 ( .C ( clk ), .D ( signal_23700 ), .Q ( signal_23701 ) ) ;
    buf_clk cell_9016 ( .C ( clk ), .D ( signal_23708 ), .Q ( signal_23709 ) ) ;
    buf_clk cell_9024 ( .C ( clk ), .D ( signal_23716 ), .Q ( signal_23717 ) ) ;
    buf_clk cell_9032 ( .C ( clk ), .D ( signal_23724 ), .Q ( signal_23725 ) ) ;
    buf_clk cell_9040 ( .C ( clk ), .D ( signal_23732 ), .Q ( signal_23733 ) ) ;
    buf_clk cell_9048 ( .C ( clk ), .D ( signal_23740 ), .Q ( signal_23741 ) ) ;
    buf_clk cell_9076 ( .C ( clk ), .D ( signal_23768 ), .Q ( signal_23769 ) ) ;
    buf_clk cell_9086 ( .C ( clk ), .D ( signal_23778 ), .Q ( signal_23779 ) ) ;
    buf_clk cell_9096 ( .C ( clk ), .D ( signal_23788 ), .Q ( signal_23789 ) ) ;
    buf_clk cell_9106 ( .C ( clk ), .D ( signal_23798 ), .Q ( signal_23799 ) ) ;
    buf_clk cell_9116 ( .C ( clk ), .D ( signal_23808 ), .Q ( signal_23809 ) ) ;
    buf_clk cell_9152 ( .C ( clk ), .D ( signal_23844 ), .Q ( signal_23845 ) ) ;
    buf_clk cell_9168 ( .C ( clk ), .D ( signal_23860 ), .Q ( signal_23861 ) ) ;
    buf_clk cell_9184 ( .C ( clk ), .D ( signal_23876 ), .Q ( signal_23877 ) ) ;
    buf_clk cell_9200 ( .C ( clk ), .D ( signal_23892 ), .Q ( signal_23893 ) ) ;
    buf_clk cell_9216 ( .C ( clk ), .D ( signal_23908 ), .Q ( signal_23909 ) ) ;
    buf_clk cell_9252 ( .C ( clk ), .D ( signal_23944 ), .Q ( signal_23945 ) ) ;
    buf_clk cell_9268 ( .C ( clk ), .D ( signal_23960 ), .Q ( signal_23961 ) ) ;
    buf_clk cell_9284 ( .C ( clk ), .D ( signal_23976 ), .Q ( signal_23977 ) ) ;
    buf_clk cell_9300 ( .C ( clk ), .D ( signal_23992 ), .Q ( signal_23993 ) ) ;
    buf_clk cell_9316 ( .C ( clk ), .D ( signal_24008 ), .Q ( signal_24009 ) ) ;
    buf_clk cell_9326 ( .C ( clk ), .D ( signal_24018 ), .Q ( signal_24019 ) ) ;
    buf_clk cell_9336 ( .C ( clk ), .D ( signal_24028 ), .Q ( signal_24029 ) ) ;
    buf_clk cell_9346 ( .C ( clk ), .D ( signal_24038 ), .Q ( signal_24039 ) ) ;
    buf_clk cell_9356 ( .C ( clk ), .D ( signal_24048 ), .Q ( signal_24049 ) ) ;
    buf_clk cell_9366 ( .C ( clk ), .D ( signal_24058 ), .Q ( signal_24059 ) ) ;
    buf_clk cell_9560 ( .C ( clk ), .D ( signal_24252 ), .Q ( signal_24253 ) ) ;
    buf_clk cell_9576 ( .C ( clk ), .D ( signal_24268 ), .Q ( signal_24269 ) ) ;
    buf_clk cell_9592 ( .C ( clk ), .D ( signal_24284 ), .Q ( signal_24285 ) ) ;
    buf_clk cell_9608 ( .C ( clk ), .D ( signal_24300 ), .Q ( signal_24301 ) ) ;
    buf_clk cell_9624 ( .C ( clk ), .D ( signal_24316 ), .Q ( signal_24317 ) ) ;
    buf_clk cell_9642 ( .C ( clk ), .D ( signal_24334 ), .Q ( signal_24335 ) ) ;
    buf_clk cell_9660 ( .C ( clk ), .D ( signal_24352 ), .Q ( signal_24353 ) ) ;
    buf_clk cell_9678 ( .C ( clk ), .D ( signal_24370 ), .Q ( signal_24371 ) ) ;
    buf_clk cell_9696 ( .C ( clk ), .D ( signal_24388 ), .Q ( signal_24389 ) ) ;
    buf_clk cell_9714 ( .C ( clk ), .D ( signal_24406 ), .Q ( signal_24407 ) ) ;
    buf_clk cell_9892 ( .C ( clk ), .D ( signal_24584 ), .Q ( signal_24585 ) ) ;
    buf_clk cell_9912 ( .C ( clk ), .D ( signal_24604 ), .Q ( signal_24605 ) ) ;
    buf_clk cell_9932 ( .C ( clk ), .D ( signal_24624 ), .Q ( signal_24625 ) ) ;
    buf_clk cell_9952 ( .C ( clk ), .D ( signal_24644 ), .Q ( signal_24645 ) ) ;
    buf_clk cell_9972 ( .C ( clk ), .D ( signal_24664 ), .Q ( signal_24665 ) ) ;

    /* cells in depth 15 */
    buf_clk cell_7529 ( .C ( clk ), .D ( signal_22221 ), .Q ( signal_22222 ) ) ;
    buf_clk cell_7535 ( .C ( clk ), .D ( signal_22227 ), .Q ( signal_22228 ) ) ;
    buf_clk cell_7541 ( .C ( clk ), .D ( signal_22233 ), .Q ( signal_22234 ) ) ;
    buf_clk cell_7547 ( .C ( clk ), .D ( signal_22239 ), .Q ( signal_22240 ) ) ;
    buf_clk cell_7553 ( .C ( clk ), .D ( signal_22245 ), .Q ( signal_22246 ) ) ;
    buf_clk cell_7561 ( .C ( clk ), .D ( signal_22253 ), .Q ( signal_22254 ) ) ;
    buf_clk cell_7569 ( .C ( clk ), .D ( signal_22261 ), .Q ( signal_22262 ) ) ;
    buf_clk cell_7577 ( .C ( clk ), .D ( signal_22269 ), .Q ( signal_22270 ) ) ;
    buf_clk cell_7585 ( .C ( clk ), .D ( signal_22277 ), .Q ( signal_22278 ) ) ;
    buf_clk cell_7593 ( .C ( clk ), .D ( signal_22285 ), .Q ( signal_22286 ) ) ;
    buf_clk cell_7599 ( .C ( clk ), .D ( signal_22291 ), .Q ( signal_22292 ) ) ;
    buf_clk cell_7605 ( .C ( clk ), .D ( signal_22297 ), .Q ( signal_22298 ) ) ;
    buf_clk cell_7611 ( .C ( clk ), .D ( signal_22303 ), .Q ( signal_22304 ) ) ;
    buf_clk cell_7617 ( .C ( clk ), .D ( signal_22309 ), .Q ( signal_22310 ) ) ;
    buf_clk cell_7623 ( .C ( clk ), .D ( signal_22315 ), .Q ( signal_22316 ) ) ;
    buf_clk cell_7629 ( .C ( clk ), .D ( signal_22321 ), .Q ( signal_22322 ) ) ;
    buf_clk cell_7635 ( .C ( clk ), .D ( signal_22327 ), .Q ( signal_22328 ) ) ;
    buf_clk cell_7641 ( .C ( clk ), .D ( signal_22333 ), .Q ( signal_22334 ) ) ;
    buf_clk cell_7647 ( .C ( clk ), .D ( signal_22339 ), .Q ( signal_22340 ) ) ;
    buf_clk cell_7653 ( .C ( clk ), .D ( signal_22345 ), .Q ( signal_22346 ) ) ;
    buf_clk cell_7661 ( .C ( clk ), .D ( signal_22353 ), .Q ( signal_22354 ) ) ;
    buf_clk cell_7669 ( .C ( clk ), .D ( signal_22361 ), .Q ( signal_22362 ) ) ;
    buf_clk cell_7677 ( .C ( clk ), .D ( signal_22369 ), .Q ( signal_22370 ) ) ;
    buf_clk cell_7685 ( .C ( clk ), .D ( signal_22377 ), .Q ( signal_22378 ) ) ;
    buf_clk cell_7693 ( .C ( clk ), .D ( signal_22385 ), .Q ( signal_22386 ) ) ;
    buf_clk cell_7703 ( .C ( clk ), .D ( signal_22395 ), .Q ( signal_22396 ) ) ;
    buf_clk cell_7713 ( .C ( clk ), .D ( signal_22405 ), .Q ( signal_22406 ) ) ;
    buf_clk cell_7723 ( .C ( clk ), .D ( signal_22415 ), .Q ( signal_22416 ) ) ;
    buf_clk cell_7733 ( .C ( clk ), .D ( signal_22425 ), .Q ( signal_22426 ) ) ;
    buf_clk cell_7743 ( .C ( clk ), .D ( signal_22435 ), .Q ( signal_22436 ) ) ;
    buf_clk cell_7745 ( .C ( clk ), .D ( signal_2258 ), .Q ( signal_22438 ) ) ;
    buf_clk cell_7747 ( .C ( clk ), .D ( signal_7688 ), .Q ( signal_22440 ) ) ;
    buf_clk cell_7749 ( .C ( clk ), .D ( signal_7689 ), .Q ( signal_22442 ) ) ;
    buf_clk cell_7751 ( .C ( clk ), .D ( signal_7690 ), .Q ( signal_22444 ) ) ;
    buf_clk cell_7753 ( .C ( clk ), .D ( signal_7691 ), .Q ( signal_22446 ) ) ;
    buf_clk cell_7759 ( .C ( clk ), .D ( signal_22451 ), .Q ( signal_22452 ) ) ;
    buf_clk cell_7765 ( .C ( clk ), .D ( signal_22457 ), .Q ( signal_22458 ) ) ;
    buf_clk cell_7771 ( .C ( clk ), .D ( signal_22463 ), .Q ( signal_22464 ) ) ;
    buf_clk cell_7777 ( .C ( clk ), .D ( signal_22469 ), .Q ( signal_22470 ) ) ;
    buf_clk cell_7783 ( .C ( clk ), .D ( signal_22475 ), .Q ( signal_22476 ) ) ;
    buf_clk cell_7791 ( .C ( clk ), .D ( signal_22483 ), .Q ( signal_22484 ) ) ;
    buf_clk cell_7799 ( .C ( clk ), .D ( signal_22491 ), .Q ( signal_22492 ) ) ;
    buf_clk cell_7807 ( .C ( clk ), .D ( signal_22499 ), .Q ( signal_22500 ) ) ;
    buf_clk cell_7815 ( .C ( clk ), .D ( signal_22507 ), .Q ( signal_22508 ) ) ;
    buf_clk cell_7823 ( .C ( clk ), .D ( signal_22515 ), .Q ( signal_22516 ) ) ;
    buf_clk cell_7833 ( .C ( clk ), .D ( signal_22525 ), .Q ( signal_22526 ) ) ;
    buf_clk cell_7843 ( .C ( clk ), .D ( signal_22535 ), .Q ( signal_22536 ) ) ;
    buf_clk cell_7853 ( .C ( clk ), .D ( signal_22545 ), .Q ( signal_22546 ) ) ;
    buf_clk cell_7863 ( .C ( clk ), .D ( signal_22555 ), .Q ( signal_22556 ) ) ;
    buf_clk cell_7873 ( .C ( clk ), .D ( signal_22565 ), .Q ( signal_22566 ) ) ;
    buf_clk cell_7881 ( .C ( clk ), .D ( signal_22573 ), .Q ( signal_22574 ) ) ;
    buf_clk cell_7889 ( .C ( clk ), .D ( signal_22581 ), .Q ( signal_22582 ) ) ;
    buf_clk cell_7897 ( .C ( clk ), .D ( signal_22589 ), .Q ( signal_22590 ) ) ;
    buf_clk cell_7905 ( .C ( clk ), .D ( signal_22597 ), .Q ( signal_22598 ) ) ;
    buf_clk cell_7913 ( .C ( clk ), .D ( signal_22605 ), .Q ( signal_22606 ) ) ;
    buf_clk cell_7919 ( .C ( clk ), .D ( signal_22611 ), .Q ( signal_22612 ) ) ;
    buf_clk cell_7925 ( .C ( clk ), .D ( signal_22617 ), .Q ( signal_22618 ) ) ;
    buf_clk cell_7931 ( .C ( clk ), .D ( signal_22623 ), .Q ( signal_22624 ) ) ;
    buf_clk cell_7937 ( .C ( clk ), .D ( signal_22629 ), .Q ( signal_22630 ) ) ;
    buf_clk cell_7943 ( .C ( clk ), .D ( signal_22635 ), .Q ( signal_22636 ) ) ;
    buf_clk cell_7949 ( .C ( clk ), .D ( signal_22641 ), .Q ( signal_22642 ) ) ;
    buf_clk cell_7955 ( .C ( clk ), .D ( signal_22647 ), .Q ( signal_22648 ) ) ;
    buf_clk cell_7961 ( .C ( clk ), .D ( signal_22653 ), .Q ( signal_22654 ) ) ;
    buf_clk cell_7967 ( .C ( clk ), .D ( signal_22659 ), .Q ( signal_22660 ) ) ;
    buf_clk cell_7973 ( .C ( clk ), .D ( signal_22665 ), .Q ( signal_22666 ) ) ;
    buf_clk cell_7975 ( .C ( clk ), .D ( signal_21639 ), .Q ( signal_22668 ) ) ;
    buf_clk cell_7977 ( .C ( clk ), .D ( signal_21641 ), .Q ( signal_22670 ) ) ;
    buf_clk cell_7979 ( .C ( clk ), .D ( signal_21643 ), .Q ( signal_22672 ) ) ;
    buf_clk cell_7981 ( .C ( clk ), .D ( signal_21645 ), .Q ( signal_22674 ) ) ;
    buf_clk cell_7983 ( .C ( clk ), .D ( signal_21647 ), .Q ( signal_22676 ) ) ;
    buf_clk cell_7987 ( .C ( clk ), .D ( signal_22679 ), .Q ( signal_22680 ) ) ;
    buf_clk cell_7991 ( .C ( clk ), .D ( signal_22683 ), .Q ( signal_22684 ) ) ;
    buf_clk cell_7995 ( .C ( clk ), .D ( signal_22687 ), .Q ( signal_22688 ) ) ;
    buf_clk cell_7999 ( .C ( clk ), .D ( signal_22691 ), .Q ( signal_22692 ) ) ;
    buf_clk cell_8003 ( .C ( clk ), .D ( signal_22695 ), .Q ( signal_22696 ) ) ;
    buf_clk cell_8007 ( .C ( clk ), .D ( signal_22699 ), .Q ( signal_22700 ) ) ;
    buf_clk cell_8011 ( .C ( clk ), .D ( signal_22703 ), .Q ( signal_22704 ) ) ;
    buf_clk cell_8015 ( .C ( clk ), .D ( signal_22707 ), .Q ( signal_22708 ) ) ;
    buf_clk cell_8019 ( .C ( clk ), .D ( signal_22711 ), .Q ( signal_22712 ) ) ;
    buf_clk cell_8023 ( .C ( clk ), .D ( signal_22715 ), .Q ( signal_22716 ) ) ;
    buf_clk cell_8029 ( .C ( clk ), .D ( signal_22721 ), .Q ( signal_22722 ) ) ;
    buf_clk cell_8035 ( .C ( clk ), .D ( signal_22727 ), .Q ( signal_22728 ) ) ;
    buf_clk cell_8041 ( .C ( clk ), .D ( signal_22733 ), .Q ( signal_22734 ) ) ;
    buf_clk cell_8047 ( .C ( clk ), .D ( signal_22739 ), .Q ( signal_22740 ) ) ;
    buf_clk cell_8053 ( .C ( clk ), .D ( signal_22745 ), .Q ( signal_22746 ) ) ;
    buf_clk cell_8055 ( .C ( clk ), .D ( signal_2287 ), .Q ( signal_22748 ) ) ;
    buf_clk cell_8057 ( .C ( clk ), .D ( signal_7804 ), .Q ( signal_22750 ) ) ;
    buf_clk cell_8059 ( .C ( clk ), .D ( signal_7805 ), .Q ( signal_22752 ) ) ;
    buf_clk cell_8061 ( .C ( clk ), .D ( signal_7806 ), .Q ( signal_22754 ) ) ;
    buf_clk cell_8063 ( .C ( clk ), .D ( signal_7807 ), .Q ( signal_22756 ) ) ;
    buf_clk cell_8069 ( .C ( clk ), .D ( signal_22761 ), .Q ( signal_22762 ) ) ;
    buf_clk cell_8075 ( .C ( clk ), .D ( signal_22767 ), .Q ( signal_22768 ) ) ;
    buf_clk cell_8081 ( .C ( clk ), .D ( signal_22773 ), .Q ( signal_22774 ) ) ;
    buf_clk cell_8087 ( .C ( clk ), .D ( signal_22779 ), .Q ( signal_22780 ) ) ;
    buf_clk cell_8093 ( .C ( clk ), .D ( signal_22785 ), .Q ( signal_22786 ) ) ;
    buf_clk cell_8097 ( .C ( clk ), .D ( signal_22789 ), .Q ( signal_22790 ) ) ;
    buf_clk cell_8101 ( .C ( clk ), .D ( signal_22793 ), .Q ( signal_22794 ) ) ;
    buf_clk cell_8105 ( .C ( clk ), .D ( signal_22797 ), .Q ( signal_22798 ) ) ;
    buf_clk cell_8109 ( .C ( clk ), .D ( signal_22801 ), .Q ( signal_22802 ) ) ;
    buf_clk cell_8113 ( .C ( clk ), .D ( signal_22805 ), .Q ( signal_22806 ) ) ;
    buf_clk cell_8119 ( .C ( clk ), .D ( signal_22811 ), .Q ( signal_22812 ) ) ;
    buf_clk cell_8125 ( .C ( clk ), .D ( signal_22817 ), .Q ( signal_22818 ) ) ;
    buf_clk cell_8131 ( .C ( clk ), .D ( signal_22823 ), .Q ( signal_22824 ) ) ;
    buf_clk cell_8137 ( .C ( clk ), .D ( signal_22829 ), .Q ( signal_22830 ) ) ;
    buf_clk cell_8143 ( .C ( clk ), .D ( signal_22835 ), .Q ( signal_22836 ) ) ;
    buf_clk cell_8145 ( .C ( clk ), .D ( signal_2312 ), .Q ( signal_22838 ) ) ;
    buf_clk cell_8147 ( .C ( clk ), .D ( signal_7904 ), .Q ( signal_22840 ) ) ;
    buf_clk cell_8149 ( .C ( clk ), .D ( signal_7905 ), .Q ( signal_22842 ) ) ;
    buf_clk cell_8151 ( .C ( clk ), .D ( signal_7906 ), .Q ( signal_22844 ) ) ;
    buf_clk cell_8153 ( .C ( clk ), .D ( signal_7907 ), .Q ( signal_22846 ) ) ;
    buf_clk cell_8157 ( .C ( clk ), .D ( signal_22849 ), .Q ( signal_22850 ) ) ;
    buf_clk cell_8161 ( .C ( clk ), .D ( signal_22853 ), .Q ( signal_22854 ) ) ;
    buf_clk cell_8165 ( .C ( clk ), .D ( signal_22857 ), .Q ( signal_22858 ) ) ;
    buf_clk cell_8169 ( .C ( clk ), .D ( signal_22861 ), .Q ( signal_22862 ) ) ;
    buf_clk cell_8173 ( .C ( clk ), .D ( signal_22865 ), .Q ( signal_22866 ) ) ;
    buf_clk cell_8177 ( .C ( clk ), .D ( signal_22869 ), .Q ( signal_22870 ) ) ;
    buf_clk cell_8183 ( .C ( clk ), .D ( signal_22875 ), .Q ( signal_22876 ) ) ;
    buf_clk cell_8189 ( .C ( clk ), .D ( signal_22881 ), .Q ( signal_22882 ) ) ;
    buf_clk cell_8195 ( .C ( clk ), .D ( signal_22887 ), .Q ( signal_22888 ) ) ;
    buf_clk cell_8201 ( .C ( clk ), .D ( signal_22893 ), .Q ( signal_22894 ) ) ;
    buf_clk cell_8209 ( .C ( clk ), .D ( signal_22901 ), .Q ( signal_22902 ) ) ;
    buf_clk cell_8217 ( .C ( clk ), .D ( signal_22909 ), .Q ( signal_22910 ) ) ;
    buf_clk cell_8225 ( .C ( clk ), .D ( signal_22917 ), .Q ( signal_22918 ) ) ;
    buf_clk cell_8233 ( .C ( clk ), .D ( signal_22925 ), .Q ( signal_22926 ) ) ;
    buf_clk cell_8241 ( .C ( clk ), .D ( signal_22933 ), .Q ( signal_22934 ) ) ;
    buf_clk cell_8247 ( .C ( clk ), .D ( signal_22939 ), .Q ( signal_22940 ) ) ;
    buf_clk cell_8253 ( .C ( clk ), .D ( signal_22945 ), .Q ( signal_22946 ) ) ;
    buf_clk cell_8259 ( .C ( clk ), .D ( signal_22951 ), .Q ( signal_22952 ) ) ;
    buf_clk cell_8265 ( .C ( clk ), .D ( signal_22957 ), .Q ( signal_22958 ) ) ;
    buf_clk cell_8271 ( .C ( clk ), .D ( signal_22963 ), .Q ( signal_22964 ) ) ;
    buf_clk cell_8281 ( .C ( clk ), .D ( signal_22973 ), .Q ( signal_22974 ) ) ;
    buf_clk cell_8291 ( .C ( clk ), .D ( signal_22983 ), .Q ( signal_22984 ) ) ;
    buf_clk cell_8301 ( .C ( clk ), .D ( signal_22993 ), .Q ( signal_22994 ) ) ;
    buf_clk cell_8311 ( .C ( clk ), .D ( signal_23003 ), .Q ( signal_23004 ) ) ;
    buf_clk cell_8321 ( .C ( clk ), .D ( signal_23013 ), .Q ( signal_23014 ) ) ;
    buf_clk cell_8327 ( .C ( clk ), .D ( signal_23019 ), .Q ( signal_23020 ) ) ;
    buf_clk cell_8333 ( .C ( clk ), .D ( signal_23025 ), .Q ( signal_23026 ) ) ;
    buf_clk cell_8339 ( .C ( clk ), .D ( signal_23031 ), .Q ( signal_23032 ) ) ;
    buf_clk cell_8345 ( .C ( clk ), .D ( signal_23037 ), .Q ( signal_23038 ) ) ;
    buf_clk cell_8351 ( .C ( clk ), .D ( signal_23043 ), .Q ( signal_23044 ) ) ;
    buf_clk cell_8355 ( .C ( clk ), .D ( signal_2288 ), .Q ( signal_23048 ) ) ;
    buf_clk cell_8359 ( .C ( clk ), .D ( signal_7808 ), .Q ( signal_23052 ) ) ;
    buf_clk cell_8363 ( .C ( clk ), .D ( signal_7809 ), .Q ( signal_23056 ) ) ;
    buf_clk cell_8367 ( .C ( clk ), .D ( signal_7810 ), .Q ( signal_23060 ) ) ;
    buf_clk cell_8371 ( .C ( clk ), .D ( signal_7811 ), .Q ( signal_23064 ) ) ;
    buf_clk cell_8379 ( .C ( clk ), .D ( signal_23071 ), .Q ( signal_23072 ) ) ;
    buf_clk cell_8387 ( .C ( clk ), .D ( signal_23079 ), .Q ( signal_23080 ) ) ;
    buf_clk cell_8395 ( .C ( clk ), .D ( signal_23087 ), .Q ( signal_23088 ) ) ;
    buf_clk cell_8403 ( .C ( clk ), .D ( signal_23095 ), .Q ( signal_23096 ) ) ;
    buf_clk cell_8411 ( .C ( clk ), .D ( signal_23103 ), .Q ( signal_23104 ) ) ;
    buf_clk cell_8417 ( .C ( clk ), .D ( signal_23109 ), .Q ( signal_23110 ) ) ;
    buf_clk cell_8423 ( .C ( clk ), .D ( signal_23115 ), .Q ( signal_23116 ) ) ;
    buf_clk cell_8429 ( .C ( clk ), .D ( signal_23121 ), .Q ( signal_23122 ) ) ;
    buf_clk cell_8435 ( .C ( clk ), .D ( signal_23127 ), .Q ( signal_23128 ) ) ;
    buf_clk cell_8441 ( .C ( clk ), .D ( signal_23133 ), .Q ( signal_23134 ) ) ;
    buf_clk cell_8449 ( .C ( clk ), .D ( signal_23141 ), .Q ( signal_23142 ) ) ;
    buf_clk cell_8457 ( .C ( clk ), .D ( signal_23149 ), .Q ( signal_23150 ) ) ;
    buf_clk cell_8465 ( .C ( clk ), .D ( signal_23157 ), .Q ( signal_23158 ) ) ;
    buf_clk cell_8473 ( .C ( clk ), .D ( signal_23165 ), .Q ( signal_23166 ) ) ;
    buf_clk cell_8481 ( .C ( clk ), .D ( signal_23173 ), .Q ( signal_23174 ) ) ;
    buf_clk cell_8487 ( .C ( clk ), .D ( signal_23179 ), .Q ( signal_23180 ) ) ;
    buf_clk cell_8493 ( .C ( clk ), .D ( signal_23185 ), .Q ( signal_23186 ) ) ;
    buf_clk cell_8499 ( .C ( clk ), .D ( signal_23191 ), .Q ( signal_23192 ) ) ;
    buf_clk cell_8505 ( .C ( clk ), .D ( signal_23197 ), .Q ( signal_23198 ) ) ;
    buf_clk cell_8511 ( .C ( clk ), .D ( signal_23203 ), .Q ( signal_23204 ) ) ;
    buf_clk cell_8519 ( .C ( clk ), .D ( signal_23211 ), .Q ( signal_23212 ) ) ;
    buf_clk cell_8527 ( .C ( clk ), .D ( signal_23219 ), .Q ( signal_23220 ) ) ;
    buf_clk cell_8535 ( .C ( clk ), .D ( signal_23227 ), .Q ( signal_23228 ) ) ;
    buf_clk cell_8543 ( .C ( clk ), .D ( signal_23235 ), .Q ( signal_23236 ) ) ;
    buf_clk cell_8551 ( .C ( clk ), .D ( signal_23243 ), .Q ( signal_23244 ) ) ;
    buf_clk cell_8555 ( .C ( clk ), .D ( signal_2213 ), .Q ( signal_23248 ) ) ;
    buf_clk cell_8559 ( .C ( clk ), .D ( signal_7508 ), .Q ( signal_23252 ) ) ;
    buf_clk cell_8563 ( .C ( clk ), .D ( signal_7509 ), .Q ( signal_23256 ) ) ;
    buf_clk cell_8567 ( .C ( clk ), .D ( signal_7510 ), .Q ( signal_23260 ) ) ;
    buf_clk cell_8571 ( .C ( clk ), .D ( signal_7511 ), .Q ( signal_23264 ) ) ;
    buf_clk cell_8577 ( .C ( clk ), .D ( signal_23269 ), .Q ( signal_23270 ) ) ;
    buf_clk cell_8583 ( .C ( clk ), .D ( signal_23275 ), .Q ( signal_23276 ) ) ;
    buf_clk cell_8589 ( .C ( clk ), .D ( signal_23281 ), .Q ( signal_23282 ) ) ;
    buf_clk cell_8595 ( .C ( clk ), .D ( signal_23287 ), .Q ( signal_23288 ) ) ;
    buf_clk cell_8601 ( .C ( clk ), .D ( signal_23293 ), .Q ( signal_23294 ) ) ;
    buf_clk cell_8607 ( .C ( clk ), .D ( signal_23299 ), .Q ( signal_23300 ) ) ;
    buf_clk cell_8613 ( .C ( clk ), .D ( signal_23305 ), .Q ( signal_23306 ) ) ;
    buf_clk cell_8619 ( .C ( clk ), .D ( signal_23311 ), .Q ( signal_23312 ) ) ;
    buf_clk cell_8625 ( .C ( clk ), .D ( signal_23317 ), .Q ( signal_23318 ) ) ;
    buf_clk cell_8631 ( .C ( clk ), .D ( signal_23323 ), .Q ( signal_23324 ) ) ;
    buf_clk cell_8635 ( .C ( clk ), .D ( signal_2189 ), .Q ( signal_23328 ) ) ;
    buf_clk cell_8639 ( .C ( clk ), .D ( signal_7412 ), .Q ( signal_23332 ) ) ;
    buf_clk cell_8643 ( .C ( clk ), .D ( signal_7413 ), .Q ( signal_23336 ) ) ;
    buf_clk cell_8647 ( .C ( clk ), .D ( signal_7414 ), .Q ( signal_23340 ) ) ;
    buf_clk cell_8651 ( .C ( clk ), .D ( signal_7415 ), .Q ( signal_23344 ) ) ;
    buf_clk cell_8655 ( .C ( clk ), .D ( signal_2138 ), .Q ( signal_23348 ) ) ;
    buf_clk cell_8659 ( .C ( clk ), .D ( signal_7208 ), .Q ( signal_23352 ) ) ;
    buf_clk cell_8663 ( .C ( clk ), .D ( signal_7209 ), .Q ( signal_23356 ) ) ;
    buf_clk cell_8667 ( .C ( clk ), .D ( signal_7210 ), .Q ( signal_23360 ) ) ;
    buf_clk cell_8671 ( .C ( clk ), .D ( signal_7211 ), .Q ( signal_23364 ) ) ;
    buf_clk cell_8677 ( .C ( clk ), .D ( signal_23369 ), .Q ( signal_23370 ) ) ;
    buf_clk cell_8685 ( .C ( clk ), .D ( signal_23377 ), .Q ( signal_23378 ) ) ;
    buf_clk cell_8693 ( .C ( clk ), .D ( signal_23385 ), .Q ( signal_23386 ) ) ;
    buf_clk cell_8701 ( .C ( clk ), .D ( signal_23393 ), .Q ( signal_23394 ) ) ;
    buf_clk cell_8709 ( .C ( clk ), .D ( signal_23401 ), .Q ( signal_23402 ) ) ;
    buf_clk cell_8721 ( .C ( clk ), .D ( signal_23413 ), .Q ( signal_23414 ) ) ;
    buf_clk cell_8733 ( .C ( clk ), .D ( signal_23425 ), .Q ( signal_23426 ) ) ;
    buf_clk cell_8745 ( .C ( clk ), .D ( signal_23437 ), .Q ( signal_23438 ) ) ;
    buf_clk cell_8757 ( .C ( clk ), .D ( signal_23449 ), .Q ( signal_23450 ) ) ;
    buf_clk cell_8769 ( .C ( clk ), .D ( signal_23461 ), .Q ( signal_23462 ) ) ;
    buf_clk cell_8775 ( .C ( clk ), .D ( signal_2238 ), .Q ( signal_23468 ) ) ;
    buf_clk cell_8781 ( .C ( clk ), .D ( signal_7608 ), .Q ( signal_23474 ) ) ;
    buf_clk cell_8787 ( .C ( clk ), .D ( signal_7609 ), .Q ( signal_23480 ) ) ;
    buf_clk cell_8793 ( .C ( clk ), .D ( signal_7610 ), .Q ( signal_23486 ) ) ;
    buf_clk cell_8799 ( .C ( clk ), .D ( signal_7611 ), .Q ( signal_23492 ) ) ;
    buf_clk cell_8805 ( .C ( clk ), .D ( signal_2210 ), .Q ( signal_23498 ) ) ;
    buf_clk cell_8811 ( .C ( clk ), .D ( signal_7496 ), .Q ( signal_23504 ) ) ;
    buf_clk cell_8817 ( .C ( clk ), .D ( signal_7497 ), .Q ( signal_23510 ) ) ;
    buf_clk cell_8823 ( .C ( clk ), .D ( signal_7498 ), .Q ( signal_23516 ) ) ;
    buf_clk cell_8829 ( .C ( clk ), .D ( signal_7499 ), .Q ( signal_23522 ) ) ;
    buf_clk cell_8843 ( .C ( clk ), .D ( signal_23535 ), .Q ( signal_23536 ) ) ;
    buf_clk cell_8857 ( .C ( clk ), .D ( signal_23549 ), .Q ( signal_23550 ) ) ;
    buf_clk cell_8871 ( .C ( clk ), .D ( signal_23563 ), .Q ( signal_23564 ) ) ;
    buf_clk cell_8885 ( .C ( clk ), .D ( signal_23577 ), .Q ( signal_23578 ) ) ;
    buf_clk cell_8899 ( .C ( clk ), .D ( signal_23591 ), .Q ( signal_23592 ) ) ;
    buf_clk cell_8907 ( .C ( clk ), .D ( signal_23599 ), .Q ( signal_23600 ) ) ;
    buf_clk cell_8915 ( .C ( clk ), .D ( signal_23607 ), .Q ( signal_23608 ) ) ;
    buf_clk cell_8923 ( .C ( clk ), .D ( signal_23615 ), .Q ( signal_23616 ) ) ;
    buf_clk cell_8931 ( .C ( clk ), .D ( signal_23623 ), .Q ( signal_23624 ) ) ;
    buf_clk cell_8939 ( .C ( clk ), .D ( signal_23631 ), .Q ( signal_23632 ) ) ;
    buf_clk cell_8953 ( .C ( clk ), .D ( signal_23645 ), .Q ( signal_23646 ) ) ;
    buf_clk cell_8967 ( .C ( clk ), .D ( signal_23659 ), .Q ( signal_23660 ) ) ;
    buf_clk cell_8981 ( .C ( clk ), .D ( signal_23673 ), .Q ( signal_23674 ) ) ;
    buf_clk cell_8995 ( .C ( clk ), .D ( signal_23687 ), .Q ( signal_23688 ) ) ;
    buf_clk cell_9009 ( .C ( clk ), .D ( signal_23701 ), .Q ( signal_23702 ) ) ;
    buf_clk cell_9017 ( .C ( clk ), .D ( signal_23709 ), .Q ( signal_23710 ) ) ;
    buf_clk cell_9025 ( .C ( clk ), .D ( signal_23717 ), .Q ( signal_23718 ) ) ;
    buf_clk cell_9033 ( .C ( clk ), .D ( signal_23725 ), .Q ( signal_23726 ) ) ;
    buf_clk cell_9041 ( .C ( clk ), .D ( signal_23733 ), .Q ( signal_23734 ) ) ;
    buf_clk cell_9049 ( .C ( clk ), .D ( signal_23741 ), .Q ( signal_23742 ) ) ;
    buf_clk cell_9077 ( .C ( clk ), .D ( signal_23769 ), .Q ( signal_23770 ) ) ;
    buf_clk cell_9087 ( .C ( clk ), .D ( signal_23779 ), .Q ( signal_23780 ) ) ;
    buf_clk cell_9097 ( .C ( clk ), .D ( signal_23789 ), .Q ( signal_23790 ) ) ;
    buf_clk cell_9107 ( .C ( clk ), .D ( signal_23799 ), .Q ( signal_23800 ) ) ;
    buf_clk cell_9117 ( .C ( clk ), .D ( signal_23809 ), .Q ( signal_23810 ) ) ;
    buf_clk cell_9153 ( .C ( clk ), .D ( signal_23845 ), .Q ( signal_23846 ) ) ;
    buf_clk cell_9169 ( .C ( clk ), .D ( signal_23861 ), .Q ( signal_23862 ) ) ;
    buf_clk cell_9185 ( .C ( clk ), .D ( signal_23877 ), .Q ( signal_23878 ) ) ;
    buf_clk cell_9201 ( .C ( clk ), .D ( signal_23893 ), .Q ( signal_23894 ) ) ;
    buf_clk cell_9217 ( .C ( clk ), .D ( signal_23909 ), .Q ( signal_23910 ) ) ;
    buf_clk cell_9253 ( .C ( clk ), .D ( signal_23945 ), .Q ( signal_23946 ) ) ;
    buf_clk cell_9269 ( .C ( clk ), .D ( signal_23961 ), .Q ( signal_23962 ) ) ;
    buf_clk cell_9285 ( .C ( clk ), .D ( signal_23977 ), .Q ( signal_23978 ) ) ;
    buf_clk cell_9301 ( .C ( clk ), .D ( signal_23993 ), .Q ( signal_23994 ) ) ;
    buf_clk cell_9317 ( .C ( clk ), .D ( signal_24009 ), .Q ( signal_24010 ) ) ;
    buf_clk cell_9327 ( .C ( clk ), .D ( signal_24019 ), .Q ( signal_24020 ) ) ;
    buf_clk cell_9337 ( .C ( clk ), .D ( signal_24029 ), .Q ( signal_24030 ) ) ;
    buf_clk cell_9347 ( .C ( clk ), .D ( signal_24039 ), .Q ( signal_24040 ) ) ;
    buf_clk cell_9357 ( .C ( clk ), .D ( signal_24049 ), .Q ( signal_24050 ) ) ;
    buf_clk cell_9367 ( .C ( clk ), .D ( signal_24059 ), .Q ( signal_24060 ) ) ;
    buf_clk cell_9425 ( .C ( clk ), .D ( signal_2289 ), .Q ( signal_24118 ) ) ;
    buf_clk cell_9435 ( .C ( clk ), .D ( signal_7812 ), .Q ( signal_24128 ) ) ;
    buf_clk cell_9445 ( .C ( clk ), .D ( signal_7813 ), .Q ( signal_24138 ) ) ;
    buf_clk cell_9455 ( .C ( clk ), .D ( signal_7814 ), .Q ( signal_24148 ) ) ;
    buf_clk cell_9465 ( .C ( clk ), .D ( signal_7815 ), .Q ( signal_24158 ) ) ;
    buf_clk cell_9505 ( .C ( clk ), .D ( signal_2265 ), .Q ( signal_24198 ) ) ;
    buf_clk cell_9515 ( .C ( clk ), .D ( signal_7716 ), .Q ( signal_24208 ) ) ;
    buf_clk cell_9525 ( .C ( clk ), .D ( signal_7717 ), .Q ( signal_24218 ) ) ;
    buf_clk cell_9535 ( .C ( clk ), .D ( signal_7718 ), .Q ( signal_24228 ) ) ;
    buf_clk cell_9545 ( .C ( clk ), .D ( signal_7719 ), .Q ( signal_24238 ) ) ;
    buf_clk cell_9561 ( .C ( clk ), .D ( signal_24253 ), .Q ( signal_24254 ) ) ;
    buf_clk cell_9577 ( .C ( clk ), .D ( signal_24269 ), .Q ( signal_24270 ) ) ;
    buf_clk cell_9593 ( .C ( clk ), .D ( signal_24285 ), .Q ( signal_24286 ) ) ;
    buf_clk cell_9609 ( .C ( clk ), .D ( signal_24301 ), .Q ( signal_24302 ) ) ;
    buf_clk cell_9625 ( .C ( clk ), .D ( signal_24317 ), .Q ( signal_24318 ) ) ;
    buf_clk cell_9643 ( .C ( clk ), .D ( signal_24335 ), .Q ( signal_24336 ) ) ;
    buf_clk cell_9661 ( .C ( clk ), .D ( signal_24353 ), .Q ( signal_24354 ) ) ;
    buf_clk cell_9679 ( .C ( clk ), .D ( signal_24371 ), .Q ( signal_24372 ) ) ;
    buf_clk cell_9697 ( .C ( clk ), .D ( signal_24389 ), .Q ( signal_24390 ) ) ;
    buf_clk cell_9715 ( .C ( clk ), .D ( signal_24407 ), .Q ( signal_24408 ) ) ;
    buf_clk cell_9893 ( .C ( clk ), .D ( signal_24585 ), .Q ( signal_24586 ) ) ;
    buf_clk cell_9913 ( .C ( clk ), .D ( signal_24605 ), .Q ( signal_24606 ) ) ;
    buf_clk cell_9933 ( .C ( clk ), .D ( signal_24625 ), .Q ( signal_24626 ) ) ;
    buf_clk cell_9953 ( .C ( clk ), .D ( signal_24645 ), .Q ( signal_24646 ) ) ;
    buf_clk cell_9973 ( .C ( clk ), .D ( signal_24665 ), .Q ( signal_24666 ) ) ;

    /* cells in depth 16 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2180 ( .a ({signal_21487, signal_21477, signal_21467, signal_21457, signal_21447}), .b ({signal_7183, signal_7182, signal_7181, signal_7180, signal_2131}), .clk ( clk ), .r ({Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720]}), .c ({signal_7439, signal_7438, signal_7437, signal_7436, signal_2195}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2181 ( .a ({signal_21517, signal_21511, signal_21505, signal_21499, signal_21493}), .b ({signal_7191, signal_7190, signal_7189, signal_7188, signal_2133}), .clk ( clk ), .r ({Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730]}), .c ({signal_7443, signal_7442, signal_7441, signal_7440, signal_2196}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2182 ( .a ({signal_21557, signal_21549, signal_21541, signal_21533, signal_21525}), .b ({signal_7203, signal_7202, signal_7201, signal_7200, signal_2136}), .clk ( clk ), .r ({Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740]}), .c ({signal_7447, signal_7446, signal_7445, signal_7444, signal_2197}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2183 ( .a ({signal_21597, signal_21589, signal_21581, signal_21573, signal_21565}), .b ({signal_7207, signal_7206, signal_7205, signal_7204, signal_2137}), .clk ( clk ), .r ({Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750]}), .c ({signal_7451, signal_7450, signal_7449, signal_7448, signal_2198}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2199 ( .a ({signal_7439, signal_7438, signal_7437, signal_7436, signal_2195}), .b ({signal_7515, signal_7514, signal_7513, signal_7512, signal_2214}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2225 ( .a ({signal_21617, signal_21613, signal_21609, signal_21605, signal_21601}), .b ({signal_7399, signal_7398, signal_7397, signal_7396, signal_2185}), .clk ( clk ), .r ({Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760]}), .c ({signal_7619, signal_7618, signal_7617, signal_7616, signal_2240}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2226 ( .a ({signal_21637, signal_21633, signal_21629, signal_21625, signal_21621}), .b ({signal_7407, signal_7406, signal_7405, signal_7404, signal_2187}), .clk ( clk ), .r ({Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770]}), .c ({signal_7623, signal_7622, signal_7621, signal_7620, signal_2241}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2227 ( .a ({signal_21647, signal_21645, signal_21643, signal_21641, signal_21639}), .b ({signal_7279, signal_7278, signal_7277, signal_7276, signal_2155}), .clk ( clk ), .r ({Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780]}), .c ({signal_7627, signal_7626, signal_7625, signal_7624, signal_2242}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2228 ( .a ({signal_7427, signal_7426, signal_7425, signal_7424, signal_2192}), .b ({signal_21657, signal_21655, signal_21653, signal_21651, signal_21649}), .clk ( clk ), .r ({Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790]}), .c ({signal_7631, signal_7630, signal_7629, signal_7628, signal_2243}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2229 ( .a ({signal_21677, signal_21673, signal_21669, signal_21665, signal_21661}), .b ({signal_7435, signal_7434, signal_7433, signal_7432, signal_2194}), .clk ( clk ), .r ({Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800]}), .c ({signal_7635, signal_7634, signal_7633, signal_7632, signal_2244}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2244 ( .a ({signal_7619, signal_7618, signal_7617, signal_7616, signal_2240}), .b ({signal_7695, signal_7694, signal_7693, signal_7692, signal_2259}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2245 ( .a ({signal_7627, signal_7626, signal_7625, signal_7624, signal_2242}), .b ({signal_7699, signal_7698, signal_7697, signal_7696, signal_2260}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2246 ( .a ({signal_7635, signal_7634, signal_7633, signal_7632, signal_2244}), .b ({signal_7703, signal_7702, signal_7701, signal_7700, signal_2261}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2247 ( .a ({signal_21727, signal_21717, signal_21707, signal_21697, signal_21687}), .b ({signal_7519, signal_7518, signal_7517, signal_7516, signal_2215}), .clk ( clk ), .r ({Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810]}), .c ({signal_7707, signal_7706, signal_7705, signal_7704, signal_2262}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2255 ( .a ({signal_21757, signal_21751, signal_21745, signal_21739, signal_21733}), .b ({signal_7555, signal_7554, signal_7553, signal_7552, signal_2224}), .clk ( clk ), .r ({Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820]}), .c ({signal_7739, signal_7738, signal_7737, signal_7736, signal_2270}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2256 ( .a ({signal_21767, signal_21765, signal_21763, signal_21761, signal_21759}), .b ({signal_7559, signal_7558, signal_7557, signal_7556, signal_2225}), .clk ( clk ), .r ({Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830]}), .c ({signal_7743, signal_7742, signal_7741, signal_7740, signal_2271}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2257 ( .a ({signal_21807, signal_21799, signal_21791, signal_21783, signal_21775}), .b ({signal_7563, signal_7562, signal_7561, signal_7560, signal_2226}), .clk ( clk ), .r ({Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840]}), .c ({signal_7747, signal_7746, signal_7745, signal_7744, signal_2272}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2258 ( .a ({signal_21837, signal_21831, signal_21825, signal_21819, signal_21813}), .b ({signal_7567, signal_7566, signal_7565, signal_7564, signal_2227}), .clk ( clk ), .r ({Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850]}), .c ({signal_7751, signal_7750, signal_7749, signal_7748, signal_2273}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2259 ( .a ({signal_21877, signal_21869, signal_21861, signal_21853, signal_21845}), .b ({signal_7575, signal_7574, signal_7573, signal_7572, signal_2229}), .clk ( clk ), .r ({Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860]}), .c ({signal_7755, signal_7754, signal_7753, signal_7752, signal_2274}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2260 ( .a ({signal_21917, signal_21909, signal_21901, signal_21893, signal_21885}), .b ({signal_7579, signal_7578, signal_7577, signal_7576, signal_2230}), .clk ( clk ), .r ({Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870]}), .c ({signal_7759, signal_7758, signal_7757, signal_7756, signal_2275}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2261 ( .a ({signal_21957, signal_21949, signal_21941, signal_21933, signal_21925}), .b ({signal_7583, signal_7582, signal_7581, signal_7580, signal_2231}), .clk ( clk ), .r ({Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880]}), .c ({signal_7763, signal_7762, signal_7761, signal_7760, signal_2276}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2262 ( .a ({signal_21617, signal_21613, signal_21609, signal_21605, signal_21601}), .b ({signal_7503, signal_7502, signal_7501, signal_7500, signal_2211}), .clk ( clk ), .r ({Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890]}), .c ({signal_7767, signal_7766, signal_7765, signal_7764, signal_2277}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2263 ( .a ({signal_22007, signal_21997, signal_21987, signal_21977, signal_21967}), .b ({signal_7595, signal_7594, signal_7593, signal_7592, signal_2234}), .clk ( clk ), .r ({Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900]}), .c ({signal_7771, signal_7770, signal_7769, signal_7768, signal_2278}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2264 ( .a ({signal_7479, signal_7478, signal_7477, signal_7476, signal_2205}), .b ({signal_7599, signal_7598, signal_7597, signal_7596, signal_2235}), .clk ( clk ), .r ({Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910]}), .c ({signal_7775, signal_7774, signal_7773, signal_7772, signal_2279}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2265 ( .a ({signal_22047, signal_22039, signal_22031, signal_22023, signal_22015}), .b ({signal_7507, signal_7506, signal_7505, signal_7504, signal_2212}), .clk ( clk ), .r ({Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920]}), .c ({signal_7779, signal_7778, signal_7777, signal_7776, signal_2280}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2266 ( .a ({signal_22087, signal_22079, signal_22071, signal_22063, signal_22055}), .b ({signal_7607, signal_7606, signal_7605, signal_7604, signal_2237}), .clk ( clk ), .r ({Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930]}), .c ({signal_7783, signal_7782, signal_7781, signal_7780, signal_2281}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2275 ( .a ({signal_7743, signal_7742, signal_7741, signal_7740, signal_2271}), .b ({signal_7819, signal_7818, signal_7817, signal_7816, signal_2290}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2276 ( .a ({signal_7747, signal_7746, signal_7745, signal_7744, signal_2272}), .b ({signal_7823, signal_7822, signal_7821, signal_7820, signal_2291}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2277 ( .a ({signal_7755, signal_7754, signal_7753, signal_7752, signal_2274}), .b ({signal_7827, signal_7826, signal_7825, signal_7824, signal_2292}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2278 ( .a ({signal_7763, signal_7762, signal_7761, signal_7760, signal_2276}), .b ({signal_7831, signal_7830, signal_7829, signal_7828, signal_2293}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2279 ( .a ({signal_7767, signal_7766, signal_7765, signal_7764, signal_2277}), .b ({signal_7835, signal_7834, signal_7833, signal_7832, signal_2294}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2280 ( .a ({signal_7779, signal_7778, signal_7777, signal_7776, signal_2280}), .b ({signal_7839, signal_7838, signal_7837, signal_7836, signal_2295}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2287 ( .a ({signal_7715, signal_7714, signal_7713, signal_7712, signal_2264}), .b ({signal_7547, signal_7546, signal_7545, signal_7544, signal_2222}), .clk ( clk ), .r ({Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940]}), .c ({signal_7867, signal_7866, signal_7865, signal_7864, signal_2302}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2288 ( .a ({signal_22097, signal_22095, signal_22093, signal_22091, signal_22089}), .b ({signal_7675, signal_7674, signal_7673, signal_7672, signal_2254}), .clk ( clk ), .r ({Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950]}), .c ({signal_7871, signal_7870, signal_7869, signal_7868, signal_2303}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2290 ( .a ({signal_22097, signal_22095, signal_22093, signal_22091, signal_22089}), .b ({signal_7683, signal_7682, signal_7681, signal_7680, signal_2256}), .clk ( clk ), .r ({Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960]}), .c ({signal_7879, signal_7878, signal_7877, signal_7876, signal_2305}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2299 ( .a ({signal_7871, signal_7870, signal_7869, signal_7868, signal_2303}), .b ({signal_7915, signal_7914, signal_7913, signal_7912, signal_2314}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2301 ( .a ({signal_7879, signal_7878, signal_7877, signal_7876, signal_2305}), .b ({signal_7923, signal_7922, signal_7921, signal_7920, signal_2316}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2304 ( .a ({signal_22137, signal_22129, signal_22121, signal_22113, signal_22105}), .b ({signal_7847, signal_7846, signal_7845, signal_7844, signal_2297}), .clk ( clk ), .r ({Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970]}), .c ({signal_7935, signal_7934, signal_7933, signal_7932, signal_2319}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2305 ( .a ({signal_22177, signal_22169, signal_22161, signal_22153, signal_22145}), .b ({signal_7859, signal_7858, signal_7857, signal_7856, signal_2300}), .clk ( clk ), .r ({Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980]}), .c ({signal_7939, signal_7938, signal_7937, signal_7936, signal_2320}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2306 ( .a ({signal_22217, signal_22209, signal_22201, signal_22193, signal_22185}), .b ({signal_7863, signal_7862, signal_7861, signal_7860, signal_2301}), .clk ( clk ), .r ({Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990]}), .c ({signal_7943, signal_7942, signal_7941, signal_7940, signal_2321}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2307 ( .a ({signal_7803, signal_7802, signal_7801, signal_7800, signal_2286}), .b ({signal_7591, signal_7590, signal_7589, signal_7588, signal_2233}), .clk ( clk ), .r ({Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000]}), .c ({signal_7947, signal_7946, signal_7945, signal_7944, signal_2322}) ) ;
    buf_clk cell_7530 ( .C ( clk ), .D ( signal_22222 ), .Q ( signal_22223 ) ) ;
    buf_clk cell_7536 ( .C ( clk ), .D ( signal_22228 ), .Q ( signal_22229 ) ) ;
    buf_clk cell_7542 ( .C ( clk ), .D ( signal_22234 ), .Q ( signal_22235 ) ) ;
    buf_clk cell_7548 ( .C ( clk ), .D ( signal_22240 ), .Q ( signal_22241 ) ) ;
    buf_clk cell_7554 ( .C ( clk ), .D ( signal_22246 ), .Q ( signal_22247 ) ) ;
    buf_clk cell_7562 ( .C ( clk ), .D ( signal_22254 ), .Q ( signal_22255 ) ) ;
    buf_clk cell_7570 ( .C ( clk ), .D ( signal_22262 ), .Q ( signal_22263 ) ) ;
    buf_clk cell_7578 ( .C ( clk ), .D ( signal_22270 ), .Q ( signal_22271 ) ) ;
    buf_clk cell_7586 ( .C ( clk ), .D ( signal_22278 ), .Q ( signal_22279 ) ) ;
    buf_clk cell_7594 ( .C ( clk ), .D ( signal_22286 ), .Q ( signal_22287 ) ) ;
    buf_clk cell_7600 ( .C ( clk ), .D ( signal_22292 ), .Q ( signal_22293 ) ) ;
    buf_clk cell_7606 ( .C ( clk ), .D ( signal_22298 ), .Q ( signal_22299 ) ) ;
    buf_clk cell_7612 ( .C ( clk ), .D ( signal_22304 ), .Q ( signal_22305 ) ) ;
    buf_clk cell_7618 ( .C ( clk ), .D ( signal_22310 ), .Q ( signal_22311 ) ) ;
    buf_clk cell_7624 ( .C ( clk ), .D ( signal_22316 ), .Q ( signal_22317 ) ) ;
    buf_clk cell_7630 ( .C ( clk ), .D ( signal_22322 ), .Q ( signal_22323 ) ) ;
    buf_clk cell_7636 ( .C ( clk ), .D ( signal_22328 ), .Q ( signal_22329 ) ) ;
    buf_clk cell_7642 ( .C ( clk ), .D ( signal_22334 ), .Q ( signal_22335 ) ) ;
    buf_clk cell_7648 ( .C ( clk ), .D ( signal_22340 ), .Q ( signal_22341 ) ) ;
    buf_clk cell_7654 ( .C ( clk ), .D ( signal_22346 ), .Q ( signal_22347 ) ) ;
    buf_clk cell_7662 ( .C ( clk ), .D ( signal_22354 ), .Q ( signal_22355 ) ) ;
    buf_clk cell_7670 ( .C ( clk ), .D ( signal_22362 ), .Q ( signal_22363 ) ) ;
    buf_clk cell_7678 ( .C ( clk ), .D ( signal_22370 ), .Q ( signal_22371 ) ) ;
    buf_clk cell_7686 ( .C ( clk ), .D ( signal_22378 ), .Q ( signal_22379 ) ) ;
    buf_clk cell_7694 ( .C ( clk ), .D ( signal_22386 ), .Q ( signal_22387 ) ) ;
    buf_clk cell_7704 ( .C ( clk ), .D ( signal_22396 ), .Q ( signal_22397 ) ) ;
    buf_clk cell_7714 ( .C ( clk ), .D ( signal_22406 ), .Q ( signal_22407 ) ) ;
    buf_clk cell_7724 ( .C ( clk ), .D ( signal_22416 ), .Q ( signal_22417 ) ) ;
    buf_clk cell_7734 ( .C ( clk ), .D ( signal_22426 ), .Q ( signal_22427 ) ) ;
    buf_clk cell_7744 ( .C ( clk ), .D ( signal_22436 ), .Q ( signal_22437 ) ) ;
    buf_clk cell_7746 ( .C ( clk ), .D ( signal_22438 ), .Q ( signal_22439 ) ) ;
    buf_clk cell_7748 ( .C ( clk ), .D ( signal_22440 ), .Q ( signal_22441 ) ) ;
    buf_clk cell_7750 ( .C ( clk ), .D ( signal_22442 ), .Q ( signal_22443 ) ) ;
    buf_clk cell_7752 ( .C ( clk ), .D ( signal_22444 ), .Q ( signal_22445 ) ) ;
    buf_clk cell_7754 ( .C ( clk ), .D ( signal_22446 ), .Q ( signal_22447 ) ) ;
    buf_clk cell_7760 ( .C ( clk ), .D ( signal_22452 ), .Q ( signal_22453 ) ) ;
    buf_clk cell_7766 ( .C ( clk ), .D ( signal_22458 ), .Q ( signal_22459 ) ) ;
    buf_clk cell_7772 ( .C ( clk ), .D ( signal_22464 ), .Q ( signal_22465 ) ) ;
    buf_clk cell_7778 ( .C ( clk ), .D ( signal_22470 ), .Q ( signal_22471 ) ) ;
    buf_clk cell_7784 ( .C ( clk ), .D ( signal_22476 ), .Q ( signal_22477 ) ) ;
    buf_clk cell_7792 ( .C ( clk ), .D ( signal_22484 ), .Q ( signal_22485 ) ) ;
    buf_clk cell_7800 ( .C ( clk ), .D ( signal_22492 ), .Q ( signal_22493 ) ) ;
    buf_clk cell_7808 ( .C ( clk ), .D ( signal_22500 ), .Q ( signal_22501 ) ) ;
    buf_clk cell_7816 ( .C ( clk ), .D ( signal_22508 ), .Q ( signal_22509 ) ) ;
    buf_clk cell_7824 ( .C ( clk ), .D ( signal_22516 ), .Q ( signal_22517 ) ) ;
    buf_clk cell_7834 ( .C ( clk ), .D ( signal_22526 ), .Q ( signal_22527 ) ) ;
    buf_clk cell_7844 ( .C ( clk ), .D ( signal_22536 ), .Q ( signal_22537 ) ) ;
    buf_clk cell_7854 ( .C ( clk ), .D ( signal_22546 ), .Q ( signal_22547 ) ) ;
    buf_clk cell_7864 ( .C ( clk ), .D ( signal_22556 ), .Q ( signal_22557 ) ) ;
    buf_clk cell_7874 ( .C ( clk ), .D ( signal_22566 ), .Q ( signal_22567 ) ) ;
    buf_clk cell_7882 ( .C ( clk ), .D ( signal_22574 ), .Q ( signal_22575 ) ) ;
    buf_clk cell_7890 ( .C ( clk ), .D ( signal_22582 ), .Q ( signal_22583 ) ) ;
    buf_clk cell_7898 ( .C ( clk ), .D ( signal_22590 ), .Q ( signal_22591 ) ) ;
    buf_clk cell_7906 ( .C ( clk ), .D ( signal_22598 ), .Q ( signal_22599 ) ) ;
    buf_clk cell_7914 ( .C ( clk ), .D ( signal_22606 ), .Q ( signal_22607 ) ) ;
    buf_clk cell_7920 ( .C ( clk ), .D ( signal_22612 ), .Q ( signal_22613 ) ) ;
    buf_clk cell_7926 ( .C ( clk ), .D ( signal_22618 ), .Q ( signal_22619 ) ) ;
    buf_clk cell_7932 ( .C ( clk ), .D ( signal_22624 ), .Q ( signal_22625 ) ) ;
    buf_clk cell_7938 ( .C ( clk ), .D ( signal_22630 ), .Q ( signal_22631 ) ) ;
    buf_clk cell_7944 ( .C ( clk ), .D ( signal_22636 ), .Q ( signal_22637 ) ) ;
    buf_clk cell_7950 ( .C ( clk ), .D ( signal_22642 ), .Q ( signal_22643 ) ) ;
    buf_clk cell_7956 ( .C ( clk ), .D ( signal_22648 ), .Q ( signal_22649 ) ) ;
    buf_clk cell_7962 ( .C ( clk ), .D ( signal_22654 ), .Q ( signal_22655 ) ) ;
    buf_clk cell_7968 ( .C ( clk ), .D ( signal_22660 ), .Q ( signal_22661 ) ) ;
    buf_clk cell_7974 ( .C ( clk ), .D ( signal_22666 ), .Q ( signal_22667 ) ) ;
    buf_clk cell_7976 ( .C ( clk ), .D ( signal_22668 ), .Q ( signal_22669 ) ) ;
    buf_clk cell_7978 ( .C ( clk ), .D ( signal_22670 ), .Q ( signal_22671 ) ) ;
    buf_clk cell_7980 ( .C ( clk ), .D ( signal_22672 ), .Q ( signal_22673 ) ) ;
    buf_clk cell_7982 ( .C ( clk ), .D ( signal_22674 ), .Q ( signal_22675 ) ) ;
    buf_clk cell_7984 ( .C ( clk ), .D ( signal_22676 ), .Q ( signal_22677 ) ) ;
    buf_clk cell_7988 ( .C ( clk ), .D ( signal_22680 ), .Q ( signal_22681 ) ) ;
    buf_clk cell_7992 ( .C ( clk ), .D ( signal_22684 ), .Q ( signal_22685 ) ) ;
    buf_clk cell_7996 ( .C ( clk ), .D ( signal_22688 ), .Q ( signal_22689 ) ) ;
    buf_clk cell_8000 ( .C ( clk ), .D ( signal_22692 ), .Q ( signal_22693 ) ) ;
    buf_clk cell_8004 ( .C ( clk ), .D ( signal_22696 ), .Q ( signal_22697 ) ) ;
    buf_clk cell_8008 ( .C ( clk ), .D ( signal_22700 ), .Q ( signal_22701 ) ) ;
    buf_clk cell_8012 ( .C ( clk ), .D ( signal_22704 ), .Q ( signal_22705 ) ) ;
    buf_clk cell_8016 ( .C ( clk ), .D ( signal_22708 ), .Q ( signal_22709 ) ) ;
    buf_clk cell_8020 ( .C ( clk ), .D ( signal_22712 ), .Q ( signal_22713 ) ) ;
    buf_clk cell_8024 ( .C ( clk ), .D ( signal_22716 ), .Q ( signal_22717 ) ) ;
    buf_clk cell_8030 ( .C ( clk ), .D ( signal_22722 ), .Q ( signal_22723 ) ) ;
    buf_clk cell_8036 ( .C ( clk ), .D ( signal_22728 ), .Q ( signal_22729 ) ) ;
    buf_clk cell_8042 ( .C ( clk ), .D ( signal_22734 ), .Q ( signal_22735 ) ) ;
    buf_clk cell_8048 ( .C ( clk ), .D ( signal_22740 ), .Q ( signal_22741 ) ) ;
    buf_clk cell_8054 ( .C ( clk ), .D ( signal_22746 ), .Q ( signal_22747 ) ) ;
    buf_clk cell_8056 ( .C ( clk ), .D ( signal_22748 ), .Q ( signal_22749 ) ) ;
    buf_clk cell_8058 ( .C ( clk ), .D ( signal_22750 ), .Q ( signal_22751 ) ) ;
    buf_clk cell_8060 ( .C ( clk ), .D ( signal_22752 ), .Q ( signal_22753 ) ) ;
    buf_clk cell_8062 ( .C ( clk ), .D ( signal_22754 ), .Q ( signal_22755 ) ) ;
    buf_clk cell_8064 ( .C ( clk ), .D ( signal_22756 ), .Q ( signal_22757 ) ) ;
    buf_clk cell_8070 ( .C ( clk ), .D ( signal_22762 ), .Q ( signal_22763 ) ) ;
    buf_clk cell_8076 ( .C ( clk ), .D ( signal_22768 ), .Q ( signal_22769 ) ) ;
    buf_clk cell_8082 ( .C ( clk ), .D ( signal_22774 ), .Q ( signal_22775 ) ) ;
    buf_clk cell_8088 ( .C ( clk ), .D ( signal_22780 ), .Q ( signal_22781 ) ) ;
    buf_clk cell_8094 ( .C ( clk ), .D ( signal_22786 ), .Q ( signal_22787 ) ) ;
    buf_clk cell_8098 ( .C ( clk ), .D ( signal_22790 ), .Q ( signal_22791 ) ) ;
    buf_clk cell_8102 ( .C ( clk ), .D ( signal_22794 ), .Q ( signal_22795 ) ) ;
    buf_clk cell_8106 ( .C ( clk ), .D ( signal_22798 ), .Q ( signal_22799 ) ) ;
    buf_clk cell_8110 ( .C ( clk ), .D ( signal_22802 ), .Q ( signal_22803 ) ) ;
    buf_clk cell_8114 ( .C ( clk ), .D ( signal_22806 ), .Q ( signal_22807 ) ) ;
    buf_clk cell_8120 ( .C ( clk ), .D ( signal_22812 ), .Q ( signal_22813 ) ) ;
    buf_clk cell_8126 ( .C ( clk ), .D ( signal_22818 ), .Q ( signal_22819 ) ) ;
    buf_clk cell_8132 ( .C ( clk ), .D ( signal_22824 ), .Q ( signal_22825 ) ) ;
    buf_clk cell_8138 ( .C ( clk ), .D ( signal_22830 ), .Q ( signal_22831 ) ) ;
    buf_clk cell_8144 ( .C ( clk ), .D ( signal_22836 ), .Q ( signal_22837 ) ) ;
    buf_clk cell_8146 ( .C ( clk ), .D ( signal_22838 ), .Q ( signal_22839 ) ) ;
    buf_clk cell_8148 ( .C ( clk ), .D ( signal_22840 ), .Q ( signal_22841 ) ) ;
    buf_clk cell_8150 ( .C ( clk ), .D ( signal_22842 ), .Q ( signal_22843 ) ) ;
    buf_clk cell_8152 ( .C ( clk ), .D ( signal_22844 ), .Q ( signal_22845 ) ) ;
    buf_clk cell_8154 ( .C ( clk ), .D ( signal_22846 ), .Q ( signal_22847 ) ) ;
    buf_clk cell_8158 ( .C ( clk ), .D ( signal_22850 ), .Q ( signal_22851 ) ) ;
    buf_clk cell_8162 ( .C ( clk ), .D ( signal_22854 ), .Q ( signal_22855 ) ) ;
    buf_clk cell_8166 ( .C ( clk ), .D ( signal_22858 ), .Q ( signal_22859 ) ) ;
    buf_clk cell_8170 ( .C ( clk ), .D ( signal_22862 ), .Q ( signal_22863 ) ) ;
    buf_clk cell_8174 ( .C ( clk ), .D ( signal_22866 ), .Q ( signal_22867 ) ) ;
    buf_clk cell_8178 ( .C ( clk ), .D ( signal_22870 ), .Q ( signal_22871 ) ) ;
    buf_clk cell_8184 ( .C ( clk ), .D ( signal_22876 ), .Q ( signal_22877 ) ) ;
    buf_clk cell_8190 ( .C ( clk ), .D ( signal_22882 ), .Q ( signal_22883 ) ) ;
    buf_clk cell_8196 ( .C ( clk ), .D ( signal_22888 ), .Q ( signal_22889 ) ) ;
    buf_clk cell_8202 ( .C ( clk ), .D ( signal_22894 ), .Q ( signal_22895 ) ) ;
    buf_clk cell_8210 ( .C ( clk ), .D ( signal_22902 ), .Q ( signal_22903 ) ) ;
    buf_clk cell_8218 ( .C ( clk ), .D ( signal_22910 ), .Q ( signal_22911 ) ) ;
    buf_clk cell_8226 ( .C ( clk ), .D ( signal_22918 ), .Q ( signal_22919 ) ) ;
    buf_clk cell_8234 ( .C ( clk ), .D ( signal_22926 ), .Q ( signal_22927 ) ) ;
    buf_clk cell_8242 ( .C ( clk ), .D ( signal_22934 ), .Q ( signal_22935 ) ) ;
    buf_clk cell_8248 ( .C ( clk ), .D ( signal_22940 ), .Q ( signal_22941 ) ) ;
    buf_clk cell_8254 ( .C ( clk ), .D ( signal_22946 ), .Q ( signal_22947 ) ) ;
    buf_clk cell_8260 ( .C ( clk ), .D ( signal_22952 ), .Q ( signal_22953 ) ) ;
    buf_clk cell_8266 ( .C ( clk ), .D ( signal_22958 ), .Q ( signal_22959 ) ) ;
    buf_clk cell_8272 ( .C ( clk ), .D ( signal_22964 ), .Q ( signal_22965 ) ) ;
    buf_clk cell_8282 ( .C ( clk ), .D ( signal_22974 ), .Q ( signal_22975 ) ) ;
    buf_clk cell_8292 ( .C ( clk ), .D ( signal_22984 ), .Q ( signal_22985 ) ) ;
    buf_clk cell_8302 ( .C ( clk ), .D ( signal_22994 ), .Q ( signal_22995 ) ) ;
    buf_clk cell_8312 ( .C ( clk ), .D ( signal_23004 ), .Q ( signal_23005 ) ) ;
    buf_clk cell_8322 ( .C ( clk ), .D ( signal_23014 ), .Q ( signal_23015 ) ) ;
    buf_clk cell_8328 ( .C ( clk ), .D ( signal_23020 ), .Q ( signal_23021 ) ) ;
    buf_clk cell_8334 ( .C ( clk ), .D ( signal_23026 ), .Q ( signal_23027 ) ) ;
    buf_clk cell_8340 ( .C ( clk ), .D ( signal_23032 ), .Q ( signal_23033 ) ) ;
    buf_clk cell_8346 ( .C ( clk ), .D ( signal_23038 ), .Q ( signal_23039 ) ) ;
    buf_clk cell_8352 ( .C ( clk ), .D ( signal_23044 ), .Q ( signal_23045 ) ) ;
    buf_clk cell_8356 ( .C ( clk ), .D ( signal_23048 ), .Q ( signal_23049 ) ) ;
    buf_clk cell_8360 ( .C ( clk ), .D ( signal_23052 ), .Q ( signal_23053 ) ) ;
    buf_clk cell_8364 ( .C ( clk ), .D ( signal_23056 ), .Q ( signal_23057 ) ) ;
    buf_clk cell_8368 ( .C ( clk ), .D ( signal_23060 ), .Q ( signal_23061 ) ) ;
    buf_clk cell_8372 ( .C ( clk ), .D ( signal_23064 ), .Q ( signal_23065 ) ) ;
    buf_clk cell_8380 ( .C ( clk ), .D ( signal_23072 ), .Q ( signal_23073 ) ) ;
    buf_clk cell_8388 ( .C ( clk ), .D ( signal_23080 ), .Q ( signal_23081 ) ) ;
    buf_clk cell_8396 ( .C ( clk ), .D ( signal_23088 ), .Q ( signal_23089 ) ) ;
    buf_clk cell_8404 ( .C ( clk ), .D ( signal_23096 ), .Q ( signal_23097 ) ) ;
    buf_clk cell_8412 ( .C ( clk ), .D ( signal_23104 ), .Q ( signal_23105 ) ) ;
    buf_clk cell_8418 ( .C ( clk ), .D ( signal_23110 ), .Q ( signal_23111 ) ) ;
    buf_clk cell_8424 ( .C ( clk ), .D ( signal_23116 ), .Q ( signal_23117 ) ) ;
    buf_clk cell_8430 ( .C ( clk ), .D ( signal_23122 ), .Q ( signal_23123 ) ) ;
    buf_clk cell_8436 ( .C ( clk ), .D ( signal_23128 ), .Q ( signal_23129 ) ) ;
    buf_clk cell_8442 ( .C ( clk ), .D ( signal_23134 ), .Q ( signal_23135 ) ) ;
    buf_clk cell_8450 ( .C ( clk ), .D ( signal_23142 ), .Q ( signal_23143 ) ) ;
    buf_clk cell_8458 ( .C ( clk ), .D ( signal_23150 ), .Q ( signal_23151 ) ) ;
    buf_clk cell_8466 ( .C ( clk ), .D ( signal_23158 ), .Q ( signal_23159 ) ) ;
    buf_clk cell_8474 ( .C ( clk ), .D ( signal_23166 ), .Q ( signal_23167 ) ) ;
    buf_clk cell_8482 ( .C ( clk ), .D ( signal_23174 ), .Q ( signal_23175 ) ) ;
    buf_clk cell_8488 ( .C ( clk ), .D ( signal_23180 ), .Q ( signal_23181 ) ) ;
    buf_clk cell_8494 ( .C ( clk ), .D ( signal_23186 ), .Q ( signal_23187 ) ) ;
    buf_clk cell_8500 ( .C ( clk ), .D ( signal_23192 ), .Q ( signal_23193 ) ) ;
    buf_clk cell_8506 ( .C ( clk ), .D ( signal_23198 ), .Q ( signal_23199 ) ) ;
    buf_clk cell_8512 ( .C ( clk ), .D ( signal_23204 ), .Q ( signal_23205 ) ) ;
    buf_clk cell_8520 ( .C ( clk ), .D ( signal_23212 ), .Q ( signal_23213 ) ) ;
    buf_clk cell_8528 ( .C ( clk ), .D ( signal_23220 ), .Q ( signal_23221 ) ) ;
    buf_clk cell_8536 ( .C ( clk ), .D ( signal_23228 ), .Q ( signal_23229 ) ) ;
    buf_clk cell_8544 ( .C ( clk ), .D ( signal_23236 ), .Q ( signal_23237 ) ) ;
    buf_clk cell_8552 ( .C ( clk ), .D ( signal_23244 ), .Q ( signal_23245 ) ) ;
    buf_clk cell_8556 ( .C ( clk ), .D ( signal_23248 ), .Q ( signal_23249 ) ) ;
    buf_clk cell_8560 ( .C ( clk ), .D ( signal_23252 ), .Q ( signal_23253 ) ) ;
    buf_clk cell_8564 ( .C ( clk ), .D ( signal_23256 ), .Q ( signal_23257 ) ) ;
    buf_clk cell_8568 ( .C ( clk ), .D ( signal_23260 ), .Q ( signal_23261 ) ) ;
    buf_clk cell_8572 ( .C ( clk ), .D ( signal_23264 ), .Q ( signal_23265 ) ) ;
    buf_clk cell_8578 ( .C ( clk ), .D ( signal_23270 ), .Q ( signal_23271 ) ) ;
    buf_clk cell_8584 ( .C ( clk ), .D ( signal_23276 ), .Q ( signal_23277 ) ) ;
    buf_clk cell_8590 ( .C ( clk ), .D ( signal_23282 ), .Q ( signal_23283 ) ) ;
    buf_clk cell_8596 ( .C ( clk ), .D ( signal_23288 ), .Q ( signal_23289 ) ) ;
    buf_clk cell_8602 ( .C ( clk ), .D ( signal_23294 ), .Q ( signal_23295 ) ) ;
    buf_clk cell_8608 ( .C ( clk ), .D ( signal_23300 ), .Q ( signal_23301 ) ) ;
    buf_clk cell_8614 ( .C ( clk ), .D ( signal_23306 ), .Q ( signal_23307 ) ) ;
    buf_clk cell_8620 ( .C ( clk ), .D ( signal_23312 ), .Q ( signal_23313 ) ) ;
    buf_clk cell_8626 ( .C ( clk ), .D ( signal_23318 ), .Q ( signal_23319 ) ) ;
    buf_clk cell_8632 ( .C ( clk ), .D ( signal_23324 ), .Q ( signal_23325 ) ) ;
    buf_clk cell_8636 ( .C ( clk ), .D ( signal_23328 ), .Q ( signal_23329 ) ) ;
    buf_clk cell_8640 ( .C ( clk ), .D ( signal_23332 ), .Q ( signal_23333 ) ) ;
    buf_clk cell_8644 ( .C ( clk ), .D ( signal_23336 ), .Q ( signal_23337 ) ) ;
    buf_clk cell_8648 ( .C ( clk ), .D ( signal_23340 ), .Q ( signal_23341 ) ) ;
    buf_clk cell_8652 ( .C ( clk ), .D ( signal_23344 ), .Q ( signal_23345 ) ) ;
    buf_clk cell_8656 ( .C ( clk ), .D ( signal_23348 ), .Q ( signal_23349 ) ) ;
    buf_clk cell_8660 ( .C ( clk ), .D ( signal_23352 ), .Q ( signal_23353 ) ) ;
    buf_clk cell_8664 ( .C ( clk ), .D ( signal_23356 ), .Q ( signal_23357 ) ) ;
    buf_clk cell_8668 ( .C ( clk ), .D ( signal_23360 ), .Q ( signal_23361 ) ) ;
    buf_clk cell_8672 ( .C ( clk ), .D ( signal_23364 ), .Q ( signal_23365 ) ) ;
    buf_clk cell_8678 ( .C ( clk ), .D ( signal_23370 ), .Q ( signal_23371 ) ) ;
    buf_clk cell_8686 ( .C ( clk ), .D ( signal_23378 ), .Q ( signal_23379 ) ) ;
    buf_clk cell_8694 ( .C ( clk ), .D ( signal_23386 ), .Q ( signal_23387 ) ) ;
    buf_clk cell_8702 ( .C ( clk ), .D ( signal_23394 ), .Q ( signal_23395 ) ) ;
    buf_clk cell_8710 ( .C ( clk ), .D ( signal_23402 ), .Q ( signal_23403 ) ) ;
    buf_clk cell_8722 ( .C ( clk ), .D ( signal_23414 ), .Q ( signal_23415 ) ) ;
    buf_clk cell_8734 ( .C ( clk ), .D ( signal_23426 ), .Q ( signal_23427 ) ) ;
    buf_clk cell_8746 ( .C ( clk ), .D ( signal_23438 ), .Q ( signal_23439 ) ) ;
    buf_clk cell_8758 ( .C ( clk ), .D ( signal_23450 ), .Q ( signal_23451 ) ) ;
    buf_clk cell_8770 ( .C ( clk ), .D ( signal_23462 ), .Q ( signal_23463 ) ) ;
    buf_clk cell_8776 ( .C ( clk ), .D ( signal_23468 ), .Q ( signal_23469 ) ) ;
    buf_clk cell_8782 ( .C ( clk ), .D ( signal_23474 ), .Q ( signal_23475 ) ) ;
    buf_clk cell_8788 ( .C ( clk ), .D ( signal_23480 ), .Q ( signal_23481 ) ) ;
    buf_clk cell_8794 ( .C ( clk ), .D ( signal_23486 ), .Q ( signal_23487 ) ) ;
    buf_clk cell_8800 ( .C ( clk ), .D ( signal_23492 ), .Q ( signal_23493 ) ) ;
    buf_clk cell_8806 ( .C ( clk ), .D ( signal_23498 ), .Q ( signal_23499 ) ) ;
    buf_clk cell_8812 ( .C ( clk ), .D ( signal_23504 ), .Q ( signal_23505 ) ) ;
    buf_clk cell_8818 ( .C ( clk ), .D ( signal_23510 ), .Q ( signal_23511 ) ) ;
    buf_clk cell_8824 ( .C ( clk ), .D ( signal_23516 ), .Q ( signal_23517 ) ) ;
    buf_clk cell_8830 ( .C ( clk ), .D ( signal_23522 ), .Q ( signal_23523 ) ) ;
    buf_clk cell_8844 ( .C ( clk ), .D ( signal_23536 ), .Q ( signal_23537 ) ) ;
    buf_clk cell_8858 ( .C ( clk ), .D ( signal_23550 ), .Q ( signal_23551 ) ) ;
    buf_clk cell_8872 ( .C ( clk ), .D ( signal_23564 ), .Q ( signal_23565 ) ) ;
    buf_clk cell_8886 ( .C ( clk ), .D ( signal_23578 ), .Q ( signal_23579 ) ) ;
    buf_clk cell_8900 ( .C ( clk ), .D ( signal_23592 ), .Q ( signal_23593 ) ) ;
    buf_clk cell_8908 ( .C ( clk ), .D ( signal_23600 ), .Q ( signal_23601 ) ) ;
    buf_clk cell_8916 ( .C ( clk ), .D ( signal_23608 ), .Q ( signal_23609 ) ) ;
    buf_clk cell_8924 ( .C ( clk ), .D ( signal_23616 ), .Q ( signal_23617 ) ) ;
    buf_clk cell_8932 ( .C ( clk ), .D ( signal_23624 ), .Q ( signal_23625 ) ) ;
    buf_clk cell_8940 ( .C ( clk ), .D ( signal_23632 ), .Q ( signal_23633 ) ) ;
    buf_clk cell_8954 ( .C ( clk ), .D ( signal_23646 ), .Q ( signal_23647 ) ) ;
    buf_clk cell_8968 ( .C ( clk ), .D ( signal_23660 ), .Q ( signal_23661 ) ) ;
    buf_clk cell_8982 ( .C ( clk ), .D ( signal_23674 ), .Q ( signal_23675 ) ) ;
    buf_clk cell_8996 ( .C ( clk ), .D ( signal_23688 ), .Q ( signal_23689 ) ) ;
    buf_clk cell_9010 ( .C ( clk ), .D ( signal_23702 ), .Q ( signal_23703 ) ) ;
    buf_clk cell_9018 ( .C ( clk ), .D ( signal_23710 ), .Q ( signal_23711 ) ) ;
    buf_clk cell_9026 ( .C ( clk ), .D ( signal_23718 ), .Q ( signal_23719 ) ) ;
    buf_clk cell_9034 ( .C ( clk ), .D ( signal_23726 ), .Q ( signal_23727 ) ) ;
    buf_clk cell_9042 ( .C ( clk ), .D ( signal_23734 ), .Q ( signal_23735 ) ) ;
    buf_clk cell_9050 ( .C ( clk ), .D ( signal_23742 ), .Q ( signal_23743 ) ) ;
    buf_clk cell_9078 ( .C ( clk ), .D ( signal_23770 ), .Q ( signal_23771 ) ) ;
    buf_clk cell_9088 ( .C ( clk ), .D ( signal_23780 ), .Q ( signal_23781 ) ) ;
    buf_clk cell_9098 ( .C ( clk ), .D ( signal_23790 ), .Q ( signal_23791 ) ) ;
    buf_clk cell_9108 ( .C ( clk ), .D ( signal_23800 ), .Q ( signal_23801 ) ) ;
    buf_clk cell_9118 ( .C ( clk ), .D ( signal_23810 ), .Q ( signal_23811 ) ) ;
    buf_clk cell_9154 ( .C ( clk ), .D ( signal_23846 ), .Q ( signal_23847 ) ) ;
    buf_clk cell_9170 ( .C ( clk ), .D ( signal_23862 ), .Q ( signal_23863 ) ) ;
    buf_clk cell_9186 ( .C ( clk ), .D ( signal_23878 ), .Q ( signal_23879 ) ) ;
    buf_clk cell_9202 ( .C ( clk ), .D ( signal_23894 ), .Q ( signal_23895 ) ) ;
    buf_clk cell_9218 ( .C ( clk ), .D ( signal_23910 ), .Q ( signal_23911 ) ) ;
    buf_clk cell_9254 ( .C ( clk ), .D ( signal_23946 ), .Q ( signal_23947 ) ) ;
    buf_clk cell_9270 ( .C ( clk ), .D ( signal_23962 ), .Q ( signal_23963 ) ) ;
    buf_clk cell_9286 ( .C ( clk ), .D ( signal_23978 ), .Q ( signal_23979 ) ) ;
    buf_clk cell_9302 ( .C ( clk ), .D ( signal_23994 ), .Q ( signal_23995 ) ) ;
    buf_clk cell_9318 ( .C ( clk ), .D ( signal_24010 ), .Q ( signal_24011 ) ) ;
    buf_clk cell_9328 ( .C ( clk ), .D ( signal_24020 ), .Q ( signal_24021 ) ) ;
    buf_clk cell_9338 ( .C ( clk ), .D ( signal_24030 ), .Q ( signal_24031 ) ) ;
    buf_clk cell_9348 ( .C ( clk ), .D ( signal_24040 ), .Q ( signal_24041 ) ) ;
    buf_clk cell_9358 ( .C ( clk ), .D ( signal_24050 ), .Q ( signal_24051 ) ) ;
    buf_clk cell_9368 ( .C ( clk ), .D ( signal_24060 ), .Q ( signal_24061 ) ) ;
    buf_clk cell_9426 ( .C ( clk ), .D ( signal_24118 ), .Q ( signal_24119 ) ) ;
    buf_clk cell_9436 ( .C ( clk ), .D ( signal_24128 ), .Q ( signal_24129 ) ) ;
    buf_clk cell_9446 ( .C ( clk ), .D ( signal_24138 ), .Q ( signal_24139 ) ) ;
    buf_clk cell_9456 ( .C ( clk ), .D ( signal_24148 ), .Q ( signal_24149 ) ) ;
    buf_clk cell_9466 ( .C ( clk ), .D ( signal_24158 ), .Q ( signal_24159 ) ) ;
    buf_clk cell_9506 ( .C ( clk ), .D ( signal_24198 ), .Q ( signal_24199 ) ) ;
    buf_clk cell_9516 ( .C ( clk ), .D ( signal_24208 ), .Q ( signal_24209 ) ) ;
    buf_clk cell_9526 ( .C ( clk ), .D ( signal_24218 ), .Q ( signal_24219 ) ) ;
    buf_clk cell_9536 ( .C ( clk ), .D ( signal_24228 ), .Q ( signal_24229 ) ) ;
    buf_clk cell_9546 ( .C ( clk ), .D ( signal_24238 ), .Q ( signal_24239 ) ) ;
    buf_clk cell_9562 ( .C ( clk ), .D ( signal_24254 ), .Q ( signal_24255 ) ) ;
    buf_clk cell_9578 ( .C ( clk ), .D ( signal_24270 ), .Q ( signal_24271 ) ) ;
    buf_clk cell_9594 ( .C ( clk ), .D ( signal_24286 ), .Q ( signal_24287 ) ) ;
    buf_clk cell_9610 ( .C ( clk ), .D ( signal_24302 ), .Q ( signal_24303 ) ) ;
    buf_clk cell_9626 ( .C ( clk ), .D ( signal_24318 ), .Q ( signal_24319 ) ) ;
    buf_clk cell_9644 ( .C ( clk ), .D ( signal_24336 ), .Q ( signal_24337 ) ) ;
    buf_clk cell_9662 ( .C ( clk ), .D ( signal_24354 ), .Q ( signal_24355 ) ) ;
    buf_clk cell_9680 ( .C ( clk ), .D ( signal_24372 ), .Q ( signal_24373 ) ) ;
    buf_clk cell_9698 ( .C ( clk ), .D ( signal_24390 ), .Q ( signal_24391 ) ) ;
    buf_clk cell_9716 ( .C ( clk ), .D ( signal_24408 ), .Q ( signal_24409 ) ) ;
    buf_clk cell_9894 ( .C ( clk ), .D ( signal_24586 ), .Q ( signal_24587 ) ) ;
    buf_clk cell_9914 ( .C ( clk ), .D ( signal_24606 ), .Q ( signal_24607 ) ) ;
    buf_clk cell_9934 ( .C ( clk ), .D ( signal_24626 ), .Q ( signal_24627 ) ) ;
    buf_clk cell_9954 ( .C ( clk ), .D ( signal_24646 ), .Q ( signal_24647 ) ) ;
    buf_clk cell_9974 ( .C ( clk ), .D ( signal_24666 ), .Q ( signal_24667 ) ) ;

    /* cells in depth 17 */
    buf_clk cell_8179 ( .C ( clk ), .D ( signal_22871 ), .Q ( signal_22872 ) ) ;
    buf_clk cell_8185 ( .C ( clk ), .D ( signal_22877 ), .Q ( signal_22878 ) ) ;
    buf_clk cell_8191 ( .C ( clk ), .D ( signal_22883 ), .Q ( signal_22884 ) ) ;
    buf_clk cell_8197 ( .C ( clk ), .D ( signal_22889 ), .Q ( signal_22890 ) ) ;
    buf_clk cell_8203 ( .C ( clk ), .D ( signal_22895 ), .Q ( signal_22896 ) ) ;
    buf_clk cell_8211 ( .C ( clk ), .D ( signal_22903 ), .Q ( signal_22904 ) ) ;
    buf_clk cell_8219 ( .C ( clk ), .D ( signal_22911 ), .Q ( signal_22912 ) ) ;
    buf_clk cell_8227 ( .C ( clk ), .D ( signal_22919 ), .Q ( signal_22920 ) ) ;
    buf_clk cell_8235 ( .C ( clk ), .D ( signal_22927 ), .Q ( signal_22928 ) ) ;
    buf_clk cell_8243 ( .C ( clk ), .D ( signal_22935 ), .Q ( signal_22936 ) ) ;
    buf_clk cell_8249 ( .C ( clk ), .D ( signal_22941 ), .Q ( signal_22942 ) ) ;
    buf_clk cell_8255 ( .C ( clk ), .D ( signal_22947 ), .Q ( signal_22948 ) ) ;
    buf_clk cell_8261 ( .C ( clk ), .D ( signal_22953 ), .Q ( signal_22954 ) ) ;
    buf_clk cell_8267 ( .C ( clk ), .D ( signal_22959 ), .Q ( signal_22960 ) ) ;
    buf_clk cell_8273 ( .C ( clk ), .D ( signal_22965 ), .Q ( signal_22966 ) ) ;
    buf_clk cell_8283 ( .C ( clk ), .D ( signal_22975 ), .Q ( signal_22976 ) ) ;
    buf_clk cell_8293 ( .C ( clk ), .D ( signal_22985 ), .Q ( signal_22986 ) ) ;
    buf_clk cell_8303 ( .C ( clk ), .D ( signal_22995 ), .Q ( signal_22996 ) ) ;
    buf_clk cell_8313 ( .C ( clk ), .D ( signal_23005 ), .Q ( signal_23006 ) ) ;
    buf_clk cell_8323 ( .C ( clk ), .D ( signal_23015 ), .Q ( signal_23016 ) ) ;
    buf_clk cell_8329 ( .C ( clk ), .D ( signal_23021 ), .Q ( signal_23022 ) ) ;
    buf_clk cell_8335 ( .C ( clk ), .D ( signal_23027 ), .Q ( signal_23028 ) ) ;
    buf_clk cell_8341 ( .C ( clk ), .D ( signal_23033 ), .Q ( signal_23034 ) ) ;
    buf_clk cell_8347 ( .C ( clk ), .D ( signal_23039 ), .Q ( signal_23040 ) ) ;
    buf_clk cell_8353 ( .C ( clk ), .D ( signal_23045 ), .Q ( signal_23046 ) ) ;
    buf_clk cell_8357 ( .C ( clk ), .D ( signal_23049 ), .Q ( signal_23050 ) ) ;
    buf_clk cell_8361 ( .C ( clk ), .D ( signal_23053 ), .Q ( signal_23054 ) ) ;
    buf_clk cell_8365 ( .C ( clk ), .D ( signal_23057 ), .Q ( signal_23058 ) ) ;
    buf_clk cell_8369 ( .C ( clk ), .D ( signal_23061 ), .Q ( signal_23062 ) ) ;
    buf_clk cell_8373 ( .C ( clk ), .D ( signal_23065 ), .Q ( signal_23066 ) ) ;
    buf_clk cell_8381 ( .C ( clk ), .D ( signal_23073 ), .Q ( signal_23074 ) ) ;
    buf_clk cell_8389 ( .C ( clk ), .D ( signal_23081 ), .Q ( signal_23082 ) ) ;
    buf_clk cell_8397 ( .C ( clk ), .D ( signal_23089 ), .Q ( signal_23090 ) ) ;
    buf_clk cell_8405 ( .C ( clk ), .D ( signal_23097 ), .Q ( signal_23098 ) ) ;
    buf_clk cell_8413 ( .C ( clk ), .D ( signal_23105 ), .Q ( signal_23106 ) ) ;
    buf_clk cell_8419 ( .C ( clk ), .D ( signal_23111 ), .Q ( signal_23112 ) ) ;
    buf_clk cell_8425 ( .C ( clk ), .D ( signal_23117 ), .Q ( signal_23118 ) ) ;
    buf_clk cell_8431 ( .C ( clk ), .D ( signal_23123 ), .Q ( signal_23124 ) ) ;
    buf_clk cell_8437 ( .C ( clk ), .D ( signal_23129 ), .Q ( signal_23130 ) ) ;
    buf_clk cell_8443 ( .C ( clk ), .D ( signal_23135 ), .Q ( signal_23136 ) ) ;
    buf_clk cell_8451 ( .C ( clk ), .D ( signal_23143 ), .Q ( signal_23144 ) ) ;
    buf_clk cell_8459 ( .C ( clk ), .D ( signal_23151 ), .Q ( signal_23152 ) ) ;
    buf_clk cell_8467 ( .C ( clk ), .D ( signal_23159 ), .Q ( signal_23160 ) ) ;
    buf_clk cell_8475 ( .C ( clk ), .D ( signal_23167 ), .Q ( signal_23168 ) ) ;
    buf_clk cell_8483 ( .C ( clk ), .D ( signal_23175 ), .Q ( signal_23176 ) ) ;
    buf_clk cell_8489 ( .C ( clk ), .D ( signal_23181 ), .Q ( signal_23182 ) ) ;
    buf_clk cell_8495 ( .C ( clk ), .D ( signal_23187 ), .Q ( signal_23188 ) ) ;
    buf_clk cell_8501 ( .C ( clk ), .D ( signal_23193 ), .Q ( signal_23194 ) ) ;
    buf_clk cell_8507 ( .C ( clk ), .D ( signal_23199 ), .Q ( signal_23200 ) ) ;
    buf_clk cell_8513 ( .C ( clk ), .D ( signal_23205 ), .Q ( signal_23206 ) ) ;
    buf_clk cell_8521 ( .C ( clk ), .D ( signal_23213 ), .Q ( signal_23214 ) ) ;
    buf_clk cell_8529 ( .C ( clk ), .D ( signal_23221 ), .Q ( signal_23222 ) ) ;
    buf_clk cell_8537 ( .C ( clk ), .D ( signal_23229 ), .Q ( signal_23230 ) ) ;
    buf_clk cell_8545 ( .C ( clk ), .D ( signal_23237 ), .Q ( signal_23238 ) ) ;
    buf_clk cell_8553 ( .C ( clk ), .D ( signal_23245 ), .Q ( signal_23246 ) ) ;
    buf_clk cell_8557 ( .C ( clk ), .D ( signal_23249 ), .Q ( signal_23250 ) ) ;
    buf_clk cell_8561 ( .C ( clk ), .D ( signal_23253 ), .Q ( signal_23254 ) ) ;
    buf_clk cell_8565 ( .C ( clk ), .D ( signal_23257 ), .Q ( signal_23258 ) ) ;
    buf_clk cell_8569 ( .C ( clk ), .D ( signal_23261 ), .Q ( signal_23262 ) ) ;
    buf_clk cell_8573 ( .C ( clk ), .D ( signal_23265 ), .Q ( signal_23266 ) ) ;
    buf_clk cell_8579 ( .C ( clk ), .D ( signal_23271 ), .Q ( signal_23272 ) ) ;
    buf_clk cell_8585 ( .C ( clk ), .D ( signal_23277 ), .Q ( signal_23278 ) ) ;
    buf_clk cell_8591 ( .C ( clk ), .D ( signal_23283 ), .Q ( signal_23284 ) ) ;
    buf_clk cell_8597 ( .C ( clk ), .D ( signal_23289 ), .Q ( signal_23290 ) ) ;
    buf_clk cell_8603 ( .C ( clk ), .D ( signal_23295 ), .Q ( signal_23296 ) ) ;
    buf_clk cell_8609 ( .C ( clk ), .D ( signal_23301 ), .Q ( signal_23302 ) ) ;
    buf_clk cell_8615 ( .C ( clk ), .D ( signal_23307 ), .Q ( signal_23308 ) ) ;
    buf_clk cell_8621 ( .C ( clk ), .D ( signal_23313 ), .Q ( signal_23314 ) ) ;
    buf_clk cell_8627 ( .C ( clk ), .D ( signal_23319 ), .Q ( signal_23320 ) ) ;
    buf_clk cell_8633 ( .C ( clk ), .D ( signal_23325 ), .Q ( signal_23326 ) ) ;
    buf_clk cell_8637 ( .C ( clk ), .D ( signal_23329 ), .Q ( signal_23330 ) ) ;
    buf_clk cell_8641 ( .C ( clk ), .D ( signal_23333 ), .Q ( signal_23334 ) ) ;
    buf_clk cell_8645 ( .C ( clk ), .D ( signal_23337 ), .Q ( signal_23338 ) ) ;
    buf_clk cell_8649 ( .C ( clk ), .D ( signal_23341 ), .Q ( signal_23342 ) ) ;
    buf_clk cell_8653 ( .C ( clk ), .D ( signal_23345 ), .Q ( signal_23346 ) ) ;
    buf_clk cell_8657 ( .C ( clk ), .D ( signal_23349 ), .Q ( signal_23350 ) ) ;
    buf_clk cell_8661 ( .C ( clk ), .D ( signal_23353 ), .Q ( signal_23354 ) ) ;
    buf_clk cell_8665 ( .C ( clk ), .D ( signal_23357 ), .Q ( signal_23358 ) ) ;
    buf_clk cell_8669 ( .C ( clk ), .D ( signal_23361 ), .Q ( signal_23362 ) ) ;
    buf_clk cell_8673 ( .C ( clk ), .D ( signal_23365 ), .Q ( signal_23366 ) ) ;
    buf_clk cell_8679 ( .C ( clk ), .D ( signal_23371 ), .Q ( signal_23372 ) ) ;
    buf_clk cell_8687 ( .C ( clk ), .D ( signal_23379 ), .Q ( signal_23380 ) ) ;
    buf_clk cell_8695 ( .C ( clk ), .D ( signal_23387 ), .Q ( signal_23388 ) ) ;
    buf_clk cell_8703 ( .C ( clk ), .D ( signal_23395 ), .Q ( signal_23396 ) ) ;
    buf_clk cell_8711 ( .C ( clk ), .D ( signal_23403 ), .Q ( signal_23404 ) ) ;
    buf_clk cell_8723 ( .C ( clk ), .D ( signal_23415 ), .Q ( signal_23416 ) ) ;
    buf_clk cell_8735 ( .C ( clk ), .D ( signal_23427 ), .Q ( signal_23428 ) ) ;
    buf_clk cell_8747 ( .C ( clk ), .D ( signal_23439 ), .Q ( signal_23440 ) ) ;
    buf_clk cell_8759 ( .C ( clk ), .D ( signal_23451 ), .Q ( signal_23452 ) ) ;
    buf_clk cell_8771 ( .C ( clk ), .D ( signal_23463 ), .Q ( signal_23464 ) ) ;
    buf_clk cell_8777 ( .C ( clk ), .D ( signal_23469 ), .Q ( signal_23470 ) ) ;
    buf_clk cell_8783 ( .C ( clk ), .D ( signal_23475 ), .Q ( signal_23476 ) ) ;
    buf_clk cell_8789 ( .C ( clk ), .D ( signal_23481 ), .Q ( signal_23482 ) ) ;
    buf_clk cell_8795 ( .C ( clk ), .D ( signal_23487 ), .Q ( signal_23488 ) ) ;
    buf_clk cell_8801 ( .C ( clk ), .D ( signal_23493 ), .Q ( signal_23494 ) ) ;
    buf_clk cell_8807 ( .C ( clk ), .D ( signal_23499 ), .Q ( signal_23500 ) ) ;
    buf_clk cell_8813 ( .C ( clk ), .D ( signal_23505 ), .Q ( signal_23506 ) ) ;
    buf_clk cell_8819 ( .C ( clk ), .D ( signal_23511 ), .Q ( signal_23512 ) ) ;
    buf_clk cell_8825 ( .C ( clk ), .D ( signal_23517 ), .Q ( signal_23518 ) ) ;
    buf_clk cell_8831 ( .C ( clk ), .D ( signal_23523 ), .Q ( signal_23524 ) ) ;
    buf_clk cell_8845 ( .C ( clk ), .D ( signal_23537 ), .Q ( signal_23538 ) ) ;
    buf_clk cell_8859 ( .C ( clk ), .D ( signal_23551 ), .Q ( signal_23552 ) ) ;
    buf_clk cell_8873 ( .C ( clk ), .D ( signal_23565 ), .Q ( signal_23566 ) ) ;
    buf_clk cell_8887 ( .C ( clk ), .D ( signal_23579 ), .Q ( signal_23580 ) ) ;
    buf_clk cell_8901 ( .C ( clk ), .D ( signal_23593 ), .Q ( signal_23594 ) ) ;
    buf_clk cell_8909 ( .C ( clk ), .D ( signal_23601 ), .Q ( signal_23602 ) ) ;
    buf_clk cell_8917 ( .C ( clk ), .D ( signal_23609 ), .Q ( signal_23610 ) ) ;
    buf_clk cell_8925 ( .C ( clk ), .D ( signal_23617 ), .Q ( signal_23618 ) ) ;
    buf_clk cell_8933 ( .C ( clk ), .D ( signal_23625 ), .Q ( signal_23626 ) ) ;
    buf_clk cell_8941 ( .C ( clk ), .D ( signal_23633 ), .Q ( signal_23634 ) ) ;
    buf_clk cell_8955 ( .C ( clk ), .D ( signal_23647 ), .Q ( signal_23648 ) ) ;
    buf_clk cell_8969 ( .C ( clk ), .D ( signal_23661 ), .Q ( signal_23662 ) ) ;
    buf_clk cell_8983 ( .C ( clk ), .D ( signal_23675 ), .Q ( signal_23676 ) ) ;
    buf_clk cell_8997 ( .C ( clk ), .D ( signal_23689 ), .Q ( signal_23690 ) ) ;
    buf_clk cell_9011 ( .C ( clk ), .D ( signal_23703 ), .Q ( signal_23704 ) ) ;
    buf_clk cell_9019 ( .C ( clk ), .D ( signal_23711 ), .Q ( signal_23712 ) ) ;
    buf_clk cell_9027 ( .C ( clk ), .D ( signal_23719 ), .Q ( signal_23720 ) ) ;
    buf_clk cell_9035 ( .C ( clk ), .D ( signal_23727 ), .Q ( signal_23728 ) ) ;
    buf_clk cell_9043 ( .C ( clk ), .D ( signal_23735 ), .Q ( signal_23736 ) ) ;
    buf_clk cell_9051 ( .C ( clk ), .D ( signal_23743 ), .Q ( signal_23744 ) ) ;
    buf_clk cell_9079 ( .C ( clk ), .D ( signal_23771 ), .Q ( signal_23772 ) ) ;
    buf_clk cell_9089 ( .C ( clk ), .D ( signal_23781 ), .Q ( signal_23782 ) ) ;
    buf_clk cell_9099 ( .C ( clk ), .D ( signal_23791 ), .Q ( signal_23792 ) ) ;
    buf_clk cell_9109 ( .C ( clk ), .D ( signal_23801 ), .Q ( signal_23802 ) ) ;
    buf_clk cell_9119 ( .C ( clk ), .D ( signal_23811 ), .Q ( signal_23812 ) ) ;
    buf_clk cell_9155 ( .C ( clk ), .D ( signal_23847 ), .Q ( signal_23848 ) ) ;
    buf_clk cell_9171 ( .C ( clk ), .D ( signal_23863 ), .Q ( signal_23864 ) ) ;
    buf_clk cell_9187 ( .C ( clk ), .D ( signal_23879 ), .Q ( signal_23880 ) ) ;
    buf_clk cell_9203 ( .C ( clk ), .D ( signal_23895 ), .Q ( signal_23896 ) ) ;
    buf_clk cell_9219 ( .C ( clk ), .D ( signal_23911 ), .Q ( signal_23912 ) ) ;
    buf_clk cell_9255 ( .C ( clk ), .D ( signal_23947 ), .Q ( signal_23948 ) ) ;
    buf_clk cell_9271 ( .C ( clk ), .D ( signal_23963 ), .Q ( signal_23964 ) ) ;
    buf_clk cell_9287 ( .C ( clk ), .D ( signal_23979 ), .Q ( signal_23980 ) ) ;
    buf_clk cell_9303 ( .C ( clk ), .D ( signal_23995 ), .Q ( signal_23996 ) ) ;
    buf_clk cell_9319 ( .C ( clk ), .D ( signal_24011 ), .Q ( signal_24012 ) ) ;
    buf_clk cell_9329 ( .C ( clk ), .D ( signal_24021 ), .Q ( signal_24022 ) ) ;
    buf_clk cell_9339 ( .C ( clk ), .D ( signal_24031 ), .Q ( signal_24032 ) ) ;
    buf_clk cell_9349 ( .C ( clk ), .D ( signal_24041 ), .Q ( signal_24042 ) ) ;
    buf_clk cell_9359 ( .C ( clk ), .D ( signal_24051 ), .Q ( signal_24052 ) ) ;
    buf_clk cell_9369 ( .C ( clk ), .D ( signal_24061 ), .Q ( signal_24062 ) ) ;
    buf_clk cell_9427 ( .C ( clk ), .D ( signal_24119 ), .Q ( signal_24120 ) ) ;
    buf_clk cell_9437 ( .C ( clk ), .D ( signal_24129 ), .Q ( signal_24130 ) ) ;
    buf_clk cell_9447 ( .C ( clk ), .D ( signal_24139 ), .Q ( signal_24140 ) ) ;
    buf_clk cell_9457 ( .C ( clk ), .D ( signal_24149 ), .Q ( signal_24150 ) ) ;
    buf_clk cell_9467 ( .C ( clk ), .D ( signal_24159 ), .Q ( signal_24160 ) ) ;
    buf_clk cell_9507 ( .C ( clk ), .D ( signal_24199 ), .Q ( signal_24200 ) ) ;
    buf_clk cell_9517 ( .C ( clk ), .D ( signal_24209 ), .Q ( signal_24210 ) ) ;
    buf_clk cell_9527 ( .C ( clk ), .D ( signal_24219 ), .Q ( signal_24220 ) ) ;
    buf_clk cell_9537 ( .C ( clk ), .D ( signal_24229 ), .Q ( signal_24230 ) ) ;
    buf_clk cell_9547 ( .C ( clk ), .D ( signal_24239 ), .Q ( signal_24240 ) ) ;
    buf_clk cell_9563 ( .C ( clk ), .D ( signal_24255 ), .Q ( signal_24256 ) ) ;
    buf_clk cell_9579 ( .C ( clk ), .D ( signal_24271 ), .Q ( signal_24272 ) ) ;
    buf_clk cell_9595 ( .C ( clk ), .D ( signal_24287 ), .Q ( signal_24288 ) ) ;
    buf_clk cell_9611 ( .C ( clk ), .D ( signal_24303 ), .Q ( signal_24304 ) ) ;
    buf_clk cell_9627 ( .C ( clk ), .D ( signal_24319 ), .Q ( signal_24320 ) ) ;
    buf_clk cell_9645 ( .C ( clk ), .D ( signal_24337 ), .Q ( signal_24338 ) ) ;
    buf_clk cell_9663 ( .C ( clk ), .D ( signal_24355 ), .Q ( signal_24356 ) ) ;
    buf_clk cell_9681 ( .C ( clk ), .D ( signal_24373 ), .Q ( signal_24374 ) ) ;
    buf_clk cell_9699 ( .C ( clk ), .D ( signal_24391 ), .Q ( signal_24392 ) ) ;
    buf_clk cell_9717 ( .C ( clk ), .D ( signal_24409 ), .Q ( signal_24410 ) ) ;
    buf_clk cell_9745 ( .C ( clk ), .D ( signal_2281 ), .Q ( signal_24438 ) ) ;
    buf_clk cell_9753 ( .C ( clk ), .D ( signal_7780 ), .Q ( signal_24446 ) ) ;
    buf_clk cell_9761 ( .C ( clk ), .D ( signal_7781 ), .Q ( signal_24454 ) ) ;
    buf_clk cell_9769 ( .C ( clk ), .D ( signal_7782 ), .Q ( signal_24462 ) ) ;
    buf_clk cell_9777 ( .C ( clk ), .D ( signal_7783 ), .Q ( signal_24470 ) ) ;
    buf_clk cell_9895 ( .C ( clk ), .D ( signal_24587 ), .Q ( signal_24588 ) ) ;
    buf_clk cell_9915 ( .C ( clk ), .D ( signal_24607 ), .Q ( signal_24608 ) ) ;
    buf_clk cell_9935 ( .C ( clk ), .D ( signal_24627 ), .Q ( signal_24628 ) ) ;
    buf_clk cell_9955 ( .C ( clk ), .D ( signal_24647 ), .Q ( signal_24648 ) ) ;
    buf_clk cell_9975 ( .C ( clk ), .D ( signal_24667 ), .Q ( signal_24668 ) ) ;
    buf_clk cell_10025 ( .C ( clk ), .D ( signal_2260 ), .Q ( signal_24718 ) ) ;
    buf_clk cell_10037 ( .C ( clk ), .D ( signal_7696 ), .Q ( signal_24730 ) ) ;
    buf_clk cell_10049 ( .C ( clk ), .D ( signal_7697 ), .Q ( signal_24742 ) ) ;
    buf_clk cell_10061 ( .C ( clk ), .D ( signal_7698 ), .Q ( signal_24754 ) ) ;
    buf_clk cell_10073 ( .C ( clk ), .D ( signal_7699 ), .Q ( signal_24766 ) ) ;
    buf_clk cell_10085 ( .C ( clk ), .D ( signal_2322 ), .Q ( signal_24778 ) ) ;
    buf_clk cell_10099 ( .C ( clk ), .D ( signal_7944 ), .Q ( signal_24792 ) ) ;
    buf_clk cell_10113 ( .C ( clk ), .D ( signal_7945 ), .Q ( signal_24806 ) ) ;
    buf_clk cell_10127 ( .C ( clk ), .D ( signal_7946 ), .Q ( signal_24820 ) ) ;
    buf_clk cell_10141 ( .C ( clk ), .D ( signal_7947 ), .Q ( signal_24834 ) ) ;

    /* cells in depth 18 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2230 ( .a ({signal_22247, signal_22241, signal_22235, signal_22229, signal_22223}), .b ({signal_7443, signal_7442, signal_7441, signal_7440, signal_2196}), .clk ( clk ), .r ({Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010]}), .c ({signal_7639, signal_7638, signal_7637, signal_7636, signal_2245}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2231 ( .a ({signal_22287, signal_22279, signal_22271, signal_22263, signal_22255}), .b ({signal_7447, signal_7446, signal_7445, signal_7444, signal_2197}), .clk ( clk ), .r ({Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020]}), .c ({signal_7643, signal_7642, signal_7641, signal_7640, signal_2246}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2232 ( .a ({signal_22317, signal_22311, signal_22305, signal_22299, signal_22293}), .b ({signal_7451, signal_7450, signal_7449, signal_7448, signal_2198}), .clk ( clk ), .r ({Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030]}), .c ({signal_7647, signal_7646, signal_7645, signal_7644, signal_2247}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2267 ( .a ({signal_22347, signal_22341, signal_22335, signal_22329, signal_22323}), .b ({signal_7623, signal_7622, signal_7621, signal_7620, signal_2241}), .clk ( clk ), .r ({Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040]}), .c ({signal_7787, signal_7786, signal_7785, signal_7784, signal_2282}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2268 ( .a ({signal_22387, signal_22379, signal_22371, signal_22363, signal_22355}), .b ({signal_7515, signal_7514, signal_7513, signal_7512, signal_2214}), .clk ( clk ), .r ({Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050]}), .c ({signal_7791, signal_7790, signal_7789, signal_7788, signal_2283}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2281 ( .a ({signal_7791, signal_7790, signal_7789, signal_7788, signal_2283}), .b ({signal_7843, signal_7842, signal_7841, signal_7840, signal_2296}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2284 ( .a ({signal_22437, signal_22427, signal_22417, signal_22407, signal_22397}), .b ({signal_7707, signal_7706, signal_7705, signal_7704, signal_2262}), .clk ( clk ), .r ({Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060]}), .c ({signal_7855, signal_7854, signal_7853, signal_7852, signal_2299}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2289 ( .a ({signal_22447, signal_22445, signal_22443, signal_22441, signal_22439}), .b ({signal_7695, signal_7694, signal_7693, signal_7692, signal_2259}), .clk ( clk ), .r ({Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070]}), .c ({signal_7875, signal_7874, signal_7873, signal_7872, signal_2304}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2291 ( .a ({signal_22477, signal_22471, signal_22465, signal_22459, signal_22453}), .b ({signal_7739, signal_7738, signal_7737, signal_7736, signal_2270}), .clk ( clk ), .r ({Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080]}), .c ({signal_7883, signal_7882, signal_7881, signal_7880, signal_2306}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2292 ( .a ({signal_22517, signal_22509, signal_22501, signal_22493, signal_22485}), .b ({signal_7751, signal_7750, signal_7749, signal_7748, signal_2273}), .clk ( clk ), .r ({Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090]}), .c ({signal_7887, signal_7886, signal_7885, signal_7884, signal_2307}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2293 ( .a ({signal_22567, signal_22557, signal_22547, signal_22537, signal_22527}), .b ({signal_7759, signal_7758, signal_7757, signal_7756, signal_2275}), .clk ( clk ), .r ({Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100]}), .c ({signal_7891, signal_7890, signal_7889, signal_7888, signal_2308}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2294 ( .a ({signal_22607, signal_22599, signal_22591, signal_22583, signal_22575}), .b ({signal_7771, signal_7770, signal_7769, signal_7768, signal_2278}), .clk ( clk ), .r ({Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110]}), .c ({signal_7895, signal_7894, signal_7893, signal_7892, signal_2309}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2295 ( .a ({signal_22637, signal_22631, signal_22625, signal_22619, signal_22613}), .b ({signal_7703, signal_7702, signal_7701, signal_7700, signal_2261}), .clk ( clk ), .r ({Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120]}), .c ({signal_7899, signal_7898, signal_7897, signal_7896, signal_2310}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2298 ( .a ({signal_7855, signal_7854, signal_7853, signal_7852, signal_2299}), .b ({signal_7911, signal_7910, signal_7909, signal_7908, signal_2313}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2300 ( .a ({signal_7875, signal_7874, signal_7873, signal_7872, signal_2304}), .b ({signal_7919, signal_7918, signal_7917, signal_7916, signal_2315}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2302 ( .a ({signal_7895, signal_7894, signal_7893, signal_7892, signal_2309}), .b ({signal_7927, signal_7926, signal_7925, signal_7924, signal_2317}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2303 ( .a ({signal_7899, signal_7898, signal_7897, signal_7896, signal_2310}), .b ({signal_7931, signal_7930, signal_7929, signal_7928, signal_2318}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2308 ( .a ({signal_22667, signal_22661, signal_22655, signal_22649, signal_22643}), .b ({signal_7819, signal_7818, signal_7817, signal_7816, signal_2290}), .clk ( clk ), .r ({Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130]}), .c ({signal_7951, signal_7950, signal_7949, signal_7948, signal_2323}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2309 ( .a ({signal_22677, signal_22675, signal_22673, signal_22671, signal_22669}), .b ({signal_7823, signal_7822, signal_7821, signal_7820, signal_2291}), .clk ( clk ), .r ({Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140]}), .c ({signal_7955, signal_7954, signal_7953, signal_7952, signal_2324}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2310 ( .a ({signal_22677, signal_22675, signal_22673, signal_22671, signal_22669}), .b ({signal_7827, signal_7826, signal_7825, signal_7824, signal_2292}), .clk ( clk ), .r ({Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150]}), .c ({signal_7959, signal_7958, signal_7957, signal_7956, signal_2325}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2311 ( .a ({signal_22697, signal_22693, signal_22689, signal_22685, signal_22681}), .b ({signal_7831, signal_7830, signal_7829, signal_7828, signal_2293}), .clk ( clk ), .r ({Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160]}), .c ({signal_7963, signal_7962, signal_7961, signal_7960, signal_2326}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2312 ( .a ({signal_22717, signal_22713, signal_22709, signal_22705, signal_22701}), .b ({signal_7835, signal_7834, signal_7833, signal_7832, signal_2294}), .clk ( clk ), .r ({Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175], Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170]}), .c ({signal_7967, signal_7966, signal_7965, signal_7964, signal_2327}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2313 ( .a ({signal_7867, signal_7866, signal_7865, signal_7864, signal_2302}), .b ({signal_7775, signal_7774, signal_7773, signal_7772, signal_2279}), .clk ( clk ), .r ({Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180]}), .c ({signal_7971, signal_7970, signal_7969, signal_7968, signal_2328}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2314 ( .a ({signal_22747, signal_22741, signal_22735, signal_22729, signal_22723}), .b ({signal_7839, signal_7838, signal_7837, signal_7836, signal_2295}), .clk ( clk ), .r ({Fresh[8199], Fresh[8198], Fresh[8197], Fresh[8196], Fresh[8195], Fresh[8194], Fresh[8193], Fresh[8192], Fresh[8191], Fresh[8190]}), .c ({signal_7975, signal_7974, signal_7973, signal_7972, signal_2329}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2315 ( .a ({signal_22757, signal_22755, signal_22753, signal_22751, signal_22749}), .b ({signal_7631, signal_7630, signal_7629, signal_7628, signal_2243}), .clk ( clk ), .r ({Fresh[8209], Fresh[8208], Fresh[8207], Fresh[8206], Fresh[8205], Fresh[8204], Fresh[8203], Fresh[8202], Fresh[8201], Fresh[8200]}), .c ({signal_7979, signal_7978, signal_7977, signal_7976, signal_2330}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2320 ( .a ({signal_7951, signal_7950, signal_7949, signal_7948, signal_2323}), .b ({signal_7999, signal_7998, signal_7997, signal_7996, signal_2335}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2321 ( .a ({signal_7955, signal_7954, signal_7953, signal_7952, signal_2324}), .b ({signal_8003, signal_8002, signal_8001, signal_8000, signal_2336}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2322 ( .a ({signal_7959, signal_7958, signal_7957, signal_7956, signal_2325}), .b ({signal_8007, signal_8006, signal_8005, signal_8004, signal_2337}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2323 ( .a ({signal_7963, signal_7962, signal_7961, signal_7960, signal_2326}), .b ({signal_8011, signal_8010, signal_8009, signal_8008, signal_2338}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2324 ( .a ({signal_22787, signal_22781, signal_22775, signal_22769, signal_22763}), .b ({signal_7935, signal_7934, signal_7933, signal_7932, signal_2319}), .clk ( clk ), .r ({Fresh[8219], Fresh[8218], Fresh[8217], Fresh[8216], Fresh[8215], Fresh[8214], Fresh[8213], Fresh[8212], Fresh[8211], Fresh[8210]}), .c ({signal_8015, signal_8014, signal_8013, signal_8012, signal_2339}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2326 ( .a ({signal_22807, signal_22803, signal_22799, signal_22795, signal_22791}), .b ({signal_7915, signal_7914, signal_7913, signal_7912, signal_2314}), .clk ( clk ), .r ({Fresh[8229], Fresh[8228], Fresh[8227], Fresh[8226], Fresh[8225], Fresh[8224], Fresh[8223], Fresh[8222], Fresh[8221], Fresh[8220]}), .c ({signal_8023, signal_8022, signal_8021, signal_8020, signal_2341}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2328 ( .a ({signal_22837, signal_22831, signal_22825, signal_22819, signal_22813}), .b ({signal_7939, signal_7938, signal_7937, signal_7936, signal_2320}), .clk ( clk ), .r ({Fresh[8239], Fresh[8238], Fresh[8237], Fresh[8236], Fresh[8235], Fresh[8234], Fresh[8233], Fresh[8232], Fresh[8231], Fresh[8230]}), .c ({signal_8031, signal_8030, signal_8029, signal_8028, signal_2343}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2329 ( .a ({signal_22847, signal_22845, signal_22843, signal_22841, signal_22839}), .b ({signal_7943, signal_7942, signal_7941, signal_7940, signal_2321}), .clk ( clk ), .r ({Fresh[8249], Fresh[8248], Fresh[8247], Fresh[8246], Fresh[8245], Fresh[8244], Fresh[8243], Fresh[8242], Fresh[8241], Fresh[8240]}), .c ({signal_8035, signal_8034, signal_8033, signal_8032, signal_2344}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2330 ( .a ({signal_22867, signal_22863, signal_22859, signal_22855, signal_22851}), .b ({signal_7923, signal_7922, signal_7921, signal_7920, signal_2316}), .clk ( clk ), .r ({Fresh[8259], Fresh[8258], Fresh[8257], Fresh[8256], Fresh[8255], Fresh[8254], Fresh[8253], Fresh[8252], Fresh[8251], Fresh[8250]}), .c ({signal_8039, signal_8038, signal_8037, signal_8036, signal_2345}) ) ;
    buf_clk cell_8180 ( .C ( clk ), .D ( signal_22872 ), .Q ( signal_22873 ) ) ;
    buf_clk cell_8186 ( .C ( clk ), .D ( signal_22878 ), .Q ( signal_22879 ) ) ;
    buf_clk cell_8192 ( .C ( clk ), .D ( signal_22884 ), .Q ( signal_22885 ) ) ;
    buf_clk cell_8198 ( .C ( clk ), .D ( signal_22890 ), .Q ( signal_22891 ) ) ;
    buf_clk cell_8204 ( .C ( clk ), .D ( signal_22896 ), .Q ( signal_22897 ) ) ;
    buf_clk cell_8212 ( .C ( clk ), .D ( signal_22904 ), .Q ( signal_22905 ) ) ;
    buf_clk cell_8220 ( .C ( clk ), .D ( signal_22912 ), .Q ( signal_22913 ) ) ;
    buf_clk cell_8228 ( .C ( clk ), .D ( signal_22920 ), .Q ( signal_22921 ) ) ;
    buf_clk cell_8236 ( .C ( clk ), .D ( signal_22928 ), .Q ( signal_22929 ) ) ;
    buf_clk cell_8244 ( .C ( clk ), .D ( signal_22936 ), .Q ( signal_22937 ) ) ;
    buf_clk cell_8250 ( .C ( clk ), .D ( signal_22942 ), .Q ( signal_22943 ) ) ;
    buf_clk cell_8256 ( .C ( clk ), .D ( signal_22948 ), .Q ( signal_22949 ) ) ;
    buf_clk cell_8262 ( .C ( clk ), .D ( signal_22954 ), .Q ( signal_22955 ) ) ;
    buf_clk cell_8268 ( .C ( clk ), .D ( signal_22960 ), .Q ( signal_22961 ) ) ;
    buf_clk cell_8274 ( .C ( clk ), .D ( signal_22966 ), .Q ( signal_22967 ) ) ;
    buf_clk cell_8284 ( .C ( clk ), .D ( signal_22976 ), .Q ( signal_22977 ) ) ;
    buf_clk cell_8294 ( .C ( clk ), .D ( signal_22986 ), .Q ( signal_22987 ) ) ;
    buf_clk cell_8304 ( .C ( clk ), .D ( signal_22996 ), .Q ( signal_22997 ) ) ;
    buf_clk cell_8314 ( .C ( clk ), .D ( signal_23006 ), .Q ( signal_23007 ) ) ;
    buf_clk cell_8324 ( .C ( clk ), .D ( signal_23016 ), .Q ( signal_23017 ) ) ;
    buf_clk cell_8330 ( .C ( clk ), .D ( signal_23022 ), .Q ( signal_23023 ) ) ;
    buf_clk cell_8336 ( .C ( clk ), .D ( signal_23028 ), .Q ( signal_23029 ) ) ;
    buf_clk cell_8342 ( .C ( clk ), .D ( signal_23034 ), .Q ( signal_23035 ) ) ;
    buf_clk cell_8348 ( .C ( clk ), .D ( signal_23040 ), .Q ( signal_23041 ) ) ;
    buf_clk cell_8354 ( .C ( clk ), .D ( signal_23046 ), .Q ( signal_23047 ) ) ;
    buf_clk cell_8358 ( .C ( clk ), .D ( signal_23050 ), .Q ( signal_23051 ) ) ;
    buf_clk cell_8362 ( .C ( clk ), .D ( signal_23054 ), .Q ( signal_23055 ) ) ;
    buf_clk cell_8366 ( .C ( clk ), .D ( signal_23058 ), .Q ( signal_23059 ) ) ;
    buf_clk cell_8370 ( .C ( clk ), .D ( signal_23062 ), .Q ( signal_23063 ) ) ;
    buf_clk cell_8374 ( .C ( clk ), .D ( signal_23066 ), .Q ( signal_23067 ) ) ;
    buf_clk cell_8382 ( .C ( clk ), .D ( signal_23074 ), .Q ( signal_23075 ) ) ;
    buf_clk cell_8390 ( .C ( clk ), .D ( signal_23082 ), .Q ( signal_23083 ) ) ;
    buf_clk cell_8398 ( .C ( clk ), .D ( signal_23090 ), .Q ( signal_23091 ) ) ;
    buf_clk cell_8406 ( .C ( clk ), .D ( signal_23098 ), .Q ( signal_23099 ) ) ;
    buf_clk cell_8414 ( .C ( clk ), .D ( signal_23106 ), .Q ( signal_23107 ) ) ;
    buf_clk cell_8420 ( .C ( clk ), .D ( signal_23112 ), .Q ( signal_23113 ) ) ;
    buf_clk cell_8426 ( .C ( clk ), .D ( signal_23118 ), .Q ( signal_23119 ) ) ;
    buf_clk cell_8432 ( .C ( clk ), .D ( signal_23124 ), .Q ( signal_23125 ) ) ;
    buf_clk cell_8438 ( .C ( clk ), .D ( signal_23130 ), .Q ( signal_23131 ) ) ;
    buf_clk cell_8444 ( .C ( clk ), .D ( signal_23136 ), .Q ( signal_23137 ) ) ;
    buf_clk cell_8452 ( .C ( clk ), .D ( signal_23144 ), .Q ( signal_23145 ) ) ;
    buf_clk cell_8460 ( .C ( clk ), .D ( signal_23152 ), .Q ( signal_23153 ) ) ;
    buf_clk cell_8468 ( .C ( clk ), .D ( signal_23160 ), .Q ( signal_23161 ) ) ;
    buf_clk cell_8476 ( .C ( clk ), .D ( signal_23168 ), .Q ( signal_23169 ) ) ;
    buf_clk cell_8484 ( .C ( clk ), .D ( signal_23176 ), .Q ( signal_23177 ) ) ;
    buf_clk cell_8490 ( .C ( clk ), .D ( signal_23182 ), .Q ( signal_23183 ) ) ;
    buf_clk cell_8496 ( .C ( clk ), .D ( signal_23188 ), .Q ( signal_23189 ) ) ;
    buf_clk cell_8502 ( .C ( clk ), .D ( signal_23194 ), .Q ( signal_23195 ) ) ;
    buf_clk cell_8508 ( .C ( clk ), .D ( signal_23200 ), .Q ( signal_23201 ) ) ;
    buf_clk cell_8514 ( .C ( clk ), .D ( signal_23206 ), .Q ( signal_23207 ) ) ;
    buf_clk cell_8522 ( .C ( clk ), .D ( signal_23214 ), .Q ( signal_23215 ) ) ;
    buf_clk cell_8530 ( .C ( clk ), .D ( signal_23222 ), .Q ( signal_23223 ) ) ;
    buf_clk cell_8538 ( .C ( clk ), .D ( signal_23230 ), .Q ( signal_23231 ) ) ;
    buf_clk cell_8546 ( .C ( clk ), .D ( signal_23238 ), .Q ( signal_23239 ) ) ;
    buf_clk cell_8554 ( .C ( clk ), .D ( signal_23246 ), .Q ( signal_23247 ) ) ;
    buf_clk cell_8558 ( .C ( clk ), .D ( signal_23250 ), .Q ( signal_23251 ) ) ;
    buf_clk cell_8562 ( .C ( clk ), .D ( signal_23254 ), .Q ( signal_23255 ) ) ;
    buf_clk cell_8566 ( .C ( clk ), .D ( signal_23258 ), .Q ( signal_23259 ) ) ;
    buf_clk cell_8570 ( .C ( clk ), .D ( signal_23262 ), .Q ( signal_23263 ) ) ;
    buf_clk cell_8574 ( .C ( clk ), .D ( signal_23266 ), .Q ( signal_23267 ) ) ;
    buf_clk cell_8580 ( .C ( clk ), .D ( signal_23272 ), .Q ( signal_23273 ) ) ;
    buf_clk cell_8586 ( .C ( clk ), .D ( signal_23278 ), .Q ( signal_23279 ) ) ;
    buf_clk cell_8592 ( .C ( clk ), .D ( signal_23284 ), .Q ( signal_23285 ) ) ;
    buf_clk cell_8598 ( .C ( clk ), .D ( signal_23290 ), .Q ( signal_23291 ) ) ;
    buf_clk cell_8604 ( .C ( clk ), .D ( signal_23296 ), .Q ( signal_23297 ) ) ;
    buf_clk cell_8610 ( .C ( clk ), .D ( signal_23302 ), .Q ( signal_23303 ) ) ;
    buf_clk cell_8616 ( .C ( clk ), .D ( signal_23308 ), .Q ( signal_23309 ) ) ;
    buf_clk cell_8622 ( .C ( clk ), .D ( signal_23314 ), .Q ( signal_23315 ) ) ;
    buf_clk cell_8628 ( .C ( clk ), .D ( signal_23320 ), .Q ( signal_23321 ) ) ;
    buf_clk cell_8634 ( .C ( clk ), .D ( signal_23326 ), .Q ( signal_23327 ) ) ;
    buf_clk cell_8638 ( .C ( clk ), .D ( signal_23330 ), .Q ( signal_23331 ) ) ;
    buf_clk cell_8642 ( .C ( clk ), .D ( signal_23334 ), .Q ( signal_23335 ) ) ;
    buf_clk cell_8646 ( .C ( clk ), .D ( signal_23338 ), .Q ( signal_23339 ) ) ;
    buf_clk cell_8650 ( .C ( clk ), .D ( signal_23342 ), .Q ( signal_23343 ) ) ;
    buf_clk cell_8654 ( .C ( clk ), .D ( signal_23346 ), .Q ( signal_23347 ) ) ;
    buf_clk cell_8658 ( .C ( clk ), .D ( signal_23350 ), .Q ( signal_23351 ) ) ;
    buf_clk cell_8662 ( .C ( clk ), .D ( signal_23354 ), .Q ( signal_23355 ) ) ;
    buf_clk cell_8666 ( .C ( clk ), .D ( signal_23358 ), .Q ( signal_23359 ) ) ;
    buf_clk cell_8670 ( .C ( clk ), .D ( signal_23362 ), .Q ( signal_23363 ) ) ;
    buf_clk cell_8674 ( .C ( clk ), .D ( signal_23366 ), .Q ( signal_23367 ) ) ;
    buf_clk cell_8680 ( .C ( clk ), .D ( signal_23372 ), .Q ( signal_23373 ) ) ;
    buf_clk cell_8688 ( .C ( clk ), .D ( signal_23380 ), .Q ( signal_23381 ) ) ;
    buf_clk cell_8696 ( .C ( clk ), .D ( signal_23388 ), .Q ( signal_23389 ) ) ;
    buf_clk cell_8704 ( .C ( clk ), .D ( signal_23396 ), .Q ( signal_23397 ) ) ;
    buf_clk cell_8712 ( .C ( clk ), .D ( signal_23404 ), .Q ( signal_23405 ) ) ;
    buf_clk cell_8724 ( .C ( clk ), .D ( signal_23416 ), .Q ( signal_23417 ) ) ;
    buf_clk cell_8736 ( .C ( clk ), .D ( signal_23428 ), .Q ( signal_23429 ) ) ;
    buf_clk cell_8748 ( .C ( clk ), .D ( signal_23440 ), .Q ( signal_23441 ) ) ;
    buf_clk cell_8760 ( .C ( clk ), .D ( signal_23452 ), .Q ( signal_23453 ) ) ;
    buf_clk cell_8772 ( .C ( clk ), .D ( signal_23464 ), .Q ( signal_23465 ) ) ;
    buf_clk cell_8778 ( .C ( clk ), .D ( signal_23470 ), .Q ( signal_23471 ) ) ;
    buf_clk cell_8784 ( .C ( clk ), .D ( signal_23476 ), .Q ( signal_23477 ) ) ;
    buf_clk cell_8790 ( .C ( clk ), .D ( signal_23482 ), .Q ( signal_23483 ) ) ;
    buf_clk cell_8796 ( .C ( clk ), .D ( signal_23488 ), .Q ( signal_23489 ) ) ;
    buf_clk cell_8802 ( .C ( clk ), .D ( signal_23494 ), .Q ( signal_23495 ) ) ;
    buf_clk cell_8808 ( .C ( clk ), .D ( signal_23500 ), .Q ( signal_23501 ) ) ;
    buf_clk cell_8814 ( .C ( clk ), .D ( signal_23506 ), .Q ( signal_23507 ) ) ;
    buf_clk cell_8820 ( .C ( clk ), .D ( signal_23512 ), .Q ( signal_23513 ) ) ;
    buf_clk cell_8826 ( .C ( clk ), .D ( signal_23518 ), .Q ( signal_23519 ) ) ;
    buf_clk cell_8832 ( .C ( clk ), .D ( signal_23524 ), .Q ( signal_23525 ) ) ;
    buf_clk cell_8846 ( .C ( clk ), .D ( signal_23538 ), .Q ( signal_23539 ) ) ;
    buf_clk cell_8860 ( .C ( clk ), .D ( signal_23552 ), .Q ( signal_23553 ) ) ;
    buf_clk cell_8874 ( .C ( clk ), .D ( signal_23566 ), .Q ( signal_23567 ) ) ;
    buf_clk cell_8888 ( .C ( clk ), .D ( signal_23580 ), .Q ( signal_23581 ) ) ;
    buf_clk cell_8902 ( .C ( clk ), .D ( signal_23594 ), .Q ( signal_23595 ) ) ;
    buf_clk cell_8910 ( .C ( clk ), .D ( signal_23602 ), .Q ( signal_23603 ) ) ;
    buf_clk cell_8918 ( .C ( clk ), .D ( signal_23610 ), .Q ( signal_23611 ) ) ;
    buf_clk cell_8926 ( .C ( clk ), .D ( signal_23618 ), .Q ( signal_23619 ) ) ;
    buf_clk cell_8934 ( .C ( clk ), .D ( signal_23626 ), .Q ( signal_23627 ) ) ;
    buf_clk cell_8942 ( .C ( clk ), .D ( signal_23634 ), .Q ( signal_23635 ) ) ;
    buf_clk cell_8956 ( .C ( clk ), .D ( signal_23648 ), .Q ( signal_23649 ) ) ;
    buf_clk cell_8970 ( .C ( clk ), .D ( signal_23662 ), .Q ( signal_23663 ) ) ;
    buf_clk cell_8984 ( .C ( clk ), .D ( signal_23676 ), .Q ( signal_23677 ) ) ;
    buf_clk cell_8998 ( .C ( clk ), .D ( signal_23690 ), .Q ( signal_23691 ) ) ;
    buf_clk cell_9012 ( .C ( clk ), .D ( signal_23704 ), .Q ( signal_23705 ) ) ;
    buf_clk cell_9020 ( .C ( clk ), .D ( signal_23712 ), .Q ( signal_23713 ) ) ;
    buf_clk cell_9028 ( .C ( clk ), .D ( signal_23720 ), .Q ( signal_23721 ) ) ;
    buf_clk cell_9036 ( .C ( clk ), .D ( signal_23728 ), .Q ( signal_23729 ) ) ;
    buf_clk cell_9044 ( .C ( clk ), .D ( signal_23736 ), .Q ( signal_23737 ) ) ;
    buf_clk cell_9052 ( .C ( clk ), .D ( signal_23744 ), .Q ( signal_23745 ) ) ;
    buf_clk cell_9080 ( .C ( clk ), .D ( signal_23772 ), .Q ( signal_23773 ) ) ;
    buf_clk cell_9090 ( .C ( clk ), .D ( signal_23782 ), .Q ( signal_23783 ) ) ;
    buf_clk cell_9100 ( .C ( clk ), .D ( signal_23792 ), .Q ( signal_23793 ) ) ;
    buf_clk cell_9110 ( .C ( clk ), .D ( signal_23802 ), .Q ( signal_23803 ) ) ;
    buf_clk cell_9120 ( .C ( clk ), .D ( signal_23812 ), .Q ( signal_23813 ) ) ;
    buf_clk cell_9156 ( .C ( clk ), .D ( signal_23848 ), .Q ( signal_23849 ) ) ;
    buf_clk cell_9172 ( .C ( clk ), .D ( signal_23864 ), .Q ( signal_23865 ) ) ;
    buf_clk cell_9188 ( .C ( clk ), .D ( signal_23880 ), .Q ( signal_23881 ) ) ;
    buf_clk cell_9204 ( .C ( clk ), .D ( signal_23896 ), .Q ( signal_23897 ) ) ;
    buf_clk cell_9220 ( .C ( clk ), .D ( signal_23912 ), .Q ( signal_23913 ) ) ;
    buf_clk cell_9256 ( .C ( clk ), .D ( signal_23948 ), .Q ( signal_23949 ) ) ;
    buf_clk cell_9272 ( .C ( clk ), .D ( signal_23964 ), .Q ( signal_23965 ) ) ;
    buf_clk cell_9288 ( .C ( clk ), .D ( signal_23980 ), .Q ( signal_23981 ) ) ;
    buf_clk cell_9304 ( .C ( clk ), .D ( signal_23996 ), .Q ( signal_23997 ) ) ;
    buf_clk cell_9320 ( .C ( clk ), .D ( signal_24012 ), .Q ( signal_24013 ) ) ;
    buf_clk cell_9330 ( .C ( clk ), .D ( signal_24022 ), .Q ( signal_24023 ) ) ;
    buf_clk cell_9340 ( .C ( clk ), .D ( signal_24032 ), .Q ( signal_24033 ) ) ;
    buf_clk cell_9350 ( .C ( clk ), .D ( signal_24042 ), .Q ( signal_24043 ) ) ;
    buf_clk cell_9360 ( .C ( clk ), .D ( signal_24052 ), .Q ( signal_24053 ) ) ;
    buf_clk cell_9370 ( .C ( clk ), .D ( signal_24062 ), .Q ( signal_24063 ) ) ;
    buf_clk cell_9428 ( .C ( clk ), .D ( signal_24120 ), .Q ( signal_24121 ) ) ;
    buf_clk cell_9438 ( .C ( clk ), .D ( signal_24130 ), .Q ( signal_24131 ) ) ;
    buf_clk cell_9448 ( .C ( clk ), .D ( signal_24140 ), .Q ( signal_24141 ) ) ;
    buf_clk cell_9458 ( .C ( clk ), .D ( signal_24150 ), .Q ( signal_24151 ) ) ;
    buf_clk cell_9468 ( .C ( clk ), .D ( signal_24160 ), .Q ( signal_24161 ) ) ;
    buf_clk cell_9508 ( .C ( clk ), .D ( signal_24200 ), .Q ( signal_24201 ) ) ;
    buf_clk cell_9518 ( .C ( clk ), .D ( signal_24210 ), .Q ( signal_24211 ) ) ;
    buf_clk cell_9528 ( .C ( clk ), .D ( signal_24220 ), .Q ( signal_24221 ) ) ;
    buf_clk cell_9538 ( .C ( clk ), .D ( signal_24230 ), .Q ( signal_24231 ) ) ;
    buf_clk cell_9548 ( .C ( clk ), .D ( signal_24240 ), .Q ( signal_24241 ) ) ;
    buf_clk cell_9564 ( .C ( clk ), .D ( signal_24256 ), .Q ( signal_24257 ) ) ;
    buf_clk cell_9580 ( .C ( clk ), .D ( signal_24272 ), .Q ( signal_24273 ) ) ;
    buf_clk cell_9596 ( .C ( clk ), .D ( signal_24288 ), .Q ( signal_24289 ) ) ;
    buf_clk cell_9612 ( .C ( clk ), .D ( signal_24304 ), .Q ( signal_24305 ) ) ;
    buf_clk cell_9628 ( .C ( clk ), .D ( signal_24320 ), .Q ( signal_24321 ) ) ;
    buf_clk cell_9646 ( .C ( clk ), .D ( signal_24338 ), .Q ( signal_24339 ) ) ;
    buf_clk cell_9664 ( .C ( clk ), .D ( signal_24356 ), .Q ( signal_24357 ) ) ;
    buf_clk cell_9682 ( .C ( clk ), .D ( signal_24374 ), .Q ( signal_24375 ) ) ;
    buf_clk cell_9700 ( .C ( clk ), .D ( signal_24392 ), .Q ( signal_24393 ) ) ;
    buf_clk cell_9718 ( .C ( clk ), .D ( signal_24410 ), .Q ( signal_24411 ) ) ;
    buf_clk cell_9746 ( .C ( clk ), .D ( signal_24438 ), .Q ( signal_24439 ) ) ;
    buf_clk cell_9754 ( .C ( clk ), .D ( signal_24446 ), .Q ( signal_24447 ) ) ;
    buf_clk cell_9762 ( .C ( clk ), .D ( signal_24454 ), .Q ( signal_24455 ) ) ;
    buf_clk cell_9770 ( .C ( clk ), .D ( signal_24462 ), .Q ( signal_24463 ) ) ;
    buf_clk cell_9778 ( .C ( clk ), .D ( signal_24470 ), .Q ( signal_24471 ) ) ;
    buf_clk cell_9896 ( .C ( clk ), .D ( signal_24588 ), .Q ( signal_24589 ) ) ;
    buf_clk cell_9916 ( .C ( clk ), .D ( signal_24608 ), .Q ( signal_24609 ) ) ;
    buf_clk cell_9936 ( .C ( clk ), .D ( signal_24628 ), .Q ( signal_24629 ) ) ;
    buf_clk cell_9956 ( .C ( clk ), .D ( signal_24648 ), .Q ( signal_24649 ) ) ;
    buf_clk cell_9976 ( .C ( clk ), .D ( signal_24668 ), .Q ( signal_24669 ) ) ;
    buf_clk cell_10026 ( .C ( clk ), .D ( signal_24718 ), .Q ( signal_24719 ) ) ;
    buf_clk cell_10038 ( .C ( clk ), .D ( signal_24730 ), .Q ( signal_24731 ) ) ;
    buf_clk cell_10050 ( .C ( clk ), .D ( signal_24742 ), .Q ( signal_24743 ) ) ;
    buf_clk cell_10062 ( .C ( clk ), .D ( signal_24754 ), .Q ( signal_24755 ) ) ;
    buf_clk cell_10074 ( .C ( clk ), .D ( signal_24766 ), .Q ( signal_24767 ) ) ;
    buf_clk cell_10086 ( .C ( clk ), .D ( signal_24778 ), .Q ( signal_24779 ) ) ;
    buf_clk cell_10100 ( .C ( clk ), .D ( signal_24792 ), .Q ( signal_24793 ) ) ;
    buf_clk cell_10114 ( .C ( clk ), .D ( signal_24806 ), .Q ( signal_24807 ) ) ;
    buf_clk cell_10128 ( .C ( clk ), .D ( signal_24820 ), .Q ( signal_24821 ) ) ;
    buf_clk cell_10142 ( .C ( clk ), .D ( signal_24834 ), .Q ( signal_24835 ) ) ;

    /* cells in depth 19 */
    buf_clk cell_8681 ( .C ( clk ), .D ( signal_23373 ), .Q ( signal_23374 ) ) ;
    buf_clk cell_8689 ( .C ( clk ), .D ( signal_23381 ), .Q ( signal_23382 ) ) ;
    buf_clk cell_8697 ( .C ( clk ), .D ( signal_23389 ), .Q ( signal_23390 ) ) ;
    buf_clk cell_8705 ( .C ( clk ), .D ( signal_23397 ), .Q ( signal_23398 ) ) ;
    buf_clk cell_8713 ( .C ( clk ), .D ( signal_23405 ), .Q ( signal_23406 ) ) ;
    buf_clk cell_8725 ( .C ( clk ), .D ( signal_23417 ), .Q ( signal_23418 ) ) ;
    buf_clk cell_8737 ( .C ( clk ), .D ( signal_23429 ), .Q ( signal_23430 ) ) ;
    buf_clk cell_8749 ( .C ( clk ), .D ( signal_23441 ), .Q ( signal_23442 ) ) ;
    buf_clk cell_8761 ( .C ( clk ), .D ( signal_23453 ), .Q ( signal_23454 ) ) ;
    buf_clk cell_8773 ( .C ( clk ), .D ( signal_23465 ), .Q ( signal_23466 ) ) ;
    buf_clk cell_8779 ( .C ( clk ), .D ( signal_23471 ), .Q ( signal_23472 ) ) ;
    buf_clk cell_8785 ( .C ( clk ), .D ( signal_23477 ), .Q ( signal_23478 ) ) ;
    buf_clk cell_8791 ( .C ( clk ), .D ( signal_23483 ), .Q ( signal_23484 ) ) ;
    buf_clk cell_8797 ( .C ( clk ), .D ( signal_23489 ), .Q ( signal_23490 ) ) ;
    buf_clk cell_8803 ( .C ( clk ), .D ( signal_23495 ), .Q ( signal_23496 ) ) ;
    buf_clk cell_8809 ( .C ( clk ), .D ( signal_23501 ), .Q ( signal_23502 ) ) ;
    buf_clk cell_8815 ( .C ( clk ), .D ( signal_23507 ), .Q ( signal_23508 ) ) ;
    buf_clk cell_8821 ( .C ( clk ), .D ( signal_23513 ), .Q ( signal_23514 ) ) ;
    buf_clk cell_8827 ( .C ( clk ), .D ( signal_23519 ), .Q ( signal_23520 ) ) ;
    buf_clk cell_8833 ( .C ( clk ), .D ( signal_23525 ), .Q ( signal_23526 ) ) ;
    buf_clk cell_8847 ( .C ( clk ), .D ( signal_23539 ), .Q ( signal_23540 ) ) ;
    buf_clk cell_8861 ( .C ( clk ), .D ( signal_23553 ), .Q ( signal_23554 ) ) ;
    buf_clk cell_8875 ( .C ( clk ), .D ( signal_23567 ), .Q ( signal_23568 ) ) ;
    buf_clk cell_8889 ( .C ( clk ), .D ( signal_23581 ), .Q ( signal_23582 ) ) ;
    buf_clk cell_8903 ( .C ( clk ), .D ( signal_23595 ), .Q ( signal_23596 ) ) ;
    buf_clk cell_8911 ( .C ( clk ), .D ( signal_23603 ), .Q ( signal_23604 ) ) ;
    buf_clk cell_8919 ( .C ( clk ), .D ( signal_23611 ), .Q ( signal_23612 ) ) ;
    buf_clk cell_8927 ( .C ( clk ), .D ( signal_23619 ), .Q ( signal_23620 ) ) ;
    buf_clk cell_8935 ( .C ( clk ), .D ( signal_23627 ), .Q ( signal_23628 ) ) ;
    buf_clk cell_8943 ( .C ( clk ), .D ( signal_23635 ), .Q ( signal_23636 ) ) ;
    buf_clk cell_8957 ( .C ( clk ), .D ( signal_23649 ), .Q ( signal_23650 ) ) ;
    buf_clk cell_8971 ( .C ( clk ), .D ( signal_23663 ), .Q ( signal_23664 ) ) ;
    buf_clk cell_8985 ( .C ( clk ), .D ( signal_23677 ), .Q ( signal_23678 ) ) ;
    buf_clk cell_8999 ( .C ( clk ), .D ( signal_23691 ), .Q ( signal_23692 ) ) ;
    buf_clk cell_9013 ( .C ( clk ), .D ( signal_23705 ), .Q ( signal_23706 ) ) ;
    buf_clk cell_9021 ( .C ( clk ), .D ( signal_23713 ), .Q ( signal_23714 ) ) ;
    buf_clk cell_9029 ( .C ( clk ), .D ( signal_23721 ), .Q ( signal_23722 ) ) ;
    buf_clk cell_9037 ( .C ( clk ), .D ( signal_23729 ), .Q ( signal_23730 ) ) ;
    buf_clk cell_9045 ( .C ( clk ), .D ( signal_23737 ), .Q ( signal_23738 ) ) ;
    buf_clk cell_9053 ( .C ( clk ), .D ( signal_23745 ), .Q ( signal_23746 ) ) ;
    buf_clk cell_9055 ( .C ( clk ), .D ( signal_2335 ), .Q ( signal_23748 ) ) ;
    buf_clk cell_9059 ( .C ( clk ), .D ( signal_7996 ), .Q ( signal_23752 ) ) ;
    buf_clk cell_9063 ( .C ( clk ), .D ( signal_7997 ), .Q ( signal_23756 ) ) ;
    buf_clk cell_9067 ( .C ( clk ), .D ( signal_7998 ), .Q ( signal_23760 ) ) ;
    buf_clk cell_9071 ( .C ( clk ), .D ( signal_7999 ), .Q ( signal_23764 ) ) ;
    buf_clk cell_9081 ( .C ( clk ), .D ( signal_23773 ), .Q ( signal_23774 ) ) ;
    buf_clk cell_9091 ( .C ( clk ), .D ( signal_23783 ), .Q ( signal_23784 ) ) ;
    buf_clk cell_9101 ( .C ( clk ), .D ( signal_23793 ), .Q ( signal_23794 ) ) ;
    buf_clk cell_9111 ( .C ( clk ), .D ( signal_23803 ), .Q ( signal_23804 ) ) ;
    buf_clk cell_9121 ( .C ( clk ), .D ( signal_23813 ), .Q ( signal_23814 ) ) ;
    buf_clk cell_9157 ( .C ( clk ), .D ( signal_23849 ), .Q ( signal_23850 ) ) ;
    buf_clk cell_9173 ( .C ( clk ), .D ( signal_23865 ), .Q ( signal_23866 ) ) ;
    buf_clk cell_9189 ( .C ( clk ), .D ( signal_23881 ), .Q ( signal_23882 ) ) ;
    buf_clk cell_9205 ( .C ( clk ), .D ( signal_23897 ), .Q ( signal_23898 ) ) ;
    buf_clk cell_9221 ( .C ( clk ), .D ( signal_23913 ), .Q ( signal_23914 ) ) ;
    buf_clk cell_9225 ( .C ( clk ), .D ( signal_2308 ), .Q ( signal_23918 ) ) ;
    buf_clk cell_9229 ( .C ( clk ), .D ( signal_7888 ), .Q ( signal_23922 ) ) ;
    buf_clk cell_9233 ( .C ( clk ), .D ( signal_7889 ), .Q ( signal_23926 ) ) ;
    buf_clk cell_9237 ( .C ( clk ), .D ( signal_7890 ), .Q ( signal_23930 ) ) ;
    buf_clk cell_9241 ( .C ( clk ), .D ( signal_7891 ), .Q ( signal_23934 ) ) ;
    buf_clk cell_9257 ( .C ( clk ), .D ( signal_23949 ), .Q ( signal_23950 ) ) ;
    buf_clk cell_9273 ( .C ( clk ), .D ( signal_23965 ), .Q ( signal_23966 ) ) ;
    buf_clk cell_9289 ( .C ( clk ), .D ( signal_23981 ), .Q ( signal_23982 ) ) ;
    buf_clk cell_9305 ( .C ( clk ), .D ( signal_23997 ), .Q ( signal_23998 ) ) ;
    buf_clk cell_9321 ( .C ( clk ), .D ( signal_24013 ), .Q ( signal_24014 ) ) ;
    buf_clk cell_9331 ( .C ( clk ), .D ( signal_24023 ), .Q ( signal_24024 ) ) ;
    buf_clk cell_9341 ( .C ( clk ), .D ( signal_24033 ), .Q ( signal_24034 ) ) ;
    buf_clk cell_9351 ( .C ( clk ), .D ( signal_24043 ), .Q ( signal_24044 ) ) ;
    buf_clk cell_9361 ( .C ( clk ), .D ( signal_24053 ), .Q ( signal_24054 ) ) ;
    buf_clk cell_9371 ( .C ( clk ), .D ( signal_24063 ), .Q ( signal_24064 ) ) ;
    buf_clk cell_9375 ( .C ( clk ), .D ( signal_2318 ), .Q ( signal_24068 ) ) ;
    buf_clk cell_9379 ( .C ( clk ), .D ( signal_7928 ), .Q ( signal_24072 ) ) ;
    buf_clk cell_9383 ( .C ( clk ), .D ( signal_7929 ), .Q ( signal_24076 ) ) ;
    buf_clk cell_9387 ( .C ( clk ), .D ( signal_7930 ), .Q ( signal_24080 ) ) ;
    buf_clk cell_9391 ( .C ( clk ), .D ( signal_7931 ), .Q ( signal_24084 ) ) ;
    buf_clk cell_9395 ( .C ( clk ), .D ( signal_2336 ), .Q ( signal_24088 ) ) ;
    buf_clk cell_9401 ( .C ( clk ), .D ( signal_8000 ), .Q ( signal_24094 ) ) ;
    buf_clk cell_9407 ( .C ( clk ), .D ( signal_8001 ), .Q ( signal_24100 ) ) ;
    buf_clk cell_9413 ( .C ( clk ), .D ( signal_8002 ), .Q ( signal_24106 ) ) ;
    buf_clk cell_9419 ( .C ( clk ), .D ( signal_8003 ), .Q ( signal_24112 ) ) ;
    buf_clk cell_9429 ( .C ( clk ), .D ( signal_24121 ), .Q ( signal_24122 ) ) ;
    buf_clk cell_9439 ( .C ( clk ), .D ( signal_24131 ), .Q ( signal_24132 ) ) ;
    buf_clk cell_9449 ( .C ( clk ), .D ( signal_24141 ), .Q ( signal_24142 ) ) ;
    buf_clk cell_9459 ( .C ( clk ), .D ( signal_24151 ), .Q ( signal_24152 ) ) ;
    buf_clk cell_9469 ( .C ( clk ), .D ( signal_24161 ), .Q ( signal_24162 ) ) ;
    buf_clk cell_9475 ( .C ( clk ), .D ( signal_2343 ), .Q ( signal_24168 ) ) ;
    buf_clk cell_9481 ( .C ( clk ), .D ( signal_8028 ), .Q ( signal_24174 ) ) ;
    buf_clk cell_9487 ( .C ( clk ), .D ( signal_8029 ), .Q ( signal_24180 ) ) ;
    buf_clk cell_9493 ( .C ( clk ), .D ( signal_8030 ), .Q ( signal_24186 ) ) ;
    buf_clk cell_9499 ( .C ( clk ), .D ( signal_8031 ), .Q ( signal_24192 ) ) ;
    buf_clk cell_9509 ( .C ( clk ), .D ( signal_24201 ), .Q ( signal_24202 ) ) ;
    buf_clk cell_9519 ( .C ( clk ), .D ( signal_24211 ), .Q ( signal_24212 ) ) ;
    buf_clk cell_9529 ( .C ( clk ), .D ( signal_24221 ), .Q ( signal_24222 ) ) ;
    buf_clk cell_9539 ( .C ( clk ), .D ( signal_24231 ), .Q ( signal_24232 ) ) ;
    buf_clk cell_9549 ( .C ( clk ), .D ( signal_24241 ), .Q ( signal_24242 ) ) ;
    buf_clk cell_9565 ( .C ( clk ), .D ( signal_24257 ), .Q ( signal_24258 ) ) ;
    buf_clk cell_9581 ( .C ( clk ), .D ( signal_24273 ), .Q ( signal_24274 ) ) ;
    buf_clk cell_9597 ( .C ( clk ), .D ( signal_24289 ), .Q ( signal_24290 ) ) ;
    buf_clk cell_9613 ( .C ( clk ), .D ( signal_24305 ), .Q ( signal_24306 ) ) ;
    buf_clk cell_9629 ( .C ( clk ), .D ( signal_24321 ), .Q ( signal_24322 ) ) ;
    buf_clk cell_9647 ( .C ( clk ), .D ( signal_24339 ), .Q ( signal_24340 ) ) ;
    buf_clk cell_9665 ( .C ( clk ), .D ( signal_24357 ), .Q ( signal_24358 ) ) ;
    buf_clk cell_9683 ( .C ( clk ), .D ( signal_24375 ), .Q ( signal_24376 ) ) ;
    buf_clk cell_9701 ( .C ( clk ), .D ( signal_24393 ), .Q ( signal_24394 ) ) ;
    buf_clk cell_9719 ( .C ( clk ), .D ( signal_24411 ), .Q ( signal_24412 ) ) ;
    buf_clk cell_9747 ( .C ( clk ), .D ( signal_24439 ), .Q ( signal_24440 ) ) ;
    buf_clk cell_9755 ( .C ( clk ), .D ( signal_24447 ), .Q ( signal_24448 ) ) ;
    buf_clk cell_9763 ( .C ( clk ), .D ( signal_24455 ), .Q ( signal_24456 ) ) ;
    buf_clk cell_9771 ( .C ( clk ), .D ( signal_24463 ), .Q ( signal_24464 ) ) ;
    buf_clk cell_9779 ( .C ( clk ), .D ( signal_24471 ), .Q ( signal_24472 ) ) ;
    buf_clk cell_9785 ( .C ( clk ), .D ( signal_2306 ), .Q ( signal_24478 ) ) ;
    buf_clk cell_9793 ( .C ( clk ), .D ( signal_7880 ), .Q ( signal_24486 ) ) ;
    buf_clk cell_9801 ( .C ( clk ), .D ( signal_7881 ), .Q ( signal_24494 ) ) ;
    buf_clk cell_9809 ( .C ( clk ), .D ( signal_7882 ), .Q ( signal_24502 ) ) ;
    buf_clk cell_9817 ( .C ( clk ), .D ( signal_7883 ), .Q ( signal_24510 ) ) ;
    buf_clk cell_9897 ( .C ( clk ), .D ( signal_24589 ), .Q ( signal_24590 ) ) ;
    buf_clk cell_9917 ( .C ( clk ), .D ( signal_24609 ), .Q ( signal_24610 ) ) ;
    buf_clk cell_9937 ( .C ( clk ), .D ( signal_24629 ), .Q ( signal_24630 ) ) ;
    buf_clk cell_9957 ( .C ( clk ), .D ( signal_24649 ), .Q ( signal_24650 ) ) ;
    buf_clk cell_9977 ( .C ( clk ), .D ( signal_24669 ), .Q ( signal_24670 ) ) ;
    buf_clk cell_10027 ( .C ( clk ), .D ( signal_24719 ), .Q ( signal_24720 ) ) ;
    buf_clk cell_10039 ( .C ( clk ), .D ( signal_24731 ), .Q ( signal_24732 ) ) ;
    buf_clk cell_10051 ( .C ( clk ), .D ( signal_24743 ), .Q ( signal_24744 ) ) ;
    buf_clk cell_10063 ( .C ( clk ), .D ( signal_24755 ), .Q ( signal_24756 ) ) ;
    buf_clk cell_10075 ( .C ( clk ), .D ( signal_24767 ), .Q ( signal_24768 ) ) ;
    buf_clk cell_10087 ( .C ( clk ), .D ( signal_24779 ), .Q ( signal_24780 ) ) ;
    buf_clk cell_10101 ( .C ( clk ), .D ( signal_24793 ), .Q ( signal_24794 ) ) ;
    buf_clk cell_10115 ( .C ( clk ), .D ( signal_24807 ), .Q ( signal_24808 ) ) ;
    buf_clk cell_10129 ( .C ( clk ), .D ( signal_24821 ), .Q ( signal_24822 ) ) ;
    buf_clk cell_10143 ( .C ( clk ), .D ( signal_24835 ), .Q ( signal_24836 ) ) ;
    buf_clk cell_10155 ( .C ( clk ), .D ( signal_2328 ), .Q ( signal_24848 ) ) ;
    buf_clk cell_10169 ( .C ( clk ), .D ( signal_7968 ), .Q ( signal_24862 ) ) ;
    buf_clk cell_10183 ( .C ( clk ), .D ( signal_7969 ), .Q ( signal_24876 ) ) ;
    buf_clk cell_10197 ( .C ( clk ), .D ( signal_7970 ), .Q ( signal_24890 ) ) ;
    buf_clk cell_10211 ( .C ( clk ), .D ( signal_7971 ), .Q ( signal_24904 ) ) ;

    /* cells in depth 20 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2269 ( .a ({signal_22897, signal_22891, signal_22885, signal_22879, signal_22873}), .b ({signal_7639, signal_7638, signal_7637, signal_7636, signal_2245}), .clk ( clk ), .r ({Fresh[8269], Fresh[8268], Fresh[8267], Fresh[8266], Fresh[8265], Fresh[8264], Fresh[8263], Fresh[8262], Fresh[8261], Fresh[8260]}), .c ({signal_7795, signal_7794, signal_7793, signal_7792, signal_2284}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2270 ( .a ({signal_22937, signal_22929, signal_22921, signal_22913, signal_22905}), .b ({signal_7647, signal_7646, signal_7645, signal_7644, signal_2247}), .clk ( clk ), .r ({Fresh[8279], Fresh[8278], Fresh[8277], Fresh[8276], Fresh[8275], Fresh[8274], Fresh[8273], Fresh[8272], Fresh[8271], Fresh[8270]}), .c ({signal_7799, signal_7798, signal_7797, signal_7796, signal_2285}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2296 ( .a ({signal_22967, signal_22961, signal_22955, signal_22949, signal_22943}), .b ({signal_7787, signal_7786, signal_7785, signal_7784, signal_2282}), .clk ( clk ), .r ({Fresh[8289], Fresh[8288], Fresh[8287], Fresh[8286], Fresh[8285], Fresh[8284], Fresh[8283], Fresh[8282], Fresh[8281], Fresh[8280]}), .c ({signal_7903, signal_7902, signal_7901, signal_7900, signal_2311}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2316 ( .a ({signal_23017, signal_23007, signal_22997, signal_22987, signal_22977}), .b ({signal_7887, signal_7886, signal_7885, signal_7884, signal_2307}), .clk ( clk ), .r ({Fresh[8299], Fresh[8298], Fresh[8297], Fresh[8296], Fresh[8295], Fresh[8294], Fresh[8293], Fresh[8292], Fresh[8291], Fresh[8290]}), .c ({signal_7983, signal_7982, signal_7981, signal_7980, signal_2331}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2317 ( .a ({signal_23047, signal_23041, signal_23035, signal_23029, signal_23023}), .b ({signal_7843, signal_7842, signal_7841, signal_7840, signal_2296}), .clk ( clk ), .r ({Fresh[8309], Fresh[8308], Fresh[8307], Fresh[8306], Fresh[8305], Fresh[8304], Fresh[8303], Fresh[8302], Fresh[8301], Fresh[8300]}), .c ({signal_7987, signal_7986, signal_7985, signal_7984, signal_2332}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2318 ( .a ({signal_23067, signal_23063, signal_23059, signal_23055, signal_23051}), .b ({signal_7643, signal_7642, signal_7641, signal_7640, signal_2246}), .clk ( clk ), .r ({Fresh[8319], Fresh[8318], Fresh[8317], Fresh[8316], Fresh[8315], Fresh[8314], Fresh[8313], Fresh[8312], Fresh[8311], Fresh[8310]}), .c ({signal_7991, signal_7990, signal_7989, signal_7988, signal_2333}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2325 ( .a ({signal_23107, signal_23099, signal_23091, signal_23083, signal_23075}), .b ({signal_7911, signal_7910, signal_7909, signal_7908, signal_2313}), .clk ( clk ), .r ({Fresh[8329], Fresh[8328], Fresh[8327], Fresh[8326], Fresh[8325], Fresh[8324], Fresh[8323], Fresh[8322], Fresh[8321], Fresh[8320]}), .c ({signal_8019, signal_8018, signal_8017, signal_8016, signal_2340}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2327 ( .a ({signal_23137, signal_23131, signal_23125, signal_23119, signal_23113}), .b ({signal_7919, signal_7918, signal_7917, signal_7916, signal_2315}), .clk ( clk ), .r ({Fresh[8339], Fresh[8338], Fresh[8337], Fresh[8336], Fresh[8335], Fresh[8334], Fresh[8333], Fresh[8332], Fresh[8331], Fresh[8330]}), .c ({signal_8027, signal_8026, signal_8025, signal_8024, signal_2342}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2331 ( .a ({signal_23177, signal_23169, signal_23161, signal_23153, signal_23145}), .b ({signal_7967, signal_7966, signal_7965, signal_7964, signal_2327}), .clk ( clk ), .r ({Fresh[8349], Fresh[8348], Fresh[8347], Fresh[8346], Fresh[8345], Fresh[8344], Fresh[8343], Fresh[8342], Fresh[8341], Fresh[8340]}), .c ({signal_8043, signal_8042, signal_8041, signal_8040, signal_2346}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2332 ( .a ({signal_23207, signal_23201, signal_23195, signal_23189, signal_23183}), .b ({signal_7927, signal_7926, signal_7925, signal_7924, signal_2317}), .clk ( clk ), .r ({Fresh[8359], Fresh[8358], Fresh[8357], Fresh[8356], Fresh[8355], Fresh[8354], Fresh[8353], Fresh[8352], Fresh[8351], Fresh[8350]}), .c ({signal_8047, signal_8046, signal_8045, signal_8044, signal_2347}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2333 ( .a ({signal_23247, signal_23239, signal_23231, signal_23223, signal_23215}), .b ({signal_7975, signal_7974, signal_7973, signal_7972, signal_2329}), .clk ( clk ), .r ({Fresh[8369], Fresh[8368], Fresh[8367], Fresh[8366], Fresh[8365], Fresh[8364], Fresh[8363], Fresh[8362], Fresh[8361], Fresh[8360]}), .c ({signal_8051, signal_8050, signal_8049, signal_8048, signal_2348}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2335 ( .a ({signal_8019, signal_8018, signal_8017, signal_8016, signal_2340}), .b ({signal_8059, signal_8058, signal_8057, signal_8056, signal_2350}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2336 ( .a ({signal_8047, signal_8046, signal_8045, signal_8044, signal_2347}), .b ({signal_8063, signal_8062, signal_8061, signal_8060, signal_2351}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2337 ( .a ({signal_23267, signal_23263, signal_23259, signal_23255, signal_23251}), .b ({signal_8023, signal_8022, signal_8021, signal_8020, signal_2341}), .clk ( clk ), .r ({Fresh[8379], Fresh[8378], Fresh[8377], Fresh[8376], Fresh[8375], Fresh[8374], Fresh[8373], Fresh[8372], Fresh[8371], Fresh[8370]}), .c ({signal_8067, signal_8066, signal_8065, signal_8064, signal_2352}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2339 ( .a ({signal_23297, signal_23291, signal_23285, signal_23279, signal_23273}), .b ({signal_8035, signal_8034, signal_8033, signal_8032, signal_2344}), .clk ( clk ), .r ({Fresh[8389], Fresh[8388], Fresh[8387], Fresh[8386], Fresh[8385], Fresh[8384], Fresh[8383], Fresh[8382], Fresh[8381], Fresh[8380]}), .c ({signal_8075, signal_8074, signal_8073, signal_8072, signal_2354}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2340 ( .a ({signal_23327, signal_23321, signal_23315, signal_23309, signal_23303}), .b ({signal_8007, signal_8006, signal_8005, signal_8004, signal_2337}), .clk ( clk ), .r ({Fresh[8399], Fresh[8398], Fresh[8397], Fresh[8396], Fresh[8395], Fresh[8394], Fresh[8393], Fresh[8392], Fresh[8391], Fresh[8390]}), .c ({signal_8079, signal_8078, signal_8077, signal_8076, signal_2355}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2341 ( .a ({signal_23347, signal_23343, signal_23339, signal_23335, signal_23331}), .b ({signal_8011, signal_8010, signal_8009, signal_8008, signal_2338}), .clk ( clk ), .r ({Fresh[8409], Fresh[8408], Fresh[8407], Fresh[8406], Fresh[8405], Fresh[8404], Fresh[8403], Fresh[8402], Fresh[8401], Fresh[8400]}), .c ({signal_8083, signal_8082, signal_8081, signal_8080, signal_2356}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2342 ( .a ({signal_23367, signal_23363, signal_23359, signal_23355, signal_23351}), .b ({signal_8039, signal_8038, signal_8037, signal_8036, signal_2345}), .clk ( clk ), .r ({Fresh[8419], Fresh[8418], Fresh[8417], Fresh[8416], Fresh[8415], Fresh[8414], Fresh[8413], Fresh[8412], Fresh[8411], Fresh[8410]}), .c ({signal_8087, signal_8086, signal_8085, signal_8084, signal_2357}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2343 ( .a ({signal_8015, signal_8014, signal_8013, signal_8012, signal_2339}), .b ({signal_7979, signal_7978, signal_7977, signal_7976, signal_2330}), .clk ( clk ), .r ({Fresh[8429], Fresh[8428], Fresh[8427], Fresh[8426], Fresh[8425], Fresh[8424], Fresh[8423], Fresh[8422], Fresh[8421], Fresh[8420]}), .c ({signal_8091, signal_8090, signal_8089, signal_8088, signal_2358}) ) ;
    buf_clk cell_8682 ( .C ( clk ), .D ( signal_23374 ), .Q ( signal_23375 ) ) ;
    buf_clk cell_8690 ( .C ( clk ), .D ( signal_23382 ), .Q ( signal_23383 ) ) ;
    buf_clk cell_8698 ( .C ( clk ), .D ( signal_23390 ), .Q ( signal_23391 ) ) ;
    buf_clk cell_8706 ( .C ( clk ), .D ( signal_23398 ), .Q ( signal_23399 ) ) ;
    buf_clk cell_8714 ( .C ( clk ), .D ( signal_23406 ), .Q ( signal_23407 ) ) ;
    buf_clk cell_8726 ( .C ( clk ), .D ( signal_23418 ), .Q ( signal_23419 ) ) ;
    buf_clk cell_8738 ( .C ( clk ), .D ( signal_23430 ), .Q ( signal_23431 ) ) ;
    buf_clk cell_8750 ( .C ( clk ), .D ( signal_23442 ), .Q ( signal_23443 ) ) ;
    buf_clk cell_8762 ( .C ( clk ), .D ( signal_23454 ), .Q ( signal_23455 ) ) ;
    buf_clk cell_8774 ( .C ( clk ), .D ( signal_23466 ), .Q ( signal_23467 ) ) ;
    buf_clk cell_8780 ( .C ( clk ), .D ( signal_23472 ), .Q ( signal_23473 ) ) ;
    buf_clk cell_8786 ( .C ( clk ), .D ( signal_23478 ), .Q ( signal_23479 ) ) ;
    buf_clk cell_8792 ( .C ( clk ), .D ( signal_23484 ), .Q ( signal_23485 ) ) ;
    buf_clk cell_8798 ( .C ( clk ), .D ( signal_23490 ), .Q ( signal_23491 ) ) ;
    buf_clk cell_8804 ( .C ( clk ), .D ( signal_23496 ), .Q ( signal_23497 ) ) ;
    buf_clk cell_8810 ( .C ( clk ), .D ( signal_23502 ), .Q ( signal_23503 ) ) ;
    buf_clk cell_8816 ( .C ( clk ), .D ( signal_23508 ), .Q ( signal_23509 ) ) ;
    buf_clk cell_8822 ( .C ( clk ), .D ( signal_23514 ), .Q ( signal_23515 ) ) ;
    buf_clk cell_8828 ( .C ( clk ), .D ( signal_23520 ), .Q ( signal_23521 ) ) ;
    buf_clk cell_8834 ( .C ( clk ), .D ( signal_23526 ), .Q ( signal_23527 ) ) ;
    buf_clk cell_8848 ( .C ( clk ), .D ( signal_23540 ), .Q ( signal_23541 ) ) ;
    buf_clk cell_8862 ( .C ( clk ), .D ( signal_23554 ), .Q ( signal_23555 ) ) ;
    buf_clk cell_8876 ( .C ( clk ), .D ( signal_23568 ), .Q ( signal_23569 ) ) ;
    buf_clk cell_8890 ( .C ( clk ), .D ( signal_23582 ), .Q ( signal_23583 ) ) ;
    buf_clk cell_8904 ( .C ( clk ), .D ( signal_23596 ), .Q ( signal_23597 ) ) ;
    buf_clk cell_8912 ( .C ( clk ), .D ( signal_23604 ), .Q ( signal_23605 ) ) ;
    buf_clk cell_8920 ( .C ( clk ), .D ( signal_23612 ), .Q ( signal_23613 ) ) ;
    buf_clk cell_8928 ( .C ( clk ), .D ( signal_23620 ), .Q ( signal_23621 ) ) ;
    buf_clk cell_8936 ( .C ( clk ), .D ( signal_23628 ), .Q ( signal_23629 ) ) ;
    buf_clk cell_8944 ( .C ( clk ), .D ( signal_23636 ), .Q ( signal_23637 ) ) ;
    buf_clk cell_8958 ( .C ( clk ), .D ( signal_23650 ), .Q ( signal_23651 ) ) ;
    buf_clk cell_8972 ( .C ( clk ), .D ( signal_23664 ), .Q ( signal_23665 ) ) ;
    buf_clk cell_8986 ( .C ( clk ), .D ( signal_23678 ), .Q ( signal_23679 ) ) ;
    buf_clk cell_9000 ( .C ( clk ), .D ( signal_23692 ), .Q ( signal_23693 ) ) ;
    buf_clk cell_9014 ( .C ( clk ), .D ( signal_23706 ), .Q ( signal_23707 ) ) ;
    buf_clk cell_9022 ( .C ( clk ), .D ( signal_23714 ), .Q ( signal_23715 ) ) ;
    buf_clk cell_9030 ( .C ( clk ), .D ( signal_23722 ), .Q ( signal_23723 ) ) ;
    buf_clk cell_9038 ( .C ( clk ), .D ( signal_23730 ), .Q ( signal_23731 ) ) ;
    buf_clk cell_9046 ( .C ( clk ), .D ( signal_23738 ), .Q ( signal_23739 ) ) ;
    buf_clk cell_9054 ( .C ( clk ), .D ( signal_23746 ), .Q ( signal_23747 ) ) ;
    buf_clk cell_9056 ( .C ( clk ), .D ( signal_23748 ), .Q ( signal_23749 ) ) ;
    buf_clk cell_9060 ( .C ( clk ), .D ( signal_23752 ), .Q ( signal_23753 ) ) ;
    buf_clk cell_9064 ( .C ( clk ), .D ( signal_23756 ), .Q ( signal_23757 ) ) ;
    buf_clk cell_9068 ( .C ( clk ), .D ( signal_23760 ), .Q ( signal_23761 ) ) ;
    buf_clk cell_9072 ( .C ( clk ), .D ( signal_23764 ), .Q ( signal_23765 ) ) ;
    buf_clk cell_9082 ( .C ( clk ), .D ( signal_23774 ), .Q ( signal_23775 ) ) ;
    buf_clk cell_9092 ( .C ( clk ), .D ( signal_23784 ), .Q ( signal_23785 ) ) ;
    buf_clk cell_9102 ( .C ( clk ), .D ( signal_23794 ), .Q ( signal_23795 ) ) ;
    buf_clk cell_9112 ( .C ( clk ), .D ( signal_23804 ), .Q ( signal_23805 ) ) ;
    buf_clk cell_9122 ( .C ( clk ), .D ( signal_23814 ), .Q ( signal_23815 ) ) ;
    buf_clk cell_9158 ( .C ( clk ), .D ( signal_23850 ), .Q ( signal_23851 ) ) ;
    buf_clk cell_9174 ( .C ( clk ), .D ( signal_23866 ), .Q ( signal_23867 ) ) ;
    buf_clk cell_9190 ( .C ( clk ), .D ( signal_23882 ), .Q ( signal_23883 ) ) ;
    buf_clk cell_9206 ( .C ( clk ), .D ( signal_23898 ), .Q ( signal_23899 ) ) ;
    buf_clk cell_9222 ( .C ( clk ), .D ( signal_23914 ), .Q ( signal_23915 ) ) ;
    buf_clk cell_9226 ( .C ( clk ), .D ( signal_23918 ), .Q ( signal_23919 ) ) ;
    buf_clk cell_9230 ( .C ( clk ), .D ( signal_23922 ), .Q ( signal_23923 ) ) ;
    buf_clk cell_9234 ( .C ( clk ), .D ( signal_23926 ), .Q ( signal_23927 ) ) ;
    buf_clk cell_9238 ( .C ( clk ), .D ( signal_23930 ), .Q ( signal_23931 ) ) ;
    buf_clk cell_9242 ( .C ( clk ), .D ( signal_23934 ), .Q ( signal_23935 ) ) ;
    buf_clk cell_9258 ( .C ( clk ), .D ( signal_23950 ), .Q ( signal_23951 ) ) ;
    buf_clk cell_9274 ( .C ( clk ), .D ( signal_23966 ), .Q ( signal_23967 ) ) ;
    buf_clk cell_9290 ( .C ( clk ), .D ( signal_23982 ), .Q ( signal_23983 ) ) ;
    buf_clk cell_9306 ( .C ( clk ), .D ( signal_23998 ), .Q ( signal_23999 ) ) ;
    buf_clk cell_9322 ( .C ( clk ), .D ( signal_24014 ), .Q ( signal_24015 ) ) ;
    buf_clk cell_9332 ( .C ( clk ), .D ( signal_24024 ), .Q ( signal_24025 ) ) ;
    buf_clk cell_9342 ( .C ( clk ), .D ( signal_24034 ), .Q ( signal_24035 ) ) ;
    buf_clk cell_9352 ( .C ( clk ), .D ( signal_24044 ), .Q ( signal_24045 ) ) ;
    buf_clk cell_9362 ( .C ( clk ), .D ( signal_24054 ), .Q ( signal_24055 ) ) ;
    buf_clk cell_9372 ( .C ( clk ), .D ( signal_24064 ), .Q ( signal_24065 ) ) ;
    buf_clk cell_9376 ( .C ( clk ), .D ( signal_24068 ), .Q ( signal_24069 ) ) ;
    buf_clk cell_9380 ( .C ( clk ), .D ( signal_24072 ), .Q ( signal_24073 ) ) ;
    buf_clk cell_9384 ( .C ( clk ), .D ( signal_24076 ), .Q ( signal_24077 ) ) ;
    buf_clk cell_9388 ( .C ( clk ), .D ( signal_24080 ), .Q ( signal_24081 ) ) ;
    buf_clk cell_9392 ( .C ( clk ), .D ( signal_24084 ), .Q ( signal_24085 ) ) ;
    buf_clk cell_9396 ( .C ( clk ), .D ( signal_24088 ), .Q ( signal_24089 ) ) ;
    buf_clk cell_9402 ( .C ( clk ), .D ( signal_24094 ), .Q ( signal_24095 ) ) ;
    buf_clk cell_9408 ( .C ( clk ), .D ( signal_24100 ), .Q ( signal_24101 ) ) ;
    buf_clk cell_9414 ( .C ( clk ), .D ( signal_24106 ), .Q ( signal_24107 ) ) ;
    buf_clk cell_9420 ( .C ( clk ), .D ( signal_24112 ), .Q ( signal_24113 ) ) ;
    buf_clk cell_9430 ( .C ( clk ), .D ( signal_24122 ), .Q ( signal_24123 ) ) ;
    buf_clk cell_9440 ( .C ( clk ), .D ( signal_24132 ), .Q ( signal_24133 ) ) ;
    buf_clk cell_9450 ( .C ( clk ), .D ( signal_24142 ), .Q ( signal_24143 ) ) ;
    buf_clk cell_9460 ( .C ( clk ), .D ( signal_24152 ), .Q ( signal_24153 ) ) ;
    buf_clk cell_9470 ( .C ( clk ), .D ( signal_24162 ), .Q ( signal_24163 ) ) ;
    buf_clk cell_9476 ( .C ( clk ), .D ( signal_24168 ), .Q ( signal_24169 ) ) ;
    buf_clk cell_9482 ( .C ( clk ), .D ( signal_24174 ), .Q ( signal_24175 ) ) ;
    buf_clk cell_9488 ( .C ( clk ), .D ( signal_24180 ), .Q ( signal_24181 ) ) ;
    buf_clk cell_9494 ( .C ( clk ), .D ( signal_24186 ), .Q ( signal_24187 ) ) ;
    buf_clk cell_9500 ( .C ( clk ), .D ( signal_24192 ), .Q ( signal_24193 ) ) ;
    buf_clk cell_9510 ( .C ( clk ), .D ( signal_24202 ), .Q ( signal_24203 ) ) ;
    buf_clk cell_9520 ( .C ( clk ), .D ( signal_24212 ), .Q ( signal_24213 ) ) ;
    buf_clk cell_9530 ( .C ( clk ), .D ( signal_24222 ), .Q ( signal_24223 ) ) ;
    buf_clk cell_9540 ( .C ( clk ), .D ( signal_24232 ), .Q ( signal_24233 ) ) ;
    buf_clk cell_9550 ( .C ( clk ), .D ( signal_24242 ), .Q ( signal_24243 ) ) ;
    buf_clk cell_9566 ( .C ( clk ), .D ( signal_24258 ), .Q ( signal_24259 ) ) ;
    buf_clk cell_9582 ( .C ( clk ), .D ( signal_24274 ), .Q ( signal_24275 ) ) ;
    buf_clk cell_9598 ( .C ( clk ), .D ( signal_24290 ), .Q ( signal_24291 ) ) ;
    buf_clk cell_9614 ( .C ( clk ), .D ( signal_24306 ), .Q ( signal_24307 ) ) ;
    buf_clk cell_9630 ( .C ( clk ), .D ( signal_24322 ), .Q ( signal_24323 ) ) ;
    buf_clk cell_9648 ( .C ( clk ), .D ( signal_24340 ), .Q ( signal_24341 ) ) ;
    buf_clk cell_9666 ( .C ( clk ), .D ( signal_24358 ), .Q ( signal_24359 ) ) ;
    buf_clk cell_9684 ( .C ( clk ), .D ( signal_24376 ), .Q ( signal_24377 ) ) ;
    buf_clk cell_9702 ( .C ( clk ), .D ( signal_24394 ), .Q ( signal_24395 ) ) ;
    buf_clk cell_9720 ( .C ( clk ), .D ( signal_24412 ), .Q ( signal_24413 ) ) ;
    buf_clk cell_9748 ( .C ( clk ), .D ( signal_24440 ), .Q ( signal_24441 ) ) ;
    buf_clk cell_9756 ( .C ( clk ), .D ( signal_24448 ), .Q ( signal_24449 ) ) ;
    buf_clk cell_9764 ( .C ( clk ), .D ( signal_24456 ), .Q ( signal_24457 ) ) ;
    buf_clk cell_9772 ( .C ( clk ), .D ( signal_24464 ), .Q ( signal_24465 ) ) ;
    buf_clk cell_9780 ( .C ( clk ), .D ( signal_24472 ), .Q ( signal_24473 ) ) ;
    buf_clk cell_9786 ( .C ( clk ), .D ( signal_24478 ), .Q ( signal_24479 ) ) ;
    buf_clk cell_9794 ( .C ( clk ), .D ( signal_24486 ), .Q ( signal_24487 ) ) ;
    buf_clk cell_9802 ( .C ( clk ), .D ( signal_24494 ), .Q ( signal_24495 ) ) ;
    buf_clk cell_9810 ( .C ( clk ), .D ( signal_24502 ), .Q ( signal_24503 ) ) ;
    buf_clk cell_9818 ( .C ( clk ), .D ( signal_24510 ), .Q ( signal_24511 ) ) ;
    buf_clk cell_9898 ( .C ( clk ), .D ( signal_24590 ), .Q ( signal_24591 ) ) ;
    buf_clk cell_9918 ( .C ( clk ), .D ( signal_24610 ), .Q ( signal_24611 ) ) ;
    buf_clk cell_9938 ( .C ( clk ), .D ( signal_24630 ), .Q ( signal_24631 ) ) ;
    buf_clk cell_9958 ( .C ( clk ), .D ( signal_24650 ), .Q ( signal_24651 ) ) ;
    buf_clk cell_9978 ( .C ( clk ), .D ( signal_24670 ), .Q ( signal_24671 ) ) ;
    buf_clk cell_10028 ( .C ( clk ), .D ( signal_24720 ), .Q ( signal_24721 ) ) ;
    buf_clk cell_10040 ( .C ( clk ), .D ( signal_24732 ), .Q ( signal_24733 ) ) ;
    buf_clk cell_10052 ( .C ( clk ), .D ( signal_24744 ), .Q ( signal_24745 ) ) ;
    buf_clk cell_10064 ( .C ( clk ), .D ( signal_24756 ), .Q ( signal_24757 ) ) ;
    buf_clk cell_10076 ( .C ( clk ), .D ( signal_24768 ), .Q ( signal_24769 ) ) ;
    buf_clk cell_10088 ( .C ( clk ), .D ( signal_24780 ), .Q ( signal_24781 ) ) ;
    buf_clk cell_10102 ( .C ( clk ), .D ( signal_24794 ), .Q ( signal_24795 ) ) ;
    buf_clk cell_10116 ( .C ( clk ), .D ( signal_24808 ), .Q ( signal_24809 ) ) ;
    buf_clk cell_10130 ( .C ( clk ), .D ( signal_24822 ), .Q ( signal_24823 ) ) ;
    buf_clk cell_10144 ( .C ( clk ), .D ( signal_24836 ), .Q ( signal_24837 ) ) ;
    buf_clk cell_10156 ( .C ( clk ), .D ( signal_24848 ), .Q ( signal_24849 ) ) ;
    buf_clk cell_10170 ( .C ( clk ), .D ( signal_24862 ), .Q ( signal_24863 ) ) ;
    buf_clk cell_10184 ( .C ( clk ), .D ( signal_24876 ), .Q ( signal_24877 ) ) ;
    buf_clk cell_10198 ( .C ( clk ), .D ( signal_24890 ), .Q ( signal_24891 ) ) ;
    buf_clk cell_10212 ( .C ( clk ), .D ( signal_24904 ), .Q ( signal_24905 ) ) ;

    /* cells in depth 21 */
    buf_clk cell_9057 ( .C ( clk ), .D ( signal_23749 ), .Q ( signal_23750 ) ) ;
    buf_clk cell_9061 ( .C ( clk ), .D ( signal_23753 ), .Q ( signal_23754 ) ) ;
    buf_clk cell_9065 ( .C ( clk ), .D ( signal_23757 ), .Q ( signal_23758 ) ) ;
    buf_clk cell_9069 ( .C ( clk ), .D ( signal_23761 ), .Q ( signal_23762 ) ) ;
    buf_clk cell_9073 ( .C ( clk ), .D ( signal_23765 ), .Q ( signal_23766 ) ) ;
    buf_clk cell_9083 ( .C ( clk ), .D ( signal_23775 ), .Q ( signal_23776 ) ) ;
    buf_clk cell_9093 ( .C ( clk ), .D ( signal_23785 ), .Q ( signal_23786 ) ) ;
    buf_clk cell_9103 ( .C ( clk ), .D ( signal_23795 ), .Q ( signal_23796 ) ) ;
    buf_clk cell_9113 ( .C ( clk ), .D ( signal_23805 ), .Q ( signal_23806 ) ) ;
    buf_clk cell_9123 ( .C ( clk ), .D ( signal_23815 ), .Q ( signal_23816 ) ) ;
    buf_clk cell_9125 ( .C ( clk ), .D ( signal_2354 ), .Q ( signal_23818 ) ) ;
    buf_clk cell_9127 ( .C ( clk ), .D ( signal_8072 ), .Q ( signal_23820 ) ) ;
    buf_clk cell_9129 ( .C ( clk ), .D ( signal_8073 ), .Q ( signal_23822 ) ) ;
    buf_clk cell_9131 ( .C ( clk ), .D ( signal_8074 ), .Q ( signal_23824 ) ) ;
    buf_clk cell_9133 ( .C ( clk ), .D ( signal_8075 ), .Q ( signal_23826 ) ) ;
    buf_clk cell_9135 ( .C ( clk ), .D ( signal_2357 ), .Q ( signal_23828 ) ) ;
    buf_clk cell_9137 ( .C ( clk ), .D ( signal_8084 ), .Q ( signal_23830 ) ) ;
    buf_clk cell_9139 ( .C ( clk ), .D ( signal_8085 ), .Q ( signal_23832 ) ) ;
    buf_clk cell_9141 ( .C ( clk ), .D ( signal_8086 ), .Q ( signal_23834 ) ) ;
    buf_clk cell_9143 ( .C ( clk ), .D ( signal_8087 ), .Q ( signal_23836 ) ) ;
    buf_clk cell_9159 ( .C ( clk ), .D ( signal_23851 ), .Q ( signal_23852 ) ) ;
    buf_clk cell_9175 ( .C ( clk ), .D ( signal_23867 ), .Q ( signal_23868 ) ) ;
    buf_clk cell_9191 ( .C ( clk ), .D ( signal_23883 ), .Q ( signal_23884 ) ) ;
    buf_clk cell_9207 ( .C ( clk ), .D ( signal_23899 ), .Q ( signal_23900 ) ) ;
    buf_clk cell_9223 ( .C ( clk ), .D ( signal_23915 ), .Q ( signal_23916 ) ) ;
    buf_clk cell_9227 ( .C ( clk ), .D ( signal_23919 ), .Q ( signal_23920 ) ) ;
    buf_clk cell_9231 ( .C ( clk ), .D ( signal_23923 ), .Q ( signal_23924 ) ) ;
    buf_clk cell_9235 ( .C ( clk ), .D ( signal_23927 ), .Q ( signal_23928 ) ) ;
    buf_clk cell_9239 ( .C ( clk ), .D ( signal_23931 ), .Q ( signal_23932 ) ) ;
    buf_clk cell_9243 ( .C ( clk ), .D ( signal_23935 ), .Q ( signal_23936 ) ) ;
    buf_clk cell_9259 ( .C ( clk ), .D ( signal_23951 ), .Q ( signal_23952 ) ) ;
    buf_clk cell_9275 ( .C ( clk ), .D ( signal_23967 ), .Q ( signal_23968 ) ) ;
    buf_clk cell_9291 ( .C ( clk ), .D ( signal_23983 ), .Q ( signal_23984 ) ) ;
    buf_clk cell_9307 ( .C ( clk ), .D ( signal_23999 ), .Q ( signal_24000 ) ) ;
    buf_clk cell_9323 ( .C ( clk ), .D ( signal_24015 ), .Q ( signal_24016 ) ) ;
    buf_clk cell_9333 ( .C ( clk ), .D ( signal_24025 ), .Q ( signal_24026 ) ) ;
    buf_clk cell_9343 ( .C ( clk ), .D ( signal_24035 ), .Q ( signal_24036 ) ) ;
    buf_clk cell_9353 ( .C ( clk ), .D ( signal_24045 ), .Q ( signal_24046 ) ) ;
    buf_clk cell_9363 ( .C ( clk ), .D ( signal_24055 ), .Q ( signal_24056 ) ) ;
    buf_clk cell_9373 ( .C ( clk ), .D ( signal_24065 ), .Q ( signal_24066 ) ) ;
    buf_clk cell_9377 ( .C ( clk ), .D ( signal_24069 ), .Q ( signal_24070 ) ) ;
    buf_clk cell_9381 ( .C ( clk ), .D ( signal_24073 ), .Q ( signal_24074 ) ) ;
    buf_clk cell_9385 ( .C ( clk ), .D ( signal_24077 ), .Q ( signal_24078 ) ) ;
    buf_clk cell_9389 ( .C ( clk ), .D ( signal_24081 ), .Q ( signal_24082 ) ) ;
    buf_clk cell_9393 ( .C ( clk ), .D ( signal_24085 ), .Q ( signal_24086 ) ) ;
    buf_clk cell_9397 ( .C ( clk ), .D ( signal_24089 ), .Q ( signal_24090 ) ) ;
    buf_clk cell_9403 ( .C ( clk ), .D ( signal_24095 ), .Q ( signal_24096 ) ) ;
    buf_clk cell_9409 ( .C ( clk ), .D ( signal_24101 ), .Q ( signal_24102 ) ) ;
    buf_clk cell_9415 ( .C ( clk ), .D ( signal_24107 ), .Q ( signal_24108 ) ) ;
    buf_clk cell_9421 ( .C ( clk ), .D ( signal_24113 ), .Q ( signal_24114 ) ) ;
    buf_clk cell_9431 ( .C ( clk ), .D ( signal_24123 ), .Q ( signal_24124 ) ) ;
    buf_clk cell_9441 ( .C ( clk ), .D ( signal_24133 ), .Q ( signal_24134 ) ) ;
    buf_clk cell_9451 ( .C ( clk ), .D ( signal_24143 ), .Q ( signal_24144 ) ) ;
    buf_clk cell_9461 ( .C ( clk ), .D ( signal_24153 ), .Q ( signal_24154 ) ) ;
    buf_clk cell_9471 ( .C ( clk ), .D ( signal_24163 ), .Q ( signal_24164 ) ) ;
    buf_clk cell_9477 ( .C ( clk ), .D ( signal_24169 ), .Q ( signal_24170 ) ) ;
    buf_clk cell_9483 ( .C ( clk ), .D ( signal_24175 ), .Q ( signal_24176 ) ) ;
    buf_clk cell_9489 ( .C ( clk ), .D ( signal_24181 ), .Q ( signal_24182 ) ) ;
    buf_clk cell_9495 ( .C ( clk ), .D ( signal_24187 ), .Q ( signal_24188 ) ) ;
    buf_clk cell_9501 ( .C ( clk ), .D ( signal_24193 ), .Q ( signal_24194 ) ) ;
    buf_clk cell_9511 ( .C ( clk ), .D ( signal_24203 ), .Q ( signal_24204 ) ) ;
    buf_clk cell_9521 ( .C ( clk ), .D ( signal_24213 ), .Q ( signal_24214 ) ) ;
    buf_clk cell_9531 ( .C ( clk ), .D ( signal_24223 ), .Q ( signal_24224 ) ) ;
    buf_clk cell_9541 ( .C ( clk ), .D ( signal_24233 ), .Q ( signal_24234 ) ) ;
    buf_clk cell_9551 ( .C ( clk ), .D ( signal_24243 ), .Q ( signal_24244 ) ) ;
    buf_clk cell_9567 ( .C ( clk ), .D ( signal_24259 ), .Q ( signal_24260 ) ) ;
    buf_clk cell_9583 ( .C ( clk ), .D ( signal_24275 ), .Q ( signal_24276 ) ) ;
    buf_clk cell_9599 ( .C ( clk ), .D ( signal_24291 ), .Q ( signal_24292 ) ) ;
    buf_clk cell_9615 ( .C ( clk ), .D ( signal_24307 ), .Q ( signal_24308 ) ) ;
    buf_clk cell_9631 ( .C ( clk ), .D ( signal_24323 ), .Q ( signal_24324 ) ) ;
    buf_clk cell_9649 ( .C ( clk ), .D ( signal_24341 ), .Q ( signal_24342 ) ) ;
    buf_clk cell_9667 ( .C ( clk ), .D ( signal_24359 ), .Q ( signal_24360 ) ) ;
    buf_clk cell_9685 ( .C ( clk ), .D ( signal_24377 ), .Q ( signal_24378 ) ) ;
    buf_clk cell_9703 ( .C ( clk ), .D ( signal_24395 ), .Q ( signal_24396 ) ) ;
    buf_clk cell_9721 ( .C ( clk ), .D ( signal_24413 ), .Q ( signal_24414 ) ) ;
    buf_clk cell_9725 ( .C ( clk ), .D ( signal_2348 ), .Q ( signal_24418 ) ) ;
    buf_clk cell_9729 ( .C ( clk ), .D ( signal_8048 ), .Q ( signal_24422 ) ) ;
    buf_clk cell_9733 ( .C ( clk ), .D ( signal_8049 ), .Q ( signal_24426 ) ) ;
    buf_clk cell_9737 ( .C ( clk ), .D ( signal_8050 ), .Q ( signal_24430 ) ) ;
    buf_clk cell_9741 ( .C ( clk ), .D ( signal_8051 ), .Q ( signal_24434 ) ) ;
    buf_clk cell_9749 ( .C ( clk ), .D ( signal_24441 ), .Q ( signal_24442 ) ) ;
    buf_clk cell_9757 ( .C ( clk ), .D ( signal_24449 ), .Q ( signal_24450 ) ) ;
    buf_clk cell_9765 ( .C ( clk ), .D ( signal_24457 ), .Q ( signal_24458 ) ) ;
    buf_clk cell_9773 ( .C ( clk ), .D ( signal_24465 ), .Q ( signal_24466 ) ) ;
    buf_clk cell_9781 ( .C ( clk ), .D ( signal_24473 ), .Q ( signal_24474 ) ) ;
    buf_clk cell_9787 ( .C ( clk ), .D ( signal_24479 ), .Q ( signal_24480 ) ) ;
    buf_clk cell_9795 ( .C ( clk ), .D ( signal_24487 ), .Q ( signal_24488 ) ) ;
    buf_clk cell_9803 ( .C ( clk ), .D ( signal_24495 ), .Q ( signal_24496 ) ) ;
    buf_clk cell_9811 ( .C ( clk ), .D ( signal_24503 ), .Q ( signal_24504 ) ) ;
    buf_clk cell_9819 ( .C ( clk ), .D ( signal_24511 ), .Q ( signal_24512 ) ) ;
    buf_clk cell_9825 ( .C ( clk ), .D ( signal_2285 ), .Q ( signal_24518 ) ) ;
    buf_clk cell_9831 ( .C ( clk ), .D ( signal_7796 ), .Q ( signal_24524 ) ) ;
    buf_clk cell_9837 ( .C ( clk ), .D ( signal_7797 ), .Q ( signal_24530 ) ) ;
    buf_clk cell_9843 ( .C ( clk ), .D ( signal_7798 ), .Q ( signal_24536 ) ) ;
    buf_clk cell_9849 ( .C ( clk ), .D ( signal_7799 ), .Q ( signal_24542 ) ) ;
    buf_clk cell_9899 ( .C ( clk ), .D ( signal_24591 ), .Q ( signal_24592 ) ) ;
    buf_clk cell_9919 ( .C ( clk ), .D ( signal_24611 ), .Q ( signal_24612 ) ) ;
    buf_clk cell_9939 ( .C ( clk ), .D ( signal_24631 ), .Q ( signal_24632 ) ) ;
    buf_clk cell_9959 ( .C ( clk ), .D ( signal_24651 ), .Q ( signal_24652 ) ) ;
    buf_clk cell_9979 ( .C ( clk ), .D ( signal_24671 ), .Q ( signal_24672 ) ) ;
    buf_clk cell_9985 ( .C ( clk ), .D ( signal_2332 ), .Q ( signal_24678 ) ) ;
    buf_clk cell_9993 ( .C ( clk ), .D ( signal_7984 ), .Q ( signal_24686 ) ) ;
    buf_clk cell_10001 ( .C ( clk ), .D ( signal_7985 ), .Q ( signal_24694 ) ) ;
    buf_clk cell_10009 ( .C ( clk ), .D ( signal_7986 ), .Q ( signal_24702 ) ) ;
    buf_clk cell_10017 ( .C ( clk ), .D ( signal_7987 ), .Q ( signal_24710 ) ) ;
    buf_clk cell_10029 ( .C ( clk ), .D ( signal_24721 ), .Q ( signal_24722 ) ) ;
    buf_clk cell_10041 ( .C ( clk ), .D ( signal_24733 ), .Q ( signal_24734 ) ) ;
    buf_clk cell_10053 ( .C ( clk ), .D ( signal_24745 ), .Q ( signal_24746 ) ) ;
    buf_clk cell_10065 ( .C ( clk ), .D ( signal_24757 ), .Q ( signal_24758 ) ) ;
    buf_clk cell_10077 ( .C ( clk ), .D ( signal_24769 ), .Q ( signal_24770 ) ) ;
    buf_clk cell_10089 ( .C ( clk ), .D ( signal_24781 ), .Q ( signal_24782 ) ) ;
    buf_clk cell_10103 ( .C ( clk ), .D ( signal_24795 ), .Q ( signal_24796 ) ) ;
    buf_clk cell_10117 ( .C ( clk ), .D ( signal_24809 ), .Q ( signal_24810 ) ) ;
    buf_clk cell_10131 ( .C ( clk ), .D ( signal_24823 ), .Q ( signal_24824 ) ) ;
    buf_clk cell_10145 ( .C ( clk ), .D ( signal_24837 ), .Q ( signal_24838 ) ) ;
    buf_clk cell_10157 ( .C ( clk ), .D ( signal_24849 ), .Q ( signal_24850 ) ) ;
    buf_clk cell_10171 ( .C ( clk ), .D ( signal_24863 ), .Q ( signal_24864 ) ) ;
    buf_clk cell_10185 ( .C ( clk ), .D ( signal_24877 ), .Q ( signal_24878 ) ) ;
    buf_clk cell_10199 ( .C ( clk ), .D ( signal_24891 ), .Q ( signal_24892 ) ) ;
    buf_clk cell_10213 ( .C ( clk ), .D ( signal_24905 ), .Q ( signal_24906 ) ) ;

    /* cells in depth 22 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2319 ( .a ({signal_23407, signal_23399, signal_23391, signal_23383, signal_23375}), .b ({signal_7903, signal_7902, signal_7901, signal_7900, signal_2311}), .clk ( clk ), .r ({Fresh[8439], Fresh[8438], Fresh[8437], Fresh[8436], Fresh[8435], Fresh[8434], Fresh[8433], Fresh[8432], Fresh[8431], Fresh[8430]}), .c ({signal_7995, signal_7994, signal_7993, signal_7992, signal_2334}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2334 ( .a ({signal_23467, signal_23455, signal_23443, signal_23431, signal_23419}), .b ({signal_7983, signal_7982, signal_7981, signal_7980, signal_2331}), .clk ( clk ), .r ({Fresh[8449], Fresh[8448], Fresh[8447], Fresh[8446], Fresh[8445], Fresh[8444], Fresh[8443], Fresh[8442], Fresh[8441], Fresh[8440]}), .c ({signal_8055, signal_8054, signal_8053, signal_8052, signal_2349}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2338 ( .a ({signal_23497, signal_23491, signal_23485, signal_23479, signal_23473}), .b ({signal_8027, signal_8026, signal_8025, signal_8024, signal_2342}), .clk ( clk ), .r ({Fresh[8459], Fresh[8458], Fresh[8457], Fresh[8456], Fresh[8455], Fresh[8454], Fresh[8453], Fresh[8452], Fresh[8451], Fresh[8450]}), .c ({signal_8071, signal_8070, signal_8069, signal_8068, signal_2353}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2344 ( .a ({signal_8043, signal_8042, signal_8041, signal_8040, signal_2346}), .b ({signal_7795, signal_7794, signal_7793, signal_7792, signal_2284}), .clk ( clk ), .r ({Fresh[8469], Fresh[8468], Fresh[8467], Fresh[8466], Fresh[8465], Fresh[8464], Fresh[8463], Fresh[8462], Fresh[8461], Fresh[8460]}), .c ({signal_8095, signal_8094, signal_8093, signal_8092, signal_2359}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2346 ( .a ({signal_23527, signal_23521, signal_23515, signal_23509, signal_23503}), .b ({signal_8059, signal_8058, signal_8057, signal_8056, signal_2350}), .clk ( clk ), .r ({Fresh[8479], Fresh[8478], Fresh[8477], Fresh[8476], Fresh[8475], Fresh[8474], Fresh[8473], Fresh[8472], Fresh[8471], Fresh[8470]}), .c ({signal_8103, signal_8102, signal_8101, signal_8100, signal_2361}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2348 ( .a ({signal_23597, signal_23583, signal_23569, signal_23555, signal_23541}), .b ({signal_8079, signal_8078, signal_8077, signal_8076, signal_2355}), .clk ( clk ), .r ({Fresh[8489], Fresh[8488], Fresh[8487], Fresh[8486], Fresh[8485], Fresh[8484], Fresh[8483], Fresh[8482], Fresh[8481], Fresh[8480]}), .c ({signal_8111, signal_8110, signal_8109, signal_8108, signal_2363}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2349 ( .a ({signal_23637, signal_23629, signal_23621, signal_23613, signal_23605}), .b ({signal_8083, signal_8082, signal_8081, signal_8080, signal_2356}), .clk ( clk ), .r ({Fresh[8499], Fresh[8498], Fresh[8497], Fresh[8496], Fresh[8495], Fresh[8494], Fresh[8493], Fresh[8492], Fresh[8491], Fresh[8490]}), .c ({signal_8115, signal_8114, signal_8113, signal_8112, signal_2364}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2350 ( .a ({signal_23707, signal_23693, signal_23679, signal_23665, signal_23651}), .b ({signal_8063, signal_8062, signal_8061, signal_8060, signal_2351}), .clk ( clk ), .r ({Fresh[8509], Fresh[8508], Fresh[8507], Fresh[8506], Fresh[8505], Fresh[8504], Fresh[8503], Fresh[8502], Fresh[8501], Fresh[8500]}), .c ({signal_8119, signal_8118, signal_8117, signal_8116, signal_2365}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2351 ( .a ({signal_23747, signal_23739, signal_23731, signal_23723, signal_23715}), .b ({signal_8091, signal_8090, signal_8089, signal_8088, signal_2358}), .clk ( clk ), .r ({Fresh[8519], Fresh[8518], Fresh[8517], Fresh[8516], Fresh[8515], Fresh[8514], Fresh[8513], Fresh[8512], Fresh[8511], Fresh[8510]}), .c ({signal_8123, signal_8122, signal_8121, signal_8120, signal_2366}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2352 ( .a ({signal_8067, signal_8066, signal_8065, signal_8064, signal_2352}), .b ({signal_7991, signal_7990, signal_7989, signal_7988, signal_2333}), .clk ( clk ), .r ({Fresh[8529], Fresh[8528], Fresh[8527], Fresh[8526], Fresh[8525], Fresh[8524], Fresh[8523], Fresh[8522], Fresh[8521], Fresh[8520]}), .c ({signal_8127, signal_8126, signal_8125, signal_8124, signal_2367}) ) ;
    buf_clk cell_9058 ( .C ( clk ), .D ( signal_23750 ), .Q ( signal_23751 ) ) ;
    buf_clk cell_9062 ( .C ( clk ), .D ( signal_23754 ), .Q ( signal_23755 ) ) ;
    buf_clk cell_9066 ( .C ( clk ), .D ( signal_23758 ), .Q ( signal_23759 ) ) ;
    buf_clk cell_9070 ( .C ( clk ), .D ( signal_23762 ), .Q ( signal_23763 ) ) ;
    buf_clk cell_9074 ( .C ( clk ), .D ( signal_23766 ), .Q ( signal_23767 ) ) ;
    buf_clk cell_9084 ( .C ( clk ), .D ( signal_23776 ), .Q ( signal_23777 ) ) ;
    buf_clk cell_9094 ( .C ( clk ), .D ( signal_23786 ), .Q ( signal_23787 ) ) ;
    buf_clk cell_9104 ( .C ( clk ), .D ( signal_23796 ), .Q ( signal_23797 ) ) ;
    buf_clk cell_9114 ( .C ( clk ), .D ( signal_23806 ), .Q ( signal_23807 ) ) ;
    buf_clk cell_9124 ( .C ( clk ), .D ( signal_23816 ), .Q ( signal_23817 ) ) ;
    buf_clk cell_9126 ( .C ( clk ), .D ( signal_23818 ), .Q ( signal_23819 ) ) ;
    buf_clk cell_9128 ( .C ( clk ), .D ( signal_23820 ), .Q ( signal_23821 ) ) ;
    buf_clk cell_9130 ( .C ( clk ), .D ( signal_23822 ), .Q ( signal_23823 ) ) ;
    buf_clk cell_9132 ( .C ( clk ), .D ( signal_23824 ), .Q ( signal_23825 ) ) ;
    buf_clk cell_9134 ( .C ( clk ), .D ( signal_23826 ), .Q ( signal_23827 ) ) ;
    buf_clk cell_9136 ( .C ( clk ), .D ( signal_23828 ), .Q ( signal_23829 ) ) ;
    buf_clk cell_9138 ( .C ( clk ), .D ( signal_23830 ), .Q ( signal_23831 ) ) ;
    buf_clk cell_9140 ( .C ( clk ), .D ( signal_23832 ), .Q ( signal_23833 ) ) ;
    buf_clk cell_9142 ( .C ( clk ), .D ( signal_23834 ), .Q ( signal_23835 ) ) ;
    buf_clk cell_9144 ( .C ( clk ), .D ( signal_23836 ), .Q ( signal_23837 ) ) ;
    buf_clk cell_9160 ( .C ( clk ), .D ( signal_23852 ), .Q ( signal_23853 ) ) ;
    buf_clk cell_9176 ( .C ( clk ), .D ( signal_23868 ), .Q ( signal_23869 ) ) ;
    buf_clk cell_9192 ( .C ( clk ), .D ( signal_23884 ), .Q ( signal_23885 ) ) ;
    buf_clk cell_9208 ( .C ( clk ), .D ( signal_23900 ), .Q ( signal_23901 ) ) ;
    buf_clk cell_9224 ( .C ( clk ), .D ( signal_23916 ), .Q ( signal_23917 ) ) ;
    buf_clk cell_9228 ( .C ( clk ), .D ( signal_23920 ), .Q ( signal_23921 ) ) ;
    buf_clk cell_9232 ( .C ( clk ), .D ( signal_23924 ), .Q ( signal_23925 ) ) ;
    buf_clk cell_9236 ( .C ( clk ), .D ( signal_23928 ), .Q ( signal_23929 ) ) ;
    buf_clk cell_9240 ( .C ( clk ), .D ( signal_23932 ), .Q ( signal_23933 ) ) ;
    buf_clk cell_9244 ( .C ( clk ), .D ( signal_23936 ), .Q ( signal_23937 ) ) ;
    buf_clk cell_9260 ( .C ( clk ), .D ( signal_23952 ), .Q ( signal_23953 ) ) ;
    buf_clk cell_9276 ( .C ( clk ), .D ( signal_23968 ), .Q ( signal_23969 ) ) ;
    buf_clk cell_9292 ( .C ( clk ), .D ( signal_23984 ), .Q ( signal_23985 ) ) ;
    buf_clk cell_9308 ( .C ( clk ), .D ( signal_24000 ), .Q ( signal_24001 ) ) ;
    buf_clk cell_9324 ( .C ( clk ), .D ( signal_24016 ), .Q ( signal_24017 ) ) ;
    buf_clk cell_9334 ( .C ( clk ), .D ( signal_24026 ), .Q ( signal_24027 ) ) ;
    buf_clk cell_9344 ( .C ( clk ), .D ( signal_24036 ), .Q ( signal_24037 ) ) ;
    buf_clk cell_9354 ( .C ( clk ), .D ( signal_24046 ), .Q ( signal_24047 ) ) ;
    buf_clk cell_9364 ( .C ( clk ), .D ( signal_24056 ), .Q ( signal_24057 ) ) ;
    buf_clk cell_9374 ( .C ( clk ), .D ( signal_24066 ), .Q ( signal_24067 ) ) ;
    buf_clk cell_9378 ( .C ( clk ), .D ( signal_24070 ), .Q ( signal_24071 ) ) ;
    buf_clk cell_9382 ( .C ( clk ), .D ( signal_24074 ), .Q ( signal_24075 ) ) ;
    buf_clk cell_9386 ( .C ( clk ), .D ( signal_24078 ), .Q ( signal_24079 ) ) ;
    buf_clk cell_9390 ( .C ( clk ), .D ( signal_24082 ), .Q ( signal_24083 ) ) ;
    buf_clk cell_9394 ( .C ( clk ), .D ( signal_24086 ), .Q ( signal_24087 ) ) ;
    buf_clk cell_9398 ( .C ( clk ), .D ( signal_24090 ), .Q ( signal_24091 ) ) ;
    buf_clk cell_9404 ( .C ( clk ), .D ( signal_24096 ), .Q ( signal_24097 ) ) ;
    buf_clk cell_9410 ( .C ( clk ), .D ( signal_24102 ), .Q ( signal_24103 ) ) ;
    buf_clk cell_9416 ( .C ( clk ), .D ( signal_24108 ), .Q ( signal_24109 ) ) ;
    buf_clk cell_9422 ( .C ( clk ), .D ( signal_24114 ), .Q ( signal_24115 ) ) ;
    buf_clk cell_9432 ( .C ( clk ), .D ( signal_24124 ), .Q ( signal_24125 ) ) ;
    buf_clk cell_9442 ( .C ( clk ), .D ( signal_24134 ), .Q ( signal_24135 ) ) ;
    buf_clk cell_9452 ( .C ( clk ), .D ( signal_24144 ), .Q ( signal_24145 ) ) ;
    buf_clk cell_9462 ( .C ( clk ), .D ( signal_24154 ), .Q ( signal_24155 ) ) ;
    buf_clk cell_9472 ( .C ( clk ), .D ( signal_24164 ), .Q ( signal_24165 ) ) ;
    buf_clk cell_9478 ( .C ( clk ), .D ( signal_24170 ), .Q ( signal_24171 ) ) ;
    buf_clk cell_9484 ( .C ( clk ), .D ( signal_24176 ), .Q ( signal_24177 ) ) ;
    buf_clk cell_9490 ( .C ( clk ), .D ( signal_24182 ), .Q ( signal_24183 ) ) ;
    buf_clk cell_9496 ( .C ( clk ), .D ( signal_24188 ), .Q ( signal_24189 ) ) ;
    buf_clk cell_9502 ( .C ( clk ), .D ( signal_24194 ), .Q ( signal_24195 ) ) ;
    buf_clk cell_9512 ( .C ( clk ), .D ( signal_24204 ), .Q ( signal_24205 ) ) ;
    buf_clk cell_9522 ( .C ( clk ), .D ( signal_24214 ), .Q ( signal_24215 ) ) ;
    buf_clk cell_9532 ( .C ( clk ), .D ( signal_24224 ), .Q ( signal_24225 ) ) ;
    buf_clk cell_9542 ( .C ( clk ), .D ( signal_24234 ), .Q ( signal_24235 ) ) ;
    buf_clk cell_9552 ( .C ( clk ), .D ( signal_24244 ), .Q ( signal_24245 ) ) ;
    buf_clk cell_9568 ( .C ( clk ), .D ( signal_24260 ), .Q ( signal_24261 ) ) ;
    buf_clk cell_9584 ( .C ( clk ), .D ( signal_24276 ), .Q ( signal_24277 ) ) ;
    buf_clk cell_9600 ( .C ( clk ), .D ( signal_24292 ), .Q ( signal_24293 ) ) ;
    buf_clk cell_9616 ( .C ( clk ), .D ( signal_24308 ), .Q ( signal_24309 ) ) ;
    buf_clk cell_9632 ( .C ( clk ), .D ( signal_24324 ), .Q ( signal_24325 ) ) ;
    buf_clk cell_9650 ( .C ( clk ), .D ( signal_24342 ), .Q ( signal_24343 ) ) ;
    buf_clk cell_9668 ( .C ( clk ), .D ( signal_24360 ), .Q ( signal_24361 ) ) ;
    buf_clk cell_9686 ( .C ( clk ), .D ( signal_24378 ), .Q ( signal_24379 ) ) ;
    buf_clk cell_9704 ( .C ( clk ), .D ( signal_24396 ), .Q ( signal_24397 ) ) ;
    buf_clk cell_9722 ( .C ( clk ), .D ( signal_24414 ), .Q ( signal_24415 ) ) ;
    buf_clk cell_9726 ( .C ( clk ), .D ( signal_24418 ), .Q ( signal_24419 ) ) ;
    buf_clk cell_9730 ( .C ( clk ), .D ( signal_24422 ), .Q ( signal_24423 ) ) ;
    buf_clk cell_9734 ( .C ( clk ), .D ( signal_24426 ), .Q ( signal_24427 ) ) ;
    buf_clk cell_9738 ( .C ( clk ), .D ( signal_24430 ), .Q ( signal_24431 ) ) ;
    buf_clk cell_9742 ( .C ( clk ), .D ( signal_24434 ), .Q ( signal_24435 ) ) ;
    buf_clk cell_9750 ( .C ( clk ), .D ( signal_24442 ), .Q ( signal_24443 ) ) ;
    buf_clk cell_9758 ( .C ( clk ), .D ( signal_24450 ), .Q ( signal_24451 ) ) ;
    buf_clk cell_9766 ( .C ( clk ), .D ( signal_24458 ), .Q ( signal_24459 ) ) ;
    buf_clk cell_9774 ( .C ( clk ), .D ( signal_24466 ), .Q ( signal_24467 ) ) ;
    buf_clk cell_9782 ( .C ( clk ), .D ( signal_24474 ), .Q ( signal_24475 ) ) ;
    buf_clk cell_9788 ( .C ( clk ), .D ( signal_24480 ), .Q ( signal_24481 ) ) ;
    buf_clk cell_9796 ( .C ( clk ), .D ( signal_24488 ), .Q ( signal_24489 ) ) ;
    buf_clk cell_9804 ( .C ( clk ), .D ( signal_24496 ), .Q ( signal_24497 ) ) ;
    buf_clk cell_9812 ( .C ( clk ), .D ( signal_24504 ), .Q ( signal_24505 ) ) ;
    buf_clk cell_9820 ( .C ( clk ), .D ( signal_24512 ), .Q ( signal_24513 ) ) ;
    buf_clk cell_9826 ( .C ( clk ), .D ( signal_24518 ), .Q ( signal_24519 ) ) ;
    buf_clk cell_9832 ( .C ( clk ), .D ( signal_24524 ), .Q ( signal_24525 ) ) ;
    buf_clk cell_9838 ( .C ( clk ), .D ( signal_24530 ), .Q ( signal_24531 ) ) ;
    buf_clk cell_9844 ( .C ( clk ), .D ( signal_24536 ), .Q ( signal_24537 ) ) ;
    buf_clk cell_9850 ( .C ( clk ), .D ( signal_24542 ), .Q ( signal_24543 ) ) ;
    buf_clk cell_9900 ( .C ( clk ), .D ( signal_24592 ), .Q ( signal_24593 ) ) ;
    buf_clk cell_9920 ( .C ( clk ), .D ( signal_24612 ), .Q ( signal_24613 ) ) ;
    buf_clk cell_9940 ( .C ( clk ), .D ( signal_24632 ), .Q ( signal_24633 ) ) ;
    buf_clk cell_9960 ( .C ( clk ), .D ( signal_24652 ), .Q ( signal_24653 ) ) ;
    buf_clk cell_9980 ( .C ( clk ), .D ( signal_24672 ), .Q ( signal_24673 ) ) ;
    buf_clk cell_9986 ( .C ( clk ), .D ( signal_24678 ), .Q ( signal_24679 ) ) ;
    buf_clk cell_9994 ( .C ( clk ), .D ( signal_24686 ), .Q ( signal_24687 ) ) ;
    buf_clk cell_10002 ( .C ( clk ), .D ( signal_24694 ), .Q ( signal_24695 ) ) ;
    buf_clk cell_10010 ( .C ( clk ), .D ( signal_24702 ), .Q ( signal_24703 ) ) ;
    buf_clk cell_10018 ( .C ( clk ), .D ( signal_24710 ), .Q ( signal_24711 ) ) ;
    buf_clk cell_10030 ( .C ( clk ), .D ( signal_24722 ), .Q ( signal_24723 ) ) ;
    buf_clk cell_10042 ( .C ( clk ), .D ( signal_24734 ), .Q ( signal_24735 ) ) ;
    buf_clk cell_10054 ( .C ( clk ), .D ( signal_24746 ), .Q ( signal_24747 ) ) ;
    buf_clk cell_10066 ( .C ( clk ), .D ( signal_24758 ), .Q ( signal_24759 ) ) ;
    buf_clk cell_10078 ( .C ( clk ), .D ( signal_24770 ), .Q ( signal_24771 ) ) ;
    buf_clk cell_10090 ( .C ( clk ), .D ( signal_24782 ), .Q ( signal_24783 ) ) ;
    buf_clk cell_10104 ( .C ( clk ), .D ( signal_24796 ), .Q ( signal_24797 ) ) ;
    buf_clk cell_10118 ( .C ( clk ), .D ( signal_24810 ), .Q ( signal_24811 ) ) ;
    buf_clk cell_10132 ( .C ( clk ), .D ( signal_24824 ), .Q ( signal_24825 ) ) ;
    buf_clk cell_10146 ( .C ( clk ), .D ( signal_24838 ), .Q ( signal_24839 ) ) ;
    buf_clk cell_10158 ( .C ( clk ), .D ( signal_24850 ), .Q ( signal_24851 ) ) ;
    buf_clk cell_10172 ( .C ( clk ), .D ( signal_24864 ), .Q ( signal_24865 ) ) ;
    buf_clk cell_10186 ( .C ( clk ), .D ( signal_24878 ), .Q ( signal_24879 ) ) ;
    buf_clk cell_10200 ( .C ( clk ), .D ( signal_24892 ), .Q ( signal_24893 ) ) ;
    buf_clk cell_10214 ( .C ( clk ), .D ( signal_24906 ), .Q ( signal_24907 ) ) ;

    /* cells in depth 23 */
    buf_clk cell_9399 ( .C ( clk ), .D ( signal_24091 ), .Q ( signal_24092 ) ) ;
    buf_clk cell_9405 ( .C ( clk ), .D ( signal_24097 ), .Q ( signal_24098 ) ) ;
    buf_clk cell_9411 ( .C ( clk ), .D ( signal_24103 ), .Q ( signal_24104 ) ) ;
    buf_clk cell_9417 ( .C ( clk ), .D ( signal_24109 ), .Q ( signal_24110 ) ) ;
    buf_clk cell_9423 ( .C ( clk ), .D ( signal_24115 ), .Q ( signal_24116 ) ) ;
    buf_clk cell_9433 ( .C ( clk ), .D ( signal_24125 ), .Q ( signal_24126 ) ) ;
    buf_clk cell_9443 ( .C ( clk ), .D ( signal_24135 ), .Q ( signal_24136 ) ) ;
    buf_clk cell_9453 ( .C ( clk ), .D ( signal_24145 ), .Q ( signal_24146 ) ) ;
    buf_clk cell_9463 ( .C ( clk ), .D ( signal_24155 ), .Q ( signal_24156 ) ) ;
    buf_clk cell_9473 ( .C ( clk ), .D ( signal_24165 ), .Q ( signal_24166 ) ) ;
    buf_clk cell_9479 ( .C ( clk ), .D ( signal_24171 ), .Q ( signal_24172 ) ) ;
    buf_clk cell_9485 ( .C ( clk ), .D ( signal_24177 ), .Q ( signal_24178 ) ) ;
    buf_clk cell_9491 ( .C ( clk ), .D ( signal_24183 ), .Q ( signal_24184 ) ) ;
    buf_clk cell_9497 ( .C ( clk ), .D ( signal_24189 ), .Q ( signal_24190 ) ) ;
    buf_clk cell_9503 ( .C ( clk ), .D ( signal_24195 ), .Q ( signal_24196 ) ) ;
    buf_clk cell_9513 ( .C ( clk ), .D ( signal_24205 ), .Q ( signal_24206 ) ) ;
    buf_clk cell_9523 ( .C ( clk ), .D ( signal_24215 ), .Q ( signal_24216 ) ) ;
    buf_clk cell_9533 ( .C ( clk ), .D ( signal_24225 ), .Q ( signal_24226 ) ) ;
    buf_clk cell_9543 ( .C ( clk ), .D ( signal_24235 ), .Q ( signal_24236 ) ) ;
    buf_clk cell_9553 ( .C ( clk ), .D ( signal_24245 ), .Q ( signal_24246 ) ) ;
    buf_clk cell_9569 ( .C ( clk ), .D ( signal_24261 ), .Q ( signal_24262 ) ) ;
    buf_clk cell_9585 ( .C ( clk ), .D ( signal_24277 ), .Q ( signal_24278 ) ) ;
    buf_clk cell_9601 ( .C ( clk ), .D ( signal_24293 ), .Q ( signal_24294 ) ) ;
    buf_clk cell_9617 ( .C ( clk ), .D ( signal_24309 ), .Q ( signal_24310 ) ) ;
    buf_clk cell_9633 ( .C ( clk ), .D ( signal_24325 ), .Q ( signal_24326 ) ) ;
    buf_clk cell_9651 ( .C ( clk ), .D ( signal_24343 ), .Q ( signal_24344 ) ) ;
    buf_clk cell_9669 ( .C ( clk ), .D ( signal_24361 ), .Q ( signal_24362 ) ) ;
    buf_clk cell_9687 ( .C ( clk ), .D ( signal_24379 ), .Q ( signal_24380 ) ) ;
    buf_clk cell_9705 ( .C ( clk ), .D ( signal_24397 ), .Q ( signal_24398 ) ) ;
    buf_clk cell_9723 ( .C ( clk ), .D ( signal_24415 ), .Q ( signal_24416 ) ) ;
    buf_clk cell_9727 ( .C ( clk ), .D ( signal_24419 ), .Q ( signal_24420 ) ) ;
    buf_clk cell_9731 ( .C ( clk ), .D ( signal_24423 ), .Q ( signal_24424 ) ) ;
    buf_clk cell_9735 ( .C ( clk ), .D ( signal_24427 ), .Q ( signal_24428 ) ) ;
    buf_clk cell_9739 ( .C ( clk ), .D ( signal_24431 ), .Q ( signal_24432 ) ) ;
    buf_clk cell_9743 ( .C ( clk ), .D ( signal_24435 ), .Q ( signal_24436 ) ) ;
    buf_clk cell_9751 ( .C ( clk ), .D ( signal_24443 ), .Q ( signal_24444 ) ) ;
    buf_clk cell_9759 ( .C ( clk ), .D ( signal_24451 ), .Q ( signal_24452 ) ) ;
    buf_clk cell_9767 ( .C ( clk ), .D ( signal_24459 ), .Q ( signal_24460 ) ) ;
    buf_clk cell_9775 ( .C ( clk ), .D ( signal_24467 ), .Q ( signal_24468 ) ) ;
    buf_clk cell_9783 ( .C ( clk ), .D ( signal_24475 ), .Q ( signal_24476 ) ) ;
    buf_clk cell_9789 ( .C ( clk ), .D ( signal_24481 ), .Q ( signal_24482 ) ) ;
    buf_clk cell_9797 ( .C ( clk ), .D ( signal_24489 ), .Q ( signal_24490 ) ) ;
    buf_clk cell_9805 ( .C ( clk ), .D ( signal_24497 ), .Q ( signal_24498 ) ) ;
    buf_clk cell_9813 ( .C ( clk ), .D ( signal_24505 ), .Q ( signal_24506 ) ) ;
    buf_clk cell_9821 ( .C ( clk ), .D ( signal_24513 ), .Q ( signal_24514 ) ) ;
    buf_clk cell_9827 ( .C ( clk ), .D ( signal_24519 ), .Q ( signal_24520 ) ) ;
    buf_clk cell_9833 ( .C ( clk ), .D ( signal_24525 ), .Q ( signal_24526 ) ) ;
    buf_clk cell_9839 ( .C ( clk ), .D ( signal_24531 ), .Q ( signal_24532 ) ) ;
    buf_clk cell_9845 ( .C ( clk ), .D ( signal_24537 ), .Q ( signal_24538 ) ) ;
    buf_clk cell_9851 ( .C ( clk ), .D ( signal_24543 ), .Q ( signal_24544 ) ) ;
    buf_clk cell_9855 ( .C ( clk ), .D ( signal_2361 ), .Q ( signal_24548 ) ) ;
    buf_clk cell_9859 ( .C ( clk ), .D ( signal_8100 ), .Q ( signal_24552 ) ) ;
    buf_clk cell_9863 ( .C ( clk ), .D ( signal_8101 ), .Q ( signal_24556 ) ) ;
    buf_clk cell_9867 ( .C ( clk ), .D ( signal_8102 ), .Q ( signal_24560 ) ) ;
    buf_clk cell_9871 ( .C ( clk ), .D ( signal_8103 ), .Q ( signal_24564 ) ) ;
    buf_clk cell_9901 ( .C ( clk ), .D ( signal_24593 ), .Q ( signal_24594 ) ) ;
    buf_clk cell_9921 ( .C ( clk ), .D ( signal_24613 ), .Q ( signal_24614 ) ) ;
    buf_clk cell_9941 ( .C ( clk ), .D ( signal_24633 ), .Q ( signal_24634 ) ) ;
    buf_clk cell_9961 ( .C ( clk ), .D ( signal_24653 ), .Q ( signal_24654 ) ) ;
    buf_clk cell_9981 ( .C ( clk ), .D ( signal_24673 ), .Q ( signal_24674 ) ) ;
    buf_clk cell_9987 ( .C ( clk ), .D ( signal_24679 ), .Q ( signal_24680 ) ) ;
    buf_clk cell_9995 ( .C ( clk ), .D ( signal_24687 ), .Q ( signal_24688 ) ) ;
    buf_clk cell_10003 ( .C ( clk ), .D ( signal_24695 ), .Q ( signal_24696 ) ) ;
    buf_clk cell_10011 ( .C ( clk ), .D ( signal_24703 ), .Q ( signal_24704 ) ) ;
    buf_clk cell_10019 ( .C ( clk ), .D ( signal_24711 ), .Q ( signal_24712 ) ) ;
    buf_clk cell_10031 ( .C ( clk ), .D ( signal_24723 ), .Q ( signal_24724 ) ) ;
    buf_clk cell_10043 ( .C ( clk ), .D ( signal_24735 ), .Q ( signal_24736 ) ) ;
    buf_clk cell_10055 ( .C ( clk ), .D ( signal_24747 ), .Q ( signal_24748 ) ) ;
    buf_clk cell_10067 ( .C ( clk ), .D ( signal_24759 ), .Q ( signal_24760 ) ) ;
    buf_clk cell_10079 ( .C ( clk ), .D ( signal_24771 ), .Q ( signal_24772 ) ) ;
    buf_clk cell_10091 ( .C ( clk ), .D ( signal_24783 ), .Q ( signal_24784 ) ) ;
    buf_clk cell_10105 ( .C ( clk ), .D ( signal_24797 ), .Q ( signal_24798 ) ) ;
    buf_clk cell_10119 ( .C ( clk ), .D ( signal_24811 ), .Q ( signal_24812 ) ) ;
    buf_clk cell_10133 ( .C ( clk ), .D ( signal_24825 ), .Q ( signal_24826 ) ) ;
    buf_clk cell_10147 ( .C ( clk ), .D ( signal_24839 ), .Q ( signal_24840 ) ) ;
    buf_clk cell_10159 ( .C ( clk ), .D ( signal_24851 ), .Q ( signal_24852 ) ) ;
    buf_clk cell_10173 ( .C ( clk ), .D ( signal_24865 ), .Q ( signal_24866 ) ) ;
    buf_clk cell_10187 ( .C ( clk ), .D ( signal_24879 ), .Q ( signal_24880 ) ) ;
    buf_clk cell_10201 ( .C ( clk ), .D ( signal_24893 ), .Q ( signal_24894 ) ) ;
    buf_clk cell_10215 ( .C ( clk ), .D ( signal_24907 ), .Q ( signal_24908 ) ) ;

    /* cells in depth 24 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2345 ( .a ({signal_23767, signal_23763, signal_23759, signal_23755, signal_23751}), .b ({signal_7995, signal_7994, signal_7993, signal_7992, signal_2334}), .clk ( clk ), .r ({Fresh[8539], Fresh[8538], Fresh[8537], Fresh[8536], Fresh[8535], Fresh[8534], Fresh[8533], Fresh[8532], Fresh[8531], Fresh[8530]}), .c ({signal_8099, signal_8098, signal_8097, signal_8096, signal_2360}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2347 ( .a ({signal_23817, signal_23807, signal_23797, signal_23787, signal_23777}), .b ({signal_8071, signal_8070, signal_8069, signal_8068, signal_2353}), .clk ( clk ), .r ({Fresh[8549], Fresh[8548], Fresh[8547], Fresh[8546], Fresh[8545], Fresh[8544], Fresh[8543], Fresh[8542], Fresh[8541], Fresh[8540]}), .c ({signal_8107, signal_8106, signal_8105, signal_8104, signal_2362}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2353 ( .a ({signal_23827, signal_23825, signal_23823, signal_23821, signal_23819}), .b ({signal_8055, signal_8054, signal_8053, signal_8052, signal_2349}), .clk ( clk ), .r ({Fresh[8559], Fresh[8558], Fresh[8557], Fresh[8556], Fresh[8555], Fresh[8554], Fresh[8553], Fresh[8552], Fresh[8551], Fresh[8550]}), .c ({signal_8131, signal_8130, signal_8129, signal_8128, signal_2368}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2354 ( .a ({signal_23837, signal_23835, signal_23833, signal_23831, signal_23829}), .b ({signal_8095, signal_8094, signal_8093, signal_8092, signal_2359}), .clk ( clk ), .r ({Fresh[8569], Fresh[8568], Fresh[8567], Fresh[8566], Fresh[8565], Fresh[8564], Fresh[8563], Fresh[8562], Fresh[8561], Fresh[8560]}), .c ({signal_8135, signal_8134, signal_8133, signal_8132, signal_2369}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2357 ( .a ({signal_23917, signal_23901, signal_23885, signal_23869, signal_23853}), .b ({signal_8111, signal_8110, signal_8109, signal_8108, signal_2363}), .clk ( clk ), .r ({Fresh[8579], Fresh[8578], Fresh[8577], Fresh[8576], Fresh[8575], Fresh[8574], Fresh[8573], Fresh[8572], Fresh[8571], Fresh[8570]}), .c ({signal_8147, signal_8146, signal_8145, signal_8144, signal_2372}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2358 ( .a ({signal_23937, signal_23933, signal_23929, signal_23925, signal_23921}), .b ({signal_8115, signal_8114, signal_8113, signal_8112, signal_2364}), .clk ( clk ), .r ({Fresh[8589], Fresh[8588], Fresh[8587], Fresh[8586], Fresh[8585], Fresh[8584], Fresh[8583], Fresh[8582], Fresh[8581], Fresh[8580]}), .c ({signal_8151, signal_8150, signal_8149, signal_8148, signal_2373}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2359 ( .a ({signal_24017, signal_24001, signal_23985, signal_23969, signal_23953}), .b ({signal_8119, signal_8118, signal_8117, signal_8116, signal_2365}), .clk ( clk ), .r ({Fresh[8599], Fresh[8598], Fresh[8597], Fresh[8596], Fresh[8595], Fresh[8594], Fresh[8593], Fresh[8592], Fresh[8591], Fresh[8590]}), .c ({signal_8155, signal_8154, signal_8153, signal_8152, signal_2374}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2360 ( .a ({signal_24067, signal_24057, signal_24047, signal_24037, signal_24027}), .b ({signal_8123, signal_8122, signal_8121, signal_8120, signal_2366}), .clk ( clk ), .r ({Fresh[8609], Fresh[8608], Fresh[8607], Fresh[8606], Fresh[8605], Fresh[8604], Fresh[8603], Fresh[8602], Fresh[8601], Fresh[8600]}), .c ({signal_8159, signal_8158, signal_8157, signal_8156, signal_2375}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2361 ( .a ({signal_24087, signal_24083, signal_24079, signal_24075, signal_24071}), .b ({signal_8127, signal_8126, signal_8125, signal_8124, signal_2367}), .clk ( clk ), .r ({Fresh[8619], Fresh[8618], Fresh[8617], Fresh[8616], Fresh[8615], Fresh[8614], Fresh[8613], Fresh[8612], Fresh[8611], Fresh[8610]}), .c ({signal_8163, signal_8162, signal_8161, signal_8160, signal_2376}) ) ;
    buf_clk cell_9400 ( .C ( clk ), .D ( signal_24092 ), .Q ( signal_24093 ) ) ;
    buf_clk cell_9406 ( .C ( clk ), .D ( signal_24098 ), .Q ( signal_24099 ) ) ;
    buf_clk cell_9412 ( .C ( clk ), .D ( signal_24104 ), .Q ( signal_24105 ) ) ;
    buf_clk cell_9418 ( .C ( clk ), .D ( signal_24110 ), .Q ( signal_24111 ) ) ;
    buf_clk cell_9424 ( .C ( clk ), .D ( signal_24116 ), .Q ( signal_24117 ) ) ;
    buf_clk cell_9434 ( .C ( clk ), .D ( signal_24126 ), .Q ( signal_24127 ) ) ;
    buf_clk cell_9444 ( .C ( clk ), .D ( signal_24136 ), .Q ( signal_24137 ) ) ;
    buf_clk cell_9454 ( .C ( clk ), .D ( signal_24146 ), .Q ( signal_24147 ) ) ;
    buf_clk cell_9464 ( .C ( clk ), .D ( signal_24156 ), .Q ( signal_24157 ) ) ;
    buf_clk cell_9474 ( .C ( clk ), .D ( signal_24166 ), .Q ( signal_24167 ) ) ;
    buf_clk cell_9480 ( .C ( clk ), .D ( signal_24172 ), .Q ( signal_24173 ) ) ;
    buf_clk cell_9486 ( .C ( clk ), .D ( signal_24178 ), .Q ( signal_24179 ) ) ;
    buf_clk cell_9492 ( .C ( clk ), .D ( signal_24184 ), .Q ( signal_24185 ) ) ;
    buf_clk cell_9498 ( .C ( clk ), .D ( signal_24190 ), .Q ( signal_24191 ) ) ;
    buf_clk cell_9504 ( .C ( clk ), .D ( signal_24196 ), .Q ( signal_24197 ) ) ;
    buf_clk cell_9514 ( .C ( clk ), .D ( signal_24206 ), .Q ( signal_24207 ) ) ;
    buf_clk cell_9524 ( .C ( clk ), .D ( signal_24216 ), .Q ( signal_24217 ) ) ;
    buf_clk cell_9534 ( .C ( clk ), .D ( signal_24226 ), .Q ( signal_24227 ) ) ;
    buf_clk cell_9544 ( .C ( clk ), .D ( signal_24236 ), .Q ( signal_24237 ) ) ;
    buf_clk cell_9554 ( .C ( clk ), .D ( signal_24246 ), .Q ( signal_24247 ) ) ;
    buf_clk cell_9570 ( .C ( clk ), .D ( signal_24262 ), .Q ( signal_24263 ) ) ;
    buf_clk cell_9586 ( .C ( clk ), .D ( signal_24278 ), .Q ( signal_24279 ) ) ;
    buf_clk cell_9602 ( .C ( clk ), .D ( signal_24294 ), .Q ( signal_24295 ) ) ;
    buf_clk cell_9618 ( .C ( clk ), .D ( signal_24310 ), .Q ( signal_24311 ) ) ;
    buf_clk cell_9634 ( .C ( clk ), .D ( signal_24326 ), .Q ( signal_24327 ) ) ;
    buf_clk cell_9652 ( .C ( clk ), .D ( signal_24344 ), .Q ( signal_24345 ) ) ;
    buf_clk cell_9670 ( .C ( clk ), .D ( signal_24362 ), .Q ( signal_24363 ) ) ;
    buf_clk cell_9688 ( .C ( clk ), .D ( signal_24380 ), .Q ( signal_24381 ) ) ;
    buf_clk cell_9706 ( .C ( clk ), .D ( signal_24398 ), .Q ( signal_24399 ) ) ;
    buf_clk cell_9724 ( .C ( clk ), .D ( signal_24416 ), .Q ( signal_24417 ) ) ;
    buf_clk cell_9728 ( .C ( clk ), .D ( signal_24420 ), .Q ( signal_24421 ) ) ;
    buf_clk cell_9732 ( .C ( clk ), .D ( signal_24424 ), .Q ( signal_24425 ) ) ;
    buf_clk cell_9736 ( .C ( clk ), .D ( signal_24428 ), .Q ( signal_24429 ) ) ;
    buf_clk cell_9740 ( .C ( clk ), .D ( signal_24432 ), .Q ( signal_24433 ) ) ;
    buf_clk cell_9744 ( .C ( clk ), .D ( signal_24436 ), .Q ( signal_24437 ) ) ;
    buf_clk cell_9752 ( .C ( clk ), .D ( signal_24444 ), .Q ( signal_24445 ) ) ;
    buf_clk cell_9760 ( .C ( clk ), .D ( signal_24452 ), .Q ( signal_24453 ) ) ;
    buf_clk cell_9768 ( .C ( clk ), .D ( signal_24460 ), .Q ( signal_24461 ) ) ;
    buf_clk cell_9776 ( .C ( clk ), .D ( signal_24468 ), .Q ( signal_24469 ) ) ;
    buf_clk cell_9784 ( .C ( clk ), .D ( signal_24476 ), .Q ( signal_24477 ) ) ;
    buf_clk cell_9790 ( .C ( clk ), .D ( signal_24482 ), .Q ( signal_24483 ) ) ;
    buf_clk cell_9798 ( .C ( clk ), .D ( signal_24490 ), .Q ( signal_24491 ) ) ;
    buf_clk cell_9806 ( .C ( clk ), .D ( signal_24498 ), .Q ( signal_24499 ) ) ;
    buf_clk cell_9814 ( .C ( clk ), .D ( signal_24506 ), .Q ( signal_24507 ) ) ;
    buf_clk cell_9822 ( .C ( clk ), .D ( signal_24514 ), .Q ( signal_24515 ) ) ;
    buf_clk cell_9828 ( .C ( clk ), .D ( signal_24520 ), .Q ( signal_24521 ) ) ;
    buf_clk cell_9834 ( .C ( clk ), .D ( signal_24526 ), .Q ( signal_24527 ) ) ;
    buf_clk cell_9840 ( .C ( clk ), .D ( signal_24532 ), .Q ( signal_24533 ) ) ;
    buf_clk cell_9846 ( .C ( clk ), .D ( signal_24538 ), .Q ( signal_24539 ) ) ;
    buf_clk cell_9852 ( .C ( clk ), .D ( signal_24544 ), .Q ( signal_24545 ) ) ;
    buf_clk cell_9856 ( .C ( clk ), .D ( signal_24548 ), .Q ( signal_24549 ) ) ;
    buf_clk cell_9860 ( .C ( clk ), .D ( signal_24552 ), .Q ( signal_24553 ) ) ;
    buf_clk cell_9864 ( .C ( clk ), .D ( signal_24556 ), .Q ( signal_24557 ) ) ;
    buf_clk cell_9868 ( .C ( clk ), .D ( signal_24560 ), .Q ( signal_24561 ) ) ;
    buf_clk cell_9872 ( .C ( clk ), .D ( signal_24564 ), .Q ( signal_24565 ) ) ;
    buf_clk cell_9902 ( .C ( clk ), .D ( signal_24594 ), .Q ( signal_24595 ) ) ;
    buf_clk cell_9922 ( .C ( clk ), .D ( signal_24614 ), .Q ( signal_24615 ) ) ;
    buf_clk cell_9942 ( .C ( clk ), .D ( signal_24634 ), .Q ( signal_24635 ) ) ;
    buf_clk cell_9962 ( .C ( clk ), .D ( signal_24654 ), .Q ( signal_24655 ) ) ;
    buf_clk cell_9982 ( .C ( clk ), .D ( signal_24674 ), .Q ( signal_24675 ) ) ;
    buf_clk cell_9988 ( .C ( clk ), .D ( signal_24680 ), .Q ( signal_24681 ) ) ;
    buf_clk cell_9996 ( .C ( clk ), .D ( signal_24688 ), .Q ( signal_24689 ) ) ;
    buf_clk cell_10004 ( .C ( clk ), .D ( signal_24696 ), .Q ( signal_24697 ) ) ;
    buf_clk cell_10012 ( .C ( clk ), .D ( signal_24704 ), .Q ( signal_24705 ) ) ;
    buf_clk cell_10020 ( .C ( clk ), .D ( signal_24712 ), .Q ( signal_24713 ) ) ;
    buf_clk cell_10032 ( .C ( clk ), .D ( signal_24724 ), .Q ( signal_24725 ) ) ;
    buf_clk cell_10044 ( .C ( clk ), .D ( signal_24736 ), .Q ( signal_24737 ) ) ;
    buf_clk cell_10056 ( .C ( clk ), .D ( signal_24748 ), .Q ( signal_24749 ) ) ;
    buf_clk cell_10068 ( .C ( clk ), .D ( signal_24760 ), .Q ( signal_24761 ) ) ;
    buf_clk cell_10080 ( .C ( clk ), .D ( signal_24772 ), .Q ( signal_24773 ) ) ;
    buf_clk cell_10092 ( .C ( clk ), .D ( signal_24784 ), .Q ( signal_24785 ) ) ;
    buf_clk cell_10106 ( .C ( clk ), .D ( signal_24798 ), .Q ( signal_24799 ) ) ;
    buf_clk cell_10120 ( .C ( clk ), .D ( signal_24812 ), .Q ( signal_24813 ) ) ;
    buf_clk cell_10134 ( .C ( clk ), .D ( signal_24826 ), .Q ( signal_24827 ) ) ;
    buf_clk cell_10148 ( .C ( clk ), .D ( signal_24840 ), .Q ( signal_24841 ) ) ;
    buf_clk cell_10160 ( .C ( clk ), .D ( signal_24852 ), .Q ( signal_24853 ) ) ;
    buf_clk cell_10174 ( .C ( clk ), .D ( signal_24866 ), .Q ( signal_24867 ) ) ;
    buf_clk cell_10188 ( .C ( clk ), .D ( signal_24880 ), .Q ( signal_24881 ) ) ;
    buf_clk cell_10202 ( .C ( clk ), .D ( signal_24894 ), .Q ( signal_24895 ) ) ;
    buf_clk cell_10216 ( .C ( clk ), .D ( signal_24908 ), .Q ( signal_24909 ) ) ;

    /* cells in depth 25 */
    buf_clk cell_9791 ( .C ( clk ), .D ( signal_24483 ), .Q ( signal_24484 ) ) ;
    buf_clk cell_9799 ( .C ( clk ), .D ( signal_24491 ), .Q ( signal_24492 ) ) ;
    buf_clk cell_9807 ( .C ( clk ), .D ( signal_24499 ), .Q ( signal_24500 ) ) ;
    buf_clk cell_9815 ( .C ( clk ), .D ( signal_24507 ), .Q ( signal_24508 ) ) ;
    buf_clk cell_9823 ( .C ( clk ), .D ( signal_24515 ), .Q ( signal_24516 ) ) ;
    buf_clk cell_9829 ( .C ( clk ), .D ( signal_24521 ), .Q ( signal_24522 ) ) ;
    buf_clk cell_9835 ( .C ( clk ), .D ( signal_24527 ), .Q ( signal_24528 ) ) ;
    buf_clk cell_9841 ( .C ( clk ), .D ( signal_24533 ), .Q ( signal_24534 ) ) ;
    buf_clk cell_9847 ( .C ( clk ), .D ( signal_24539 ), .Q ( signal_24540 ) ) ;
    buf_clk cell_9853 ( .C ( clk ), .D ( signal_24545 ), .Q ( signal_24546 ) ) ;
    buf_clk cell_9857 ( .C ( clk ), .D ( signal_24549 ), .Q ( signal_24550 ) ) ;
    buf_clk cell_9861 ( .C ( clk ), .D ( signal_24553 ), .Q ( signal_24554 ) ) ;
    buf_clk cell_9865 ( .C ( clk ), .D ( signal_24557 ), .Q ( signal_24558 ) ) ;
    buf_clk cell_9869 ( .C ( clk ), .D ( signal_24561 ), .Q ( signal_24562 ) ) ;
    buf_clk cell_9873 ( .C ( clk ), .D ( signal_24565 ), .Q ( signal_24566 ) ) ;
    buf_clk cell_9875 ( .C ( clk ), .D ( signal_2373 ), .Q ( signal_24568 ) ) ;
    buf_clk cell_9877 ( .C ( clk ), .D ( signal_8148 ), .Q ( signal_24570 ) ) ;
    buf_clk cell_9879 ( .C ( clk ), .D ( signal_8149 ), .Q ( signal_24572 ) ) ;
    buf_clk cell_9881 ( .C ( clk ), .D ( signal_8150 ), .Q ( signal_24574 ) ) ;
    buf_clk cell_9883 ( .C ( clk ), .D ( signal_8151 ), .Q ( signal_24576 ) ) ;
    buf_clk cell_9903 ( .C ( clk ), .D ( signal_24595 ), .Q ( signal_24596 ) ) ;
    buf_clk cell_9923 ( .C ( clk ), .D ( signal_24615 ), .Q ( signal_24616 ) ) ;
    buf_clk cell_9943 ( .C ( clk ), .D ( signal_24635 ), .Q ( signal_24636 ) ) ;
    buf_clk cell_9963 ( .C ( clk ), .D ( signal_24655 ), .Q ( signal_24656 ) ) ;
    buf_clk cell_9983 ( .C ( clk ), .D ( signal_24675 ), .Q ( signal_24676 ) ) ;
    buf_clk cell_9989 ( .C ( clk ), .D ( signal_24681 ), .Q ( signal_24682 ) ) ;
    buf_clk cell_9997 ( .C ( clk ), .D ( signal_24689 ), .Q ( signal_24690 ) ) ;
    buf_clk cell_10005 ( .C ( clk ), .D ( signal_24697 ), .Q ( signal_24698 ) ) ;
    buf_clk cell_10013 ( .C ( clk ), .D ( signal_24705 ), .Q ( signal_24706 ) ) ;
    buf_clk cell_10021 ( .C ( clk ), .D ( signal_24713 ), .Q ( signal_24714 ) ) ;
    buf_clk cell_10033 ( .C ( clk ), .D ( signal_24725 ), .Q ( signal_24726 ) ) ;
    buf_clk cell_10045 ( .C ( clk ), .D ( signal_24737 ), .Q ( signal_24738 ) ) ;
    buf_clk cell_10057 ( .C ( clk ), .D ( signal_24749 ), .Q ( signal_24750 ) ) ;
    buf_clk cell_10069 ( .C ( clk ), .D ( signal_24761 ), .Q ( signal_24762 ) ) ;
    buf_clk cell_10081 ( .C ( clk ), .D ( signal_24773 ), .Q ( signal_24774 ) ) ;
    buf_clk cell_10093 ( .C ( clk ), .D ( signal_24785 ), .Q ( signal_24786 ) ) ;
    buf_clk cell_10107 ( .C ( clk ), .D ( signal_24799 ), .Q ( signal_24800 ) ) ;
    buf_clk cell_10121 ( .C ( clk ), .D ( signal_24813 ), .Q ( signal_24814 ) ) ;
    buf_clk cell_10135 ( .C ( clk ), .D ( signal_24827 ), .Q ( signal_24828 ) ) ;
    buf_clk cell_10149 ( .C ( clk ), .D ( signal_24841 ), .Q ( signal_24842 ) ) ;
    buf_clk cell_10161 ( .C ( clk ), .D ( signal_24853 ), .Q ( signal_24854 ) ) ;
    buf_clk cell_10175 ( .C ( clk ), .D ( signal_24867 ), .Q ( signal_24868 ) ) ;
    buf_clk cell_10189 ( .C ( clk ), .D ( signal_24881 ), .Q ( signal_24882 ) ) ;
    buf_clk cell_10203 ( .C ( clk ), .D ( signal_24895 ), .Q ( signal_24896 ) ) ;
    buf_clk cell_10217 ( .C ( clk ), .D ( signal_24909 ), .Q ( signal_24910 ) ) ;

    /* cells in depth 26 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2355 ( .a ({signal_24117, signal_24111, signal_24105, signal_24099, signal_24093}), .b ({signal_8099, signal_8098, signal_8097, signal_8096, signal_2360}), .clk ( clk ), .r ({Fresh[8629], Fresh[8628], Fresh[8627], Fresh[8626], Fresh[8625], Fresh[8624], Fresh[8623], Fresh[8622], Fresh[8621], Fresh[8620]}), .c ({signal_8139, signal_8138, signal_8137, signal_8136, signal_2370}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2356 ( .a ({signal_24167, signal_24157, signal_24147, signal_24137, signal_24127}), .b ({signal_8107, signal_8106, signal_8105, signal_8104, signal_2362}), .clk ( clk ), .r ({Fresh[8639], Fresh[8638], Fresh[8637], Fresh[8636], Fresh[8635], Fresh[8634], Fresh[8633], Fresh[8632], Fresh[8631], Fresh[8630]}), .c ({signal_8143, signal_8142, signal_8141, signal_8140, signal_2371}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2362 ( .a ({signal_24197, signal_24191, signal_24185, signal_24179, signal_24173}), .b ({signal_8131, signal_8130, signal_8129, signal_8128, signal_2368}), .clk ( clk ), .r ({Fresh[8649], Fresh[8648], Fresh[8647], Fresh[8646], Fresh[8645], Fresh[8644], Fresh[8643], Fresh[8642], Fresh[8641], Fresh[8640]}), .c ({signal_8167, signal_8166, signal_8165, signal_8164, signal_2377}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2363 ( .a ({signal_24247, signal_24237, signal_24227, signal_24217, signal_24207}), .b ({signal_8135, signal_8134, signal_8133, signal_8132, signal_2369}), .clk ( clk ), .r ({Fresh[8659], Fresh[8658], Fresh[8657], Fresh[8656], Fresh[8655], Fresh[8654], Fresh[8653], Fresh[8652], Fresh[8651], Fresh[8650]}), .c ({signal_8171, signal_8170, signal_8169, signal_8168, signal_2378}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2365 ( .a ({signal_8171, signal_8170, signal_8169, signal_8168, signal_2378}), .b ({signal_8179, signal_8178, signal_8177, signal_8176, signal_26}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2368 ( .a ({signal_24327, signal_24311, signal_24295, signal_24279, signal_24263}), .b ({signal_8147, signal_8146, signal_8145, signal_8144, signal_2372}), .clk ( clk ), .r ({Fresh[8669], Fresh[8668], Fresh[8667], Fresh[8666], Fresh[8665], Fresh[8664], Fresh[8663], Fresh[8662], Fresh[8661], Fresh[8660]}), .c ({signal_8191, signal_8190, signal_8189, signal_8188, signal_2381}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2369 ( .a ({signal_24417, signal_24399, signal_24381, signal_24363, signal_24345}), .b ({signal_8155, signal_8154, signal_8153, signal_8152, signal_2374}), .clk ( clk ), .r ({Fresh[8679], Fresh[8678], Fresh[8677], Fresh[8676], Fresh[8675], Fresh[8674], Fresh[8673], Fresh[8672], Fresh[8671], Fresh[8670]}), .c ({signal_8195, signal_8194, signal_8193, signal_8192, signal_2382}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2370 ( .a ({signal_24437, signal_24433, signal_24429, signal_24425, signal_24421}), .b ({signal_8159, signal_8158, signal_8157, signal_8156, signal_2375}), .clk ( clk ), .r ({Fresh[8689], Fresh[8688], Fresh[8687], Fresh[8686], Fresh[8685], Fresh[8684], Fresh[8683], Fresh[8682], Fresh[8681], Fresh[8680]}), .c ({signal_8199, signal_8198, signal_8197, signal_8196, signal_2383}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2371 ( .a ({signal_24477, signal_24469, signal_24461, signal_24453, signal_24445}), .b ({signal_8163, signal_8162, signal_8161, signal_8160, signal_2376}), .clk ( clk ), .r ({Fresh[8699], Fresh[8698], Fresh[8697], Fresh[8696], Fresh[8695], Fresh[8694], Fresh[8693], Fresh[8692], Fresh[8691], Fresh[8690]}), .c ({signal_8203, signal_8202, signal_8201, signal_8200, signal_2384}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2374 ( .a ({signal_8199, signal_8198, signal_8197, signal_8196, signal_2383}), .b ({signal_8215, signal_8214, signal_8213, signal_8212, signal_28}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2375 ( .a ({signal_8203, signal_8202, signal_8201, signal_8200, signal_2384}), .b ({signal_8219, signal_8218, signal_8217, signal_8216, signal_29}) ) ;
    buf_clk cell_9792 ( .C ( clk ), .D ( signal_24484 ), .Q ( signal_24485 ) ) ;
    buf_clk cell_9800 ( .C ( clk ), .D ( signal_24492 ), .Q ( signal_24493 ) ) ;
    buf_clk cell_9808 ( .C ( clk ), .D ( signal_24500 ), .Q ( signal_24501 ) ) ;
    buf_clk cell_9816 ( .C ( clk ), .D ( signal_24508 ), .Q ( signal_24509 ) ) ;
    buf_clk cell_9824 ( .C ( clk ), .D ( signal_24516 ), .Q ( signal_24517 ) ) ;
    buf_clk cell_9830 ( .C ( clk ), .D ( signal_24522 ), .Q ( signal_24523 ) ) ;
    buf_clk cell_9836 ( .C ( clk ), .D ( signal_24528 ), .Q ( signal_24529 ) ) ;
    buf_clk cell_9842 ( .C ( clk ), .D ( signal_24534 ), .Q ( signal_24535 ) ) ;
    buf_clk cell_9848 ( .C ( clk ), .D ( signal_24540 ), .Q ( signal_24541 ) ) ;
    buf_clk cell_9854 ( .C ( clk ), .D ( signal_24546 ), .Q ( signal_24547 ) ) ;
    buf_clk cell_9858 ( .C ( clk ), .D ( signal_24550 ), .Q ( signal_24551 ) ) ;
    buf_clk cell_9862 ( .C ( clk ), .D ( signal_24554 ), .Q ( signal_24555 ) ) ;
    buf_clk cell_9866 ( .C ( clk ), .D ( signal_24558 ), .Q ( signal_24559 ) ) ;
    buf_clk cell_9870 ( .C ( clk ), .D ( signal_24562 ), .Q ( signal_24563 ) ) ;
    buf_clk cell_9874 ( .C ( clk ), .D ( signal_24566 ), .Q ( signal_24567 ) ) ;
    buf_clk cell_9876 ( .C ( clk ), .D ( signal_24568 ), .Q ( signal_24569 ) ) ;
    buf_clk cell_9878 ( .C ( clk ), .D ( signal_24570 ), .Q ( signal_24571 ) ) ;
    buf_clk cell_9880 ( .C ( clk ), .D ( signal_24572 ), .Q ( signal_24573 ) ) ;
    buf_clk cell_9882 ( .C ( clk ), .D ( signal_24574 ), .Q ( signal_24575 ) ) ;
    buf_clk cell_9884 ( .C ( clk ), .D ( signal_24576 ), .Q ( signal_24577 ) ) ;
    buf_clk cell_9904 ( .C ( clk ), .D ( signal_24596 ), .Q ( signal_24597 ) ) ;
    buf_clk cell_9924 ( .C ( clk ), .D ( signal_24616 ), .Q ( signal_24617 ) ) ;
    buf_clk cell_9944 ( .C ( clk ), .D ( signal_24636 ), .Q ( signal_24637 ) ) ;
    buf_clk cell_9964 ( .C ( clk ), .D ( signal_24656 ), .Q ( signal_24657 ) ) ;
    buf_clk cell_9984 ( .C ( clk ), .D ( signal_24676 ), .Q ( signal_24677 ) ) ;
    buf_clk cell_9990 ( .C ( clk ), .D ( signal_24682 ), .Q ( signal_24683 ) ) ;
    buf_clk cell_9998 ( .C ( clk ), .D ( signal_24690 ), .Q ( signal_24691 ) ) ;
    buf_clk cell_10006 ( .C ( clk ), .D ( signal_24698 ), .Q ( signal_24699 ) ) ;
    buf_clk cell_10014 ( .C ( clk ), .D ( signal_24706 ), .Q ( signal_24707 ) ) ;
    buf_clk cell_10022 ( .C ( clk ), .D ( signal_24714 ), .Q ( signal_24715 ) ) ;
    buf_clk cell_10034 ( .C ( clk ), .D ( signal_24726 ), .Q ( signal_24727 ) ) ;
    buf_clk cell_10046 ( .C ( clk ), .D ( signal_24738 ), .Q ( signal_24739 ) ) ;
    buf_clk cell_10058 ( .C ( clk ), .D ( signal_24750 ), .Q ( signal_24751 ) ) ;
    buf_clk cell_10070 ( .C ( clk ), .D ( signal_24762 ), .Q ( signal_24763 ) ) ;
    buf_clk cell_10082 ( .C ( clk ), .D ( signal_24774 ), .Q ( signal_24775 ) ) ;
    buf_clk cell_10094 ( .C ( clk ), .D ( signal_24786 ), .Q ( signal_24787 ) ) ;
    buf_clk cell_10108 ( .C ( clk ), .D ( signal_24800 ), .Q ( signal_24801 ) ) ;
    buf_clk cell_10122 ( .C ( clk ), .D ( signal_24814 ), .Q ( signal_24815 ) ) ;
    buf_clk cell_10136 ( .C ( clk ), .D ( signal_24828 ), .Q ( signal_24829 ) ) ;
    buf_clk cell_10150 ( .C ( clk ), .D ( signal_24842 ), .Q ( signal_24843 ) ) ;
    buf_clk cell_10162 ( .C ( clk ), .D ( signal_24854 ), .Q ( signal_24855 ) ) ;
    buf_clk cell_10176 ( .C ( clk ), .D ( signal_24868 ), .Q ( signal_24869 ) ) ;
    buf_clk cell_10190 ( .C ( clk ), .D ( signal_24882 ), .Q ( signal_24883 ) ) ;
    buf_clk cell_10204 ( .C ( clk ), .D ( signal_24896 ), .Q ( signal_24897 ) ) ;
    buf_clk cell_10218 ( .C ( clk ), .D ( signal_24910 ), .Q ( signal_24911 ) ) ;

    /* cells in depth 27 */
    buf_clk cell_9991 ( .C ( clk ), .D ( signal_24683 ), .Q ( signal_24684 ) ) ;
    buf_clk cell_9999 ( .C ( clk ), .D ( signal_24691 ), .Q ( signal_24692 ) ) ;
    buf_clk cell_10007 ( .C ( clk ), .D ( signal_24699 ), .Q ( signal_24700 ) ) ;
    buf_clk cell_10015 ( .C ( clk ), .D ( signal_24707 ), .Q ( signal_24708 ) ) ;
    buf_clk cell_10023 ( .C ( clk ), .D ( signal_24715 ), .Q ( signal_24716 ) ) ;
    buf_clk cell_10035 ( .C ( clk ), .D ( signal_24727 ), .Q ( signal_24728 ) ) ;
    buf_clk cell_10047 ( .C ( clk ), .D ( signal_24739 ), .Q ( signal_24740 ) ) ;
    buf_clk cell_10059 ( .C ( clk ), .D ( signal_24751 ), .Q ( signal_24752 ) ) ;
    buf_clk cell_10071 ( .C ( clk ), .D ( signal_24763 ), .Q ( signal_24764 ) ) ;
    buf_clk cell_10083 ( .C ( clk ), .D ( signal_24775 ), .Q ( signal_24776 ) ) ;
    buf_clk cell_10095 ( .C ( clk ), .D ( signal_24787 ), .Q ( signal_24788 ) ) ;
    buf_clk cell_10109 ( .C ( clk ), .D ( signal_24801 ), .Q ( signal_24802 ) ) ;
    buf_clk cell_10123 ( .C ( clk ), .D ( signal_24815 ), .Q ( signal_24816 ) ) ;
    buf_clk cell_10137 ( .C ( clk ), .D ( signal_24829 ), .Q ( signal_24830 ) ) ;
    buf_clk cell_10151 ( .C ( clk ), .D ( signal_24843 ), .Q ( signal_24844 ) ) ;
    buf_clk cell_10163 ( .C ( clk ), .D ( signal_24855 ), .Q ( signal_24856 ) ) ;
    buf_clk cell_10177 ( .C ( clk ), .D ( signal_24869 ), .Q ( signal_24870 ) ) ;
    buf_clk cell_10191 ( .C ( clk ), .D ( signal_24883 ), .Q ( signal_24884 ) ) ;
    buf_clk cell_10205 ( .C ( clk ), .D ( signal_24897 ), .Q ( signal_24898 ) ) ;
    buf_clk cell_10219 ( .C ( clk ), .D ( signal_24911 ), .Q ( signal_24912 ) ) ;
    buf_clk cell_10305 ( .C ( clk ), .D ( signal_26 ), .Q ( signal_24998 ) ) ;
    buf_clk cell_10313 ( .C ( clk ), .D ( signal_8176 ), .Q ( signal_25006 ) ) ;
    buf_clk cell_10321 ( .C ( clk ), .D ( signal_8177 ), .Q ( signal_25014 ) ) ;
    buf_clk cell_10329 ( .C ( clk ), .D ( signal_8178 ), .Q ( signal_25022 ) ) ;
    buf_clk cell_10337 ( .C ( clk ), .D ( signal_8179 ), .Q ( signal_25030 ) ) ;
    buf_clk cell_10345 ( .C ( clk ), .D ( signal_28 ), .Q ( signal_25038 ) ) ;
    buf_clk cell_10353 ( .C ( clk ), .D ( signal_8212 ), .Q ( signal_25046 ) ) ;
    buf_clk cell_10361 ( .C ( clk ), .D ( signal_8213 ), .Q ( signal_25054 ) ) ;
    buf_clk cell_10369 ( .C ( clk ), .D ( signal_8214 ), .Q ( signal_25062 ) ) ;
    buf_clk cell_10377 ( .C ( clk ), .D ( signal_8215 ), .Q ( signal_25070 ) ) ;
    buf_clk cell_10385 ( .C ( clk ), .D ( signal_29 ), .Q ( signal_25078 ) ) ;
    buf_clk cell_10393 ( .C ( clk ), .D ( signal_8216 ), .Q ( signal_25086 ) ) ;
    buf_clk cell_10401 ( .C ( clk ), .D ( signal_8217 ), .Q ( signal_25094 ) ) ;
    buf_clk cell_10409 ( .C ( clk ), .D ( signal_8218 ), .Q ( signal_25102 ) ) ;
    buf_clk cell_10417 ( .C ( clk ), .D ( signal_8219 ), .Q ( signal_25110 ) ) ;

    /* cells in depth 28 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2364 ( .a ({signal_24517, signal_24509, signal_24501, signal_24493, signal_24485}), .b ({signal_8139, signal_8138, signal_8137, signal_8136, signal_2370}), .clk ( clk ), .r ({Fresh[8709], Fresh[8708], Fresh[8707], Fresh[8706], Fresh[8705], Fresh[8704], Fresh[8703], Fresh[8702], Fresh[8701], Fresh[8700]}), .c ({signal_8175, signal_8174, signal_8173, signal_8172, signal_2379}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2366 ( .a ({signal_8175, signal_8174, signal_8173, signal_8172, signal_2379}), .b ({signal_8183, signal_8182, signal_8181, signal_8180, signal_23}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2367 ( .a ({signal_24547, signal_24541, signal_24535, signal_24529, signal_24523}), .b ({signal_8143, signal_8142, signal_8141, signal_8140, signal_2371}), .clk ( clk ), .r ({Fresh[8719], Fresh[8718], Fresh[8717], Fresh[8716], Fresh[8715], Fresh[8714], Fresh[8713], Fresh[8712], Fresh[8711], Fresh[8710]}), .c ({signal_8187, signal_8186, signal_8185, signal_8184, signal_2380}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2372 ( .a ({signal_24567, signal_24563, signal_24559, signal_24555, signal_24551}), .b ({signal_8167, signal_8166, signal_8165, signal_8164, signal_2377}), .clk ( clk ), .r ({Fresh[8729], Fresh[8728], Fresh[8727], Fresh[8726], Fresh[8725], Fresh[8724], Fresh[8723], Fresh[8722], Fresh[8721], Fresh[8720]}), .c ({signal_8207, signal_8206, signal_8205, signal_8204, signal_2385}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2373 ( .a ({signal_8187, signal_8186, signal_8185, signal_8184, signal_2380}), .b ({signal_8211, signal_8210, signal_8209, signal_8208, signal_30}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2376 ( .a ({signal_8207, signal_8206, signal_8205, signal_8204, signal_2385}), .b ({signal_8223, signal_8222, signal_8221, signal_8220, signal_24}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2377 ( .a ({signal_24577, signal_24575, signal_24573, signal_24571, signal_24569}), .b ({signal_8191, signal_8190, signal_8189, signal_8188, signal_2381}), .clk ( clk ), .r ({Fresh[8739], Fresh[8738], Fresh[8737], Fresh[8736], Fresh[8735], Fresh[8734], Fresh[8733], Fresh[8732], Fresh[8731], Fresh[8730]}), .c ({signal_8227, signal_8226, signal_8225, signal_8224, signal_2386}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2378 ( .a ({signal_24677, signal_24657, signal_24637, signal_24617, signal_24597}), .b ({signal_8195, signal_8194, signal_8193, signal_8192, signal_2382}), .clk ( clk ), .r ({Fresh[8749], Fresh[8748], Fresh[8747], Fresh[8746], Fresh[8745], Fresh[8744], Fresh[8743], Fresh[8742], Fresh[8741], Fresh[8740]}), .c ({signal_8231, signal_8230, signal_8229, signal_8228, signal_2387}) ) ;
    buf_clk cell_9992 ( .C ( clk ), .D ( signal_24684 ), .Q ( signal_24685 ) ) ;
    buf_clk cell_10000 ( .C ( clk ), .D ( signal_24692 ), .Q ( signal_24693 ) ) ;
    buf_clk cell_10008 ( .C ( clk ), .D ( signal_24700 ), .Q ( signal_24701 ) ) ;
    buf_clk cell_10016 ( .C ( clk ), .D ( signal_24708 ), .Q ( signal_24709 ) ) ;
    buf_clk cell_10024 ( .C ( clk ), .D ( signal_24716 ), .Q ( signal_24717 ) ) ;
    buf_clk cell_10036 ( .C ( clk ), .D ( signal_24728 ), .Q ( signal_24729 ) ) ;
    buf_clk cell_10048 ( .C ( clk ), .D ( signal_24740 ), .Q ( signal_24741 ) ) ;
    buf_clk cell_10060 ( .C ( clk ), .D ( signal_24752 ), .Q ( signal_24753 ) ) ;
    buf_clk cell_10072 ( .C ( clk ), .D ( signal_24764 ), .Q ( signal_24765 ) ) ;
    buf_clk cell_10084 ( .C ( clk ), .D ( signal_24776 ), .Q ( signal_24777 ) ) ;
    buf_clk cell_10096 ( .C ( clk ), .D ( signal_24788 ), .Q ( signal_24789 ) ) ;
    buf_clk cell_10110 ( .C ( clk ), .D ( signal_24802 ), .Q ( signal_24803 ) ) ;
    buf_clk cell_10124 ( .C ( clk ), .D ( signal_24816 ), .Q ( signal_24817 ) ) ;
    buf_clk cell_10138 ( .C ( clk ), .D ( signal_24830 ), .Q ( signal_24831 ) ) ;
    buf_clk cell_10152 ( .C ( clk ), .D ( signal_24844 ), .Q ( signal_24845 ) ) ;
    buf_clk cell_10164 ( .C ( clk ), .D ( signal_24856 ), .Q ( signal_24857 ) ) ;
    buf_clk cell_10178 ( .C ( clk ), .D ( signal_24870 ), .Q ( signal_24871 ) ) ;
    buf_clk cell_10192 ( .C ( clk ), .D ( signal_24884 ), .Q ( signal_24885 ) ) ;
    buf_clk cell_10206 ( .C ( clk ), .D ( signal_24898 ), .Q ( signal_24899 ) ) ;
    buf_clk cell_10220 ( .C ( clk ), .D ( signal_24912 ), .Q ( signal_24913 ) ) ;
    buf_clk cell_10306 ( .C ( clk ), .D ( signal_24998 ), .Q ( signal_24999 ) ) ;
    buf_clk cell_10314 ( .C ( clk ), .D ( signal_25006 ), .Q ( signal_25007 ) ) ;
    buf_clk cell_10322 ( .C ( clk ), .D ( signal_25014 ), .Q ( signal_25015 ) ) ;
    buf_clk cell_10330 ( .C ( clk ), .D ( signal_25022 ), .Q ( signal_25023 ) ) ;
    buf_clk cell_10338 ( .C ( clk ), .D ( signal_25030 ), .Q ( signal_25031 ) ) ;
    buf_clk cell_10346 ( .C ( clk ), .D ( signal_25038 ), .Q ( signal_25039 ) ) ;
    buf_clk cell_10354 ( .C ( clk ), .D ( signal_25046 ), .Q ( signal_25047 ) ) ;
    buf_clk cell_10362 ( .C ( clk ), .D ( signal_25054 ), .Q ( signal_25055 ) ) ;
    buf_clk cell_10370 ( .C ( clk ), .D ( signal_25062 ), .Q ( signal_25063 ) ) ;
    buf_clk cell_10378 ( .C ( clk ), .D ( signal_25070 ), .Q ( signal_25071 ) ) ;
    buf_clk cell_10386 ( .C ( clk ), .D ( signal_25078 ), .Q ( signal_25079 ) ) ;
    buf_clk cell_10394 ( .C ( clk ), .D ( signal_25086 ), .Q ( signal_25087 ) ) ;
    buf_clk cell_10402 ( .C ( clk ), .D ( signal_25094 ), .Q ( signal_25095 ) ) ;
    buf_clk cell_10410 ( .C ( clk ), .D ( signal_25102 ), .Q ( signal_25103 ) ) ;
    buf_clk cell_10418 ( .C ( clk ), .D ( signal_25110 ), .Q ( signal_25111 ) ) ;

    /* cells in depth 29 */
    buf_clk cell_10097 ( .C ( clk ), .D ( signal_24789 ), .Q ( signal_24790 ) ) ;
    buf_clk cell_10111 ( .C ( clk ), .D ( signal_24803 ), .Q ( signal_24804 ) ) ;
    buf_clk cell_10125 ( .C ( clk ), .D ( signal_24817 ), .Q ( signal_24818 ) ) ;
    buf_clk cell_10139 ( .C ( clk ), .D ( signal_24831 ), .Q ( signal_24832 ) ) ;
    buf_clk cell_10153 ( .C ( clk ), .D ( signal_24845 ), .Q ( signal_24846 ) ) ;
    buf_clk cell_10165 ( .C ( clk ), .D ( signal_24857 ), .Q ( signal_24858 ) ) ;
    buf_clk cell_10179 ( .C ( clk ), .D ( signal_24871 ), .Q ( signal_24872 ) ) ;
    buf_clk cell_10193 ( .C ( clk ), .D ( signal_24885 ), .Q ( signal_24886 ) ) ;
    buf_clk cell_10207 ( .C ( clk ), .D ( signal_24899 ), .Q ( signal_24900 ) ) ;
    buf_clk cell_10221 ( .C ( clk ), .D ( signal_24913 ), .Q ( signal_24914 ) ) ;
    buf_clk cell_10225 ( .C ( clk ), .D ( signal_23 ), .Q ( signal_24918 ) ) ;
    buf_clk cell_10231 ( .C ( clk ), .D ( signal_8180 ), .Q ( signal_24924 ) ) ;
    buf_clk cell_10237 ( .C ( clk ), .D ( signal_8181 ), .Q ( signal_24930 ) ) ;
    buf_clk cell_10243 ( .C ( clk ), .D ( signal_8182 ), .Q ( signal_24936 ) ) ;
    buf_clk cell_10249 ( .C ( clk ), .D ( signal_8183 ), .Q ( signal_24942 ) ) ;
    buf_clk cell_10255 ( .C ( clk ), .D ( signal_24 ), .Q ( signal_24948 ) ) ;
    buf_clk cell_10261 ( .C ( clk ), .D ( signal_8220 ), .Q ( signal_24954 ) ) ;
    buf_clk cell_10267 ( .C ( clk ), .D ( signal_8221 ), .Q ( signal_24960 ) ) ;
    buf_clk cell_10273 ( .C ( clk ), .D ( signal_8222 ), .Q ( signal_24966 ) ) ;
    buf_clk cell_10279 ( .C ( clk ), .D ( signal_8223 ), .Q ( signal_24972 ) ) ;
    buf_clk cell_10307 ( .C ( clk ), .D ( signal_24999 ), .Q ( signal_25000 ) ) ;
    buf_clk cell_10315 ( .C ( clk ), .D ( signal_25007 ), .Q ( signal_25008 ) ) ;
    buf_clk cell_10323 ( .C ( clk ), .D ( signal_25015 ), .Q ( signal_25016 ) ) ;
    buf_clk cell_10331 ( .C ( clk ), .D ( signal_25023 ), .Q ( signal_25024 ) ) ;
    buf_clk cell_10339 ( .C ( clk ), .D ( signal_25031 ), .Q ( signal_25032 ) ) ;
    buf_clk cell_10347 ( .C ( clk ), .D ( signal_25039 ), .Q ( signal_25040 ) ) ;
    buf_clk cell_10355 ( .C ( clk ), .D ( signal_25047 ), .Q ( signal_25048 ) ) ;
    buf_clk cell_10363 ( .C ( clk ), .D ( signal_25055 ), .Q ( signal_25056 ) ) ;
    buf_clk cell_10371 ( .C ( clk ), .D ( signal_25063 ), .Q ( signal_25064 ) ) ;
    buf_clk cell_10379 ( .C ( clk ), .D ( signal_25071 ), .Q ( signal_25072 ) ) ;
    buf_clk cell_10387 ( .C ( clk ), .D ( signal_25079 ), .Q ( signal_25080 ) ) ;
    buf_clk cell_10395 ( .C ( clk ), .D ( signal_25087 ), .Q ( signal_25088 ) ) ;
    buf_clk cell_10403 ( .C ( clk ), .D ( signal_25095 ), .Q ( signal_25096 ) ) ;
    buf_clk cell_10411 ( .C ( clk ), .D ( signal_25103 ), .Q ( signal_25104 ) ) ;
    buf_clk cell_10419 ( .C ( clk ), .D ( signal_25111 ), .Q ( signal_25112 ) ) ;
    buf_clk cell_10425 ( .C ( clk ), .D ( signal_30 ), .Q ( signal_25118 ) ) ;
    buf_clk cell_10431 ( .C ( clk ), .D ( signal_8208 ), .Q ( signal_25124 ) ) ;
    buf_clk cell_10437 ( .C ( clk ), .D ( signal_8209 ), .Q ( signal_25130 ) ) ;
    buf_clk cell_10443 ( .C ( clk ), .D ( signal_8210 ), .Q ( signal_25136 ) ) ;
    buf_clk cell_10449 ( .C ( clk ), .D ( signal_8211 ), .Q ( signal_25142 ) ) ;

    /* cells in depth 30 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2379 ( .a ({signal_24717, signal_24709, signal_24701, signal_24693, signal_24685}), .b ({signal_8227, signal_8226, signal_8225, signal_8224, signal_2386}), .clk ( clk ), .r ({Fresh[8759], Fresh[8758], Fresh[8757], Fresh[8756], Fresh[8755], Fresh[8754], Fresh[8753], Fresh[8752], Fresh[8751], Fresh[8750]}), .c ({signal_8235, signal_8234, signal_8233, signal_8232, signal_2388}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2380 ( .a ({signal_24777, signal_24765, signal_24753, signal_24741, signal_24729}), .b ({signal_8231, signal_8230, signal_8229, signal_8228, signal_2387}), .clk ( clk ), .r ({Fresh[8769], Fresh[8768], Fresh[8767], Fresh[8766], Fresh[8765], Fresh[8764], Fresh[8763], Fresh[8762], Fresh[8761], Fresh[8760]}), .c ({signal_8239, signal_8238, signal_8237, signal_8236, signal_2389}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2381 ( .a ({signal_8235, signal_8234, signal_8233, signal_8232, signal_2388}), .b ({signal_8243, signal_8242, signal_8241, signal_8240, signal_25}) ) ;
    buf_clk cell_10098 ( .C ( clk ), .D ( signal_24790 ), .Q ( signal_24791 ) ) ;
    buf_clk cell_10112 ( .C ( clk ), .D ( signal_24804 ), .Q ( signal_24805 ) ) ;
    buf_clk cell_10126 ( .C ( clk ), .D ( signal_24818 ), .Q ( signal_24819 ) ) ;
    buf_clk cell_10140 ( .C ( clk ), .D ( signal_24832 ), .Q ( signal_24833 ) ) ;
    buf_clk cell_10154 ( .C ( clk ), .D ( signal_24846 ), .Q ( signal_24847 ) ) ;
    buf_clk cell_10166 ( .C ( clk ), .D ( signal_24858 ), .Q ( signal_24859 ) ) ;
    buf_clk cell_10180 ( .C ( clk ), .D ( signal_24872 ), .Q ( signal_24873 ) ) ;
    buf_clk cell_10194 ( .C ( clk ), .D ( signal_24886 ), .Q ( signal_24887 ) ) ;
    buf_clk cell_10208 ( .C ( clk ), .D ( signal_24900 ), .Q ( signal_24901 ) ) ;
    buf_clk cell_10222 ( .C ( clk ), .D ( signal_24914 ), .Q ( signal_24915 ) ) ;
    buf_clk cell_10226 ( .C ( clk ), .D ( signal_24918 ), .Q ( signal_24919 ) ) ;
    buf_clk cell_10232 ( .C ( clk ), .D ( signal_24924 ), .Q ( signal_24925 ) ) ;
    buf_clk cell_10238 ( .C ( clk ), .D ( signal_24930 ), .Q ( signal_24931 ) ) ;
    buf_clk cell_10244 ( .C ( clk ), .D ( signal_24936 ), .Q ( signal_24937 ) ) ;
    buf_clk cell_10250 ( .C ( clk ), .D ( signal_24942 ), .Q ( signal_24943 ) ) ;
    buf_clk cell_10256 ( .C ( clk ), .D ( signal_24948 ), .Q ( signal_24949 ) ) ;
    buf_clk cell_10262 ( .C ( clk ), .D ( signal_24954 ), .Q ( signal_24955 ) ) ;
    buf_clk cell_10268 ( .C ( clk ), .D ( signal_24960 ), .Q ( signal_24961 ) ) ;
    buf_clk cell_10274 ( .C ( clk ), .D ( signal_24966 ), .Q ( signal_24967 ) ) ;
    buf_clk cell_10280 ( .C ( clk ), .D ( signal_24972 ), .Q ( signal_24973 ) ) ;
    buf_clk cell_10308 ( .C ( clk ), .D ( signal_25000 ), .Q ( signal_25001 ) ) ;
    buf_clk cell_10316 ( .C ( clk ), .D ( signal_25008 ), .Q ( signal_25009 ) ) ;
    buf_clk cell_10324 ( .C ( clk ), .D ( signal_25016 ), .Q ( signal_25017 ) ) ;
    buf_clk cell_10332 ( .C ( clk ), .D ( signal_25024 ), .Q ( signal_25025 ) ) ;
    buf_clk cell_10340 ( .C ( clk ), .D ( signal_25032 ), .Q ( signal_25033 ) ) ;
    buf_clk cell_10348 ( .C ( clk ), .D ( signal_25040 ), .Q ( signal_25041 ) ) ;
    buf_clk cell_10356 ( .C ( clk ), .D ( signal_25048 ), .Q ( signal_25049 ) ) ;
    buf_clk cell_10364 ( .C ( clk ), .D ( signal_25056 ), .Q ( signal_25057 ) ) ;
    buf_clk cell_10372 ( .C ( clk ), .D ( signal_25064 ), .Q ( signal_25065 ) ) ;
    buf_clk cell_10380 ( .C ( clk ), .D ( signal_25072 ), .Q ( signal_25073 ) ) ;
    buf_clk cell_10388 ( .C ( clk ), .D ( signal_25080 ), .Q ( signal_25081 ) ) ;
    buf_clk cell_10396 ( .C ( clk ), .D ( signal_25088 ), .Q ( signal_25089 ) ) ;
    buf_clk cell_10404 ( .C ( clk ), .D ( signal_25096 ), .Q ( signal_25097 ) ) ;
    buf_clk cell_10412 ( .C ( clk ), .D ( signal_25104 ), .Q ( signal_25105 ) ) ;
    buf_clk cell_10420 ( .C ( clk ), .D ( signal_25112 ), .Q ( signal_25113 ) ) ;
    buf_clk cell_10426 ( .C ( clk ), .D ( signal_25118 ), .Q ( signal_25119 ) ) ;
    buf_clk cell_10432 ( .C ( clk ), .D ( signal_25124 ), .Q ( signal_25125 ) ) ;
    buf_clk cell_10438 ( .C ( clk ), .D ( signal_25130 ), .Q ( signal_25131 ) ) ;
    buf_clk cell_10444 ( .C ( clk ), .D ( signal_25136 ), .Q ( signal_25137 ) ) ;
    buf_clk cell_10450 ( .C ( clk ), .D ( signal_25142 ), .Q ( signal_25143 ) ) ;

    /* cells in depth 31 */
    buf_clk cell_10167 ( .C ( clk ), .D ( signal_24859 ), .Q ( signal_24860 ) ) ;
    buf_clk cell_10181 ( .C ( clk ), .D ( signal_24873 ), .Q ( signal_24874 ) ) ;
    buf_clk cell_10195 ( .C ( clk ), .D ( signal_24887 ), .Q ( signal_24888 ) ) ;
    buf_clk cell_10209 ( .C ( clk ), .D ( signal_24901 ), .Q ( signal_24902 ) ) ;
    buf_clk cell_10223 ( .C ( clk ), .D ( signal_24915 ), .Q ( signal_24916 ) ) ;
    buf_clk cell_10227 ( .C ( clk ), .D ( signal_24919 ), .Q ( signal_24920 ) ) ;
    buf_clk cell_10233 ( .C ( clk ), .D ( signal_24925 ), .Q ( signal_24926 ) ) ;
    buf_clk cell_10239 ( .C ( clk ), .D ( signal_24931 ), .Q ( signal_24932 ) ) ;
    buf_clk cell_10245 ( .C ( clk ), .D ( signal_24937 ), .Q ( signal_24938 ) ) ;
    buf_clk cell_10251 ( .C ( clk ), .D ( signal_24943 ), .Q ( signal_24944 ) ) ;
    buf_clk cell_10257 ( .C ( clk ), .D ( signal_24949 ), .Q ( signal_24950 ) ) ;
    buf_clk cell_10263 ( .C ( clk ), .D ( signal_24955 ), .Q ( signal_24956 ) ) ;
    buf_clk cell_10269 ( .C ( clk ), .D ( signal_24961 ), .Q ( signal_24962 ) ) ;
    buf_clk cell_10275 ( .C ( clk ), .D ( signal_24967 ), .Q ( signal_24968 ) ) ;
    buf_clk cell_10281 ( .C ( clk ), .D ( signal_24973 ), .Q ( signal_24974 ) ) ;
    buf_clk cell_10285 ( .C ( clk ), .D ( signal_25 ), .Q ( signal_24978 ) ) ;
    buf_clk cell_10289 ( .C ( clk ), .D ( signal_8240 ), .Q ( signal_24982 ) ) ;
    buf_clk cell_10293 ( .C ( clk ), .D ( signal_8241 ), .Q ( signal_24986 ) ) ;
    buf_clk cell_10297 ( .C ( clk ), .D ( signal_8242 ), .Q ( signal_24990 ) ) ;
    buf_clk cell_10301 ( .C ( clk ), .D ( signal_8243 ), .Q ( signal_24994 ) ) ;
    buf_clk cell_10309 ( .C ( clk ), .D ( signal_25001 ), .Q ( signal_25002 ) ) ;
    buf_clk cell_10317 ( .C ( clk ), .D ( signal_25009 ), .Q ( signal_25010 ) ) ;
    buf_clk cell_10325 ( .C ( clk ), .D ( signal_25017 ), .Q ( signal_25018 ) ) ;
    buf_clk cell_10333 ( .C ( clk ), .D ( signal_25025 ), .Q ( signal_25026 ) ) ;
    buf_clk cell_10341 ( .C ( clk ), .D ( signal_25033 ), .Q ( signal_25034 ) ) ;
    buf_clk cell_10349 ( .C ( clk ), .D ( signal_25041 ), .Q ( signal_25042 ) ) ;
    buf_clk cell_10357 ( .C ( clk ), .D ( signal_25049 ), .Q ( signal_25050 ) ) ;
    buf_clk cell_10365 ( .C ( clk ), .D ( signal_25057 ), .Q ( signal_25058 ) ) ;
    buf_clk cell_10373 ( .C ( clk ), .D ( signal_25065 ), .Q ( signal_25066 ) ) ;
    buf_clk cell_10381 ( .C ( clk ), .D ( signal_25073 ), .Q ( signal_25074 ) ) ;
    buf_clk cell_10389 ( .C ( clk ), .D ( signal_25081 ), .Q ( signal_25082 ) ) ;
    buf_clk cell_10397 ( .C ( clk ), .D ( signal_25089 ), .Q ( signal_25090 ) ) ;
    buf_clk cell_10405 ( .C ( clk ), .D ( signal_25097 ), .Q ( signal_25098 ) ) ;
    buf_clk cell_10413 ( .C ( clk ), .D ( signal_25105 ), .Q ( signal_25106 ) ) ;
    buf_clk cell_10421 ( .C ( clk ), .D ( signal_25113 ), .Q ( signal_25114 ) ) ;
    buf_clk cell_10427 ( .C ( clk ), .D ( signal_25119 ), .Q ( signal_25120 ) ) ;
    buf_clk cell_10433 ( .C ( clk ), .D ( signal_25125 ), .Q ( signal_25126 ) ) ;
    buf_clk cell_10439 ( .C ( clk ), .D ( signal_25131 ), .Q ( signal_25132 ) ) ;
    buf_clk cell_10445 ( .C ( clk ), .D ( signal_25137 ), .Q ( signal_25138 ) ) ;
    buf_clk cell_10451 ( .C ( clk ), .D ( signal_25143 ), .Q ( signal_25144 ) ) ;

    /* cells in depth 32 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2382 ( .a ({signal_24847, signal_24833, signal_24819, signal_24805, signal_24791}), .b ({signal_8239, signal_8238, signal_8237, signal_8236, signal_2389}), .clk ( clk ), .r ({Fresh[8779], Fresh[8778], Fresh[8777], Fresh[8776], Fresh[8775], Fresh[8774], Fresh[8773], Fresh[8772], Fresh[8771], Fresh[8770]}), .c ({signal_8247, signal_8246, signal_8245, signal_8244, signal_2390}) ) ;
    buf_clk cell_10168 ( .C ( clk ), .D ( signal_24860 ), .Q ( signal_24861 ) ) ;
    buf_clk cell_10182 ( .C ( clk ), .D ( signal_24874 ), .Q ( signal_24875 ) ) ;
    buf_clk cell_10196 ( .C ( clk ), .D ( signal_24888 ), .Q ( signal_24889 ) ) ;
    buf_clk cell_10210 ( .C ( clk ), .D ( signal_24902 ), .Q ( signal_24903 ) ) ;
    buf_clk cell_10224 ( .C ( clk ), .D ( signal_24916 ), .Q ( signal_24917 ) ) ;
    buf_clk cell_10228 ( .C ( clk ), .D ( signal_24920 ), .Q ( signal_24921 ) ) ;
    buf_clk cell_10234 ( .C ( clk ), .D ( signal_24926 ), .Q ( signal_24927 ) ) ;
    buf_clk cell_10240 ( .C ( clk ), .D ( signal_24932 ), .Q ( signal_24933 ) ) ;
    buf_clk cell_10246 ( .C ( clk ), .D ( signal_24938 ), .Q ( signal_24939 ) ) ;
    buf_clk cell_10252 ( .C ( clk ), .D ( signal_24944 ), .Q ( signal_24945 ) ) ;
    buf_clk cell_10258 ( .C ( clk ), .D ( signal_24950 ), .Q ( signal_24951 ) ) ;
    buf_clk cell_10264 ( .C ( clk ), .D ( signal_24956 ), .Q ( signal_24957 ) ) ;
    buf_clk cell_10270 ( .C ( clk ), .D ( signal_24962 ), .Q ( signal_24963 ) ) ;
    buf_clk cell_10276 ( .C ( clk ), .D ( signal_24968 ), .Q ( signal_24969 ) ) ;
    buf_clk cell_10282 ( .C ( clk ), .D ( signal_24974 ), .Q ( signal_24975 ) ) ;
    buf_clk cell_10286 ( .C ( clk ), .D ( signal_24978 ), .Q ( signal_24979 ) ) ;
    buf_clk cell_10290 ( .C ( clk ), .D ( signal_24982 ), .Q ( signal_24983 ) ) ;
    buf_clk cell_10294 ( .C ( clk ), .D ( signal_24986 ), .Q ( signal_24987 ) ) ;
    buf_clk cell_10298 ( .C ( clk ), .D ( signal_24990 ), .Q ( signal_24991 ) ) ;
    buf_clk cell_10302 ( .C ( clk ), .D ( signal_24994 ), .Q ( signal_24995 ) ) ;
    buf_clk cell_10310 ( .C ( clk ), .D ( signal_25002 ), .Q ( signal_25003 ) ) ;
    buf_clk cell_10318 ( .C ( clk ), .D ( signal_25010 ), .Q ( signal_25011 ) ) ;
    buf_clk cell_10326 ( .C ( clk ), .D ( signal_25018 ), .Q ( signal_25019 ) ) ;
    buf_clk cell_10334 ( .C ( clk ), .D ( signal_25026 ), .Q ( signal_25027 ) ) ;
    buf_clk cell_10342 ( .C ( clk ), .D ( signal_25034 ), .Q ( signal_25035 ) ) ;
    buf_clk cell_10350 ( .C ( clk ), .D ( signal_25042 ), .Q ( signal_25043 ) ) ;
    buf_clk cell_10358 ( .C ( clk ), .D ( signal_25050 ), .Q ( signal_25051 ) ) ;
    buf_clk cell_10366 ( .C ( clk ), .D ( signal_25058 ), .Q ( signal_25059 ) ) ;
    buf_clk cell_10374 ( .C ( clk ), .D ( signal_25066 ), .Q ( signal_25067 ) ) ;
    buf_clk cell_10382 ( .C ( clk ), .D ( signal_25074 ), .Q ( signal_25075 ) ) ;
    buf_clk cell_10390 ( .C ( clk ), .D ( signal_25082 ), .Q ( signal_25083 ) ) ;
    buf_clk cell_10398 ( .C ( clk ), .D ( signal_25090 ), .Q ( signal_25091 ) ) ;
    buf_clk cell_10406 ( .C ( clk ), .D ( signal_25098 ), .Q ( signal_25099 ) ) ;
    buf_clk cell_10414 ( .C ( clk ), .D ( signal_25106 ), .Q ( signal_25107 ) ) ;
    buf_clk cell_10422 ( .C ( clk ), .D ( signal_25114 ), .Q ( signal_25115 ) ) ;
    buf_clk cell_10428 ( .C ( clk ), .D ( signal_25120 ), .Q ( signal_25121 ) ) ;
    buf_clk cell_10434 ( .C ( clk ), .D ( signal_25126 ), .Q ( signal_25127 ) ) ;
    buf_clk cell_10440 ( .C ( clk ), .D ( signal_25132 ), .Q ( signal_25133 ) ) ;
    buf_clk cell_10446 ( .C ( clk ), .D ( signal_25138 ), .Q ( signal_25139 ) ) ;
    buf_clk cell_10452 ( .C ( clk ), .D ( signal_25144 ), .Q ( signal_25145 ) ) ;

    /* cells in depth 33 */
    buf_clk cell_10229 ( .C ( clk ), .D ( signal_24921 ), .Q ( signal_24922 ) ) ;
    buf_clk cell_10235 ( .C ( clk ), .D ( signal_24927 ), .Q ( signal_24928 ) ) ;
    buf_clk cell_10241 ( .C ( clk ), .D ( signal_24933 ), .Q ( signal_24934 ) ) ;
    buf_clk cell_10247 ( .C ( clk ), .D ( signal_24939 ), .Q ( signal_24940 ) ) ;
    buf_clk cell_10253 ( .C ( clk ), .D ( signal_24945 ), .Q ( signal_24946 ) ) ;
    buf_clk cell_10259 ( .C ( clk ), .D ( signal_24951 ), .Q ( signal_24952 ) ) ;
    buf_clk cell_10265 ( .C ( clk ), .D ( signal_24957 ), .Q ( signal_24958 ) ) ;
    buf_clk cell_10271 ( .C ( clk ), .D ( signal_24963 ), .Q ( signal_24964 ) ) ;
    buf_clk cell_10277 ( .C ( clk ), .D ( signal_24969 ), .Q ( signal_24970 ) ) ;
    buf_clk cell_10283 ( .C ( clk ), .D ( signal_24975 ), .Q ( signal_24976 ) ) ;
    buf_clk cell_10287 ( .C ( clk ), .D ( signal_24979 ), .Q ( signal_24980 ) ) ;
    buf_clk cell_10291 ( .C ( clk ), .D ( signal_24983 ), .Q ( signal_24984 ) ) ;
    buf_clk cell_10295 ( .C ( clk ), .D ( signal_24987 ), .Q ( signal_24988 ) ) ;
    buf_clk cell_10299 ( .C ( clk ), .D ( signal_24991 ), .Q ( signal_24992 ) ) ;
    buf_clk cell_10303 ( .C ( clk ), .D ( signal_24995 ), .Q ( signal_24996 ) ) ;
    buf_clk cell_10311 ( .C ( clk ), .D ( signal_25003 ), .Q ( signal_25004 ) ) ;
    buf_clk cell_10319 ( .C ( clk ), .D ( signal_25011 ), .Q ( signal_25012 ) ) ;
    buf_clk cell_10327 ( .C ( clk ), .D ( signal_25019 ), .Q ( signal_25020 ) ) ;
    buf_clk cell_10335 ( .C ( clk ), .D ( signal_25027 ), .Q ( signal_25028 ) ) ;
    buf_clk cell_10343 ( .C ( clk ), .D ( signal_25035 ), .Q ( signal_25036 ) ) ;
    buf_clk cell_10351 ( .C ( clk ), .D ( signal_25043 ), .Q ( signal_25044 ) ) ;
    buf_clk cell_10359 ( .C ( clk ), .D ( signal_25051 ), .Q ( signal_25052 ) ) ;
    buf_clk cell_10367 ( .C ( clk ), .D ( signal_25059 ), .Q ( signal_25060 ) ) ;
    buf_clk cell_10375 ( .C ( clk ), .D ( signal_25067 ), .Q ( signal_25068 ) ) ;
    buf_clk cell_10383 ( .C ( clk ), .D ( signal_25075 ), .Q ( signal_25076 ) ) ;
    buf_clk cell_10391 ( .C ( clk ), .D ( signal_25083 ), .Q ( signal_25084 ) ) ;
    buf_clk cell_10399 ( .C ( clk ), .D ( signal_25091 ), .Q ( signal_25092 ) ) ;
    buf_clk cell_10407 ( .C ( clk ), .D ( signal_25099 ), .Q ( signal_25100 ) ) ;
    buf_clk cell_10415 ( .C ( clk ), .D ( signal_25107 ), .Q ( signal_25108 ) ) ;
    buf_clk cell_10423 ( .C ( clk ), .D ( signal_25115 ), .Q ( signal_25116 ) ) ;
    buf_clk cell_10429 ( .C ( clk ), .D ( signal_25121 ), .Q ( signal_25122 ) ) ;
    buf_clk cell_10435 ( .C ( clk ), .D ( signal_25127 ), .Q ( signal_25128 ) ) ;
    buf_clk cell_10441 ( .C ( clk ), .D ( signal_25133 ), .Q ( signal_25134 ) ) ;
    buf_clk cell_10447 ( .C ( clk ), .D ( signal_25139 ), .Q ( signal_25140 ) ) ;
    buf_clk cell_10453 ( .C ( clk ), .D ( signal_25145 ), .Q ( signal_25146 ) ) ;

    /* cells in depth 34 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_2383 ( .a ({signal_24917, signal_24903, signal_24889, signal_24875, signal_24861}), .b ({signal_8247, signal_8246, signal_8245, signal_8244, signal_2390}), .clk ( clk ), .r ({Fresh[8789], Fresh[8788], Fresh[8787], Fresh[8786], Fresh[8785], Fresh[8784], Fresh[8783], Fresh[8782], Fresh[8781], Fresh[8780]}), .c ({signal_8251, signal_8250, signal_8249, signal_8248, signal_2391}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_2384 ( .a ({signal_8251, signal_8250, signal_8249, signal_8248, signal_2391}), .b ({signal_8255, signal_8254, signal_8253, signal_8252, signal_27}) ) ;
    buf_clk cell_10230 ( .C ( clk ), .D ( signal_24922 ), .Q ( signal_24923 ) ) ;
    buf_clk cell_10236 ( .C ( clk ), .D ( signal_24928 ), .Q ( signal_24929 ) ) ;
    buf_clk cell_10242 ( .C ( clk ), .D ( signal_24934 ), .Q ( signal_24935 ) ) ;
    buf_clk cell_10248 ( .C ( clk ), .D ( signal_24940 ), .Q ( signal_24941 ) ) ;
    buf_clk cell_10254 ( .C ( clk ), .D ( signal_24946 ), .Q ( signal_24947 ) ) ;
    buf_clk cell_10260 ( .C ( clk ), .D ( signal_24952 ), .Q ( signal_24953 ) ) ;
    buf_clk cell_10266 ( .C ( clk ), .D ( signal_24958 ), .Q ( signal_24959 ) ) ;
    buf_clk cell_10272 ( .C ( clk ), .D ( signal_24964 ), .Q ( signal_24965 ) ) ;
    buf_clk cell_10278 ( .C ( clk ), .D ( signal_24970 ), .Q ( signal_24971 ) ) ;
    buf_clk cell_10284 ( .C ( clk ), .D ( signal_24976 ), .Q ( signal_24977 ) ) ;
    buf_clk cell_10288 ( .C ( clk ), .D ( signal_24980 ), .Q ( signal_24981 ) ) ;
    buf_clk cell_10292 ( .C ( clk ), .D ( signal_24984 ), .Q ( signal_24985 ) ) ;
    buf_clk cell_10296 ( .C ( clk ), .D ( signal_24988 ), .Q ( signal_24989 ) ) ;
    buf_clk cell_10300 ( .C ( clk ), .D ( signal_24992 ), .Q ( signal_24993 ) ) ;
    buf_clk cell_10304 ( .C ( clk ), .D ( signal_24996 ), .Q ( signal_24997 ) ) ;
    buf_clk cell_10312 ( .C ( clk ), .D ( signal_25004 ), .Q ( signal_25005 ) ) ;
    buf_clk cell_10320 ( .C ( clk ), .D ( signal_25012 ), .Q ( signal_25013 ) ) ;
    buf_clk cell_10328 ( .C ( clk ), .D ( signal_25020 ), .Q ( signal_25021 ) ) ;
    buf_clk cell_10336 ( .C ( clk ), .D ( signal_25028 ), .Q ( signal_25029 ) ) ;
    buf_clk cell_10344 ( .C ( clk ), .D ( signal_25036 ), .Q ( signal_25037 ) ) ;
    buf_clk cell_10352 ( .C ( clk ), .D ( signal_25044 ), .Q ( signal_25045 ) ) ;
    buf_clk cell_10360 ( .C ( clk ), .D ( signal_25052 ), .Q ( signal_25053 ) ) ;
    buf_clk cell_10368 ( .C ( clk ), .D ( signal_25060 ), .Q ( signal_25061 ) ) ;
    buf_clk cell_10376 ( .C ( clk ), .D ( signal_25068 ), .Q ( signal_25069 ) ) ;
    buf_clk cell_10384 ( .C ( clk ), .D ( signal_25076 ), .Q ( signal_25077 ) ) ;
    buf_clk cell_10392 ( .C ( clk ), .D ( signal_25084 ), .Q ( signal_25085 ) ) ;
    buf_clk cell_10400 ( .C ( clk ), .D ( signal_25092 ), .Q ( signal_25093 ) ) ;
    buf_clk cell_10408 ( .C ( clk ), .D ( signal_25100 ), .Q ( signal_25101 ) ) ;
    buf_clk cell_10416 ( .C ( clk ), .D ( signal_25108 ), .Q ( signal_25109 ) ) ;
    buf_clk cell_10424 ( .C ( clk ), .D ( signal_25116 ), .Q ( signal_25117 ) ) ;
    buf_clk cell_10430 ( .C ( clk ), .D ( signal_25122 ), .Q ( signal_25123 ) ) ;
    buf_clk cell_10436 ( .C ( clk ), .D ( signal_25128 ), .Q ( signal_25129 ) ) ;
    buf_clk cell_10442 ( .C ( clk ), .D ( signal_25134 ), .Q ( signal_25135 ) ) ;
    buf_clk cell_10448 ( .C ( clk ), .D ( signal_25140 ), .Q ( signal_25141 ) ) ;
    buf_clk cell_10454 ( .C ( clk ), .D ( signal_25146 ), .Q ( signal_25147 ) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_24947, signal_24941, signal_24935, signal_24929, signal_24923}), .Q ({SO_s4[7], SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_24977, signal_24971, signal_24965, signal_24959, signal_24953}), .Q ({SO_s4[6], SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_24997, signal_24993, signal_24989, signal_24985, signal_24981}), .Q ({SO_s4[5], SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_25037, signal_25029, signal_25021, signal_25013, signal_25005}), .Q ({SO_s4[4], SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_8255, signal_8254, signal_8253, signal_8252, signal_27}), .Q ({SO_s4[3], SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_25077, signal_25069, signal_25061, signal_25053, signal_25045}), .Q ({SO_s4[2], SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_25117, signal_25109, signal_25101, signal_25093, signal_25085}), .Q ({SO_s4[1], SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_25147, signal_25141, signal_25135, signal_25129, signal_25123}), .Q ({SO_s4[0], SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
