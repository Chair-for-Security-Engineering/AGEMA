module AES_Top(x, y);
 input [257:0] x;
 output [128:0] y;

 wire [1963:0] t;
  FX FX_inst(.x({t[668], t[667], t[666], t[665], t[664], t[663], t[662], t[661], t[660], t[659], t[658], t[657], t[656], t[655], t[654], t[653], t[652], t[651], t[650], t[649], t[648], t[647], t[646], t[645], t[644], t[643], t[642], t[641], t[640], t[639], t[638], t[637], t[636], t[635], t[634], t[633], t[632], t[631], t[630], t[629], t[628], t[627], t[626], t[625], t[624], t[623], t[622], t[621], t[620], t[619], t[618], t[617], t[616], t[615], t[614], t[613], t[612], t[611], t[610], t[609], t[608], t[607], t[606], t[605], t[604], t[603], t[602], t[601], t[600], t[599], t[598], t[597], t[596], t[595], t[594], t[593], t[592], t[591], t[590], t[589], t[588], t[587], t[586], t[585], t[584], t[583], t[582], t[581], t[580], t[579], t[578], t[577], t[576], t[575], t[574], t[573], t[572], t[571], t[570], t[569], t[568], t[567], t[566], t[565], t[564], t[563], t[562], t[561], t[560], t[559], t[558], t[557], t[556], t[555], t[554], t[553], t[552], t[551], t[550], t[549], t[548], t[547], t[546], t[545], t[544], t[543], t[542], t[541], t[540], t[539], t[538], t[537], t[536], t[535], t[534], t[533], t[532], t[531], t[530], t[529], t[528], t[527], t[526], t[525], t[524], t[523], t[522], t[521], t[520], t[519], t[518], t[517], t[516], t[515], t[514], t[513], t[512], t[511], t[510], t[509], t[508], t[507], t[506], t[505], t[504], t[503], t[502], t[501], t[500], t[499], t[498], t[497], t[496], t[495], t[494], t[493], t[492], t[491], t[490], t[489], t[488], t[487], t[486], t[485], t[484], t[483], t[482], t[481], t[480], t[479], t[478], t[477], t[476], t[475], t[474], t[473], t[472], t[471], t[470], t[469], t[468], t[467], t[466], t[465], t[464], t[463], t[462], t[461], t[460], t[459], t[458], t[457], t[456], t[455], t[454], t[453], t[452], t[451], t[450], t[449], t[448], t[447], t[446], t[445], t[444], t[443], t[442], t[441], t[440], t[439], t[438], t[437], t[436], t[435], t[434], t[433], t[432], t[431], t[430], t[429], t[428], t[427], t[426], t[425], t[424], t[423], t[422], t[421], t[420], t[419], t[418], t[417], t[416], t[415], t[414], t[413], t[412], t[411], t[410], t[409], t[408], t[407], t[406], t[405], t[404], t[403], t[402], t[401], t[400], t[399], t[398], t[397], t[396], t[395], t[394], t[393], t[392], t[391], t[390], t[389], t[388], t[387], t[386], t[385], t[384], t[383], t[382], t[381], t[380], t[379], t[378], t[377], t[376], t[375], t[374], t[373], t[372], t[371], t[370], t[369], t[368], t[367], t[366], t[365], t[364], t[363], t[362], t[361], t[360], t[359], t[358], t[357], t[356], t[355], t[354], t[353], t[352], t[351], t[350], t[349], t[348], t[347], t[346], t[345], t[344], t[343], t[342], t[341], t[340], t[339], t[338], t[337], t[336], t[335], t[334], t[333], t[332], t[331], t[330], t[329], t[328], t[327], t[326], t[325], t[324], t[323], t[322], t[321], t[320], t[319], t[318], t[317], t[316], t[315], t[314], t[313], t[312], t[311], t[310], t[309], t[308], t[307], t[306], t[305], t[304], t[303], t[302], t[301], t[300], t[299], t[298], t[297], t[296], t[295], t[294], t[293], t[292], t[291], t[290], t[289], t[288], t[287], t[286], t[285], t[284], t[283], t[282], t[281], t[280], t[279], t[278], t[277], t[276], t[275], t[274], t[273], t[272], t[271], t[270], t[269], t[268], t[267], t[266], t[265], t[264], t[263], t[262], t[261], t[260], t[259], t[258], t[257], t[256], t[255], t[254], t[253], t[252], t[251], t[250], t[249], t[248], t[247], t[246], t[245], t[244], t[243], t[242], t[241], t[240], t[239], t[238], t[237], t[236], t[235], t[234], t[233], t[232], t[231], t[230], t[229], t[228], t[227], t[226], t[225], t[224], t[223], t[222], t[221], t[220], t[219], t[218], t[217], t[216], t[215], t[214], t[213], t[212], t[211], t[210], t[209], t[208], t[207], t[206], t[205], t[204], t[203], t[202], t[201], t[200], t[199], t[198], t[197], t[196], t[195], t[194], t[193], t[192], t[191], t[190], t[189], t[188], t[187], t[186], t[185], t[184], t[183], t[182], t[181], t[180], t[179], t[178], t[177], t[176], t[175], t[174], t[173], t[172], t[171], t[170], t[169], t[168], t[167], t[166], t[165], t[164], t[163], t[162], t[161], t[160], t[159], t[158], t[157], t[156], t[155], t[154], t[153], t[152], t[151], t[150], t[149], t[148], t[147], t[146], t[145], t[144], t[143], t[142], t[141], t[140], t[139], t[138], t[137], t[136], t[135], t[134], t[133], t[132], t[131], t[130], t[129], t[128], t[127], t[126], t[125], t[124], t[123], t[122], t[121], t[120], t[119], t[118], t[117], t[116], t[115], t[114], t[113], t[112], t[111], t[110], t[109], t[108], t[107], t[106], t[105], t[104], t[103], t[102], t[101], t[100], t[99], t[98], t[97], t[96], t[95], t[94], t[93], t[92], t[91], t[90], t[89], t[88], t[87], t[86], t[85], t[84], t[83], t[82], t[81], t[80], t[79], t[78], t[77], t[76], t[75], t[74], t[73], t[72], t[71], t[70], t[69], t[68], t[67], t[66], t[65], t[64], t[63], t[62], t[61], t[60], t[59], t[58], t[57], t[56], t[55], t[54], t[53], t[52], t[51], t[50], t[49], t[48], t[47], t[46], t[45], t[44], t[43], t[42], t[41], t[40], t[39], t[38], t[37], t[36], t[35], t[34], t[33], t[32], t[31], t[30], t[29], t[28], t[27], t[26], t[25], t[24], t[23], t[22], t[21], t[20], t[19], t[18], t[17], t[16], t[15], t[14], t[13], t[12], t[11], t[10], t[9], t[8], t[7], t[6], t[5], t[4], t[3], t[2], t[1], t[0]}), .y({t[1046], t[1045], t[1044], t[1043], t[1042], t[1041], t[1040], t[1039], t[1038], t[1037], t[1036], t[1035], t[1034], t[1033], t[1032], t[1031], t[1030], t[1029], t[1028], t[1027], t[1026], t[1025], t[1024], t[1023], t[1022], t[1021], t[1020], t[1019], t[1018], t[1017], t[1016], t[1015], t[1014], t[1013], t[1012], t[1011], t[1010], t[1009], t[1008], t[1007], t[1006], t[1005], t[1004], t[1003], t[1002], t[1001], t[1000], t[999], t[998], t[997], t[996], t[995], t[994], t[993], t[992], t[991], t[990], t[989], t[988], t[987], t[986], t[985], t[984], t[983], t[982], t[981], t[980], t[979], t[978], t[977], t[976], t[975], t[974], t[973], t[972], t[971], t[970], t[969], t[968], t[967], t[966], t[965], t[964], t[963], t[962], t[961], t[960], t[959], t[958], t[957], t[956], t[955], t[954], t[953], t[952], t[951], t[950], t[949], t[948], t[947], t[946], t[945], t[944], t[943], t[942], t[941], t[940], t[939], t[938], t[937], t[936], t[935], t[934], t[933], t[932], t[931], t[930], t[929], t[928], t[927], t[926], t[925], t[924], t[923], t[922], t[921], t[920], t[919], t[918], t[917], t[916], t[915], t[914], t[913], t[912], t[911], t[910], t[909], t[908], t[907], t[906], t[905], t[904], t[903], t[902], t[901], t[900], t[899], t[898], t[897], t[896], t[895], t[894], t[893], t[892], t[891], t[890], t[889], t[888], t[887], t[886], t[885], t[884], t[883], t[882], t[881], t[880], t[879], t[878], t[877], t[876], t[875], t[874], t[873], t[872], t[871], t[870], t[869], t[868], t[867], t[866], t[865], t[864], t[863], t[862], t[861], t[860], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[852], t[851], t[850], t[849], t[848], t[847], t[846], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[803], t[802], t[801], t[800], t[799], t[798], t[797], t[796], t[795], t[794], t[793], t[792], t[791], t[790], t[789], t[788], t[787], t[786], t[785], t[784], t[783], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[761], t[760], t[759], t[758], t[757], t[756], t[755], t[754], t[753], t[752], t[751], t[750], t[749], t[748], t[747], t[746], t[745], t[744], t[743], t[742], t[741], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[719], t[718], t[717], t[716], t[715], t[714], t[713], t[712], t[711], t[710], t[709], t[708], t[707], t[706], t[705], t[704], t[703], t[702], t[701], t[700], t[699], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[684], t[683], t[682], t[681], t[680], t[679], t[678], t[677], t[676], t[675], t[674], t[673], t[672], t[671], t[670], t[669]}));
  R1_ind R1_ind_inst(.x({t[644], t[1034], t[633], t[1031], t[643], t[1035], t[634], t[1030], t[636], t[1028], t[645], t[1033], t[635], t[1029], t[1027], t[642], t[1036], t[1032], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[167], t[129], t[751], x[166], t[130], t[750], x[165], t[131], t[749], x[164], t[132], t[748], t[747], x[163], t[138], t[756], x[162], t[139], t[755], x[161], t[140], t[754], x[160], t[141], t[753], t[752], x[175], t[147], t[761], x[174], t[148], t[760], x[173], t[149], t[759], x[172], t[150], t[758], t[757], x[171], t[156], t[766], x[170], t[157], t[765], x[169], t[158], t[764], x[168], t[159], t[763], t[762], x[183], t[165], t[771], x[182], t[166], t[770], x[181], t[167], t[769], x[180], t[168], t[768], t[767], x[179], t[174], t[776], x[178], t[175], t[775], x[177], t[176], t[774], x[176], t[177], t[773], t[772], x[191], t[183], t[781], x[190], t[184], t[780], x[189], t[185], t[779], x[188], t[186], t[778], t[777], x[187], t[192], t[786], x[186], t[193], t[785], x[185], t[194], t[784], x[184], t[195], t[783], t[782], x[199], t[201], t[791], x[198], t[202], t[790], x[197], t[203], t[789], x[196], t[204], t[788], t[787], x[195], t[210], t[796], x[194], t[211], t[795], x[193], t[212], t[794], x[192], t[213], t[793], t[792], x[207], t[219], t[801], x[206], t[220], t[800], x[205], t[221], t[799], x[204], t[222], t[798], t[797], x[203], t[228], t[806], x[202], t[229], t[805], x[201], t[230], t[804], x[200], t[231], t[803], t[802], x[215], t[237], t[811], x[214], t[238], t[810], x[213], t[239], t[809], x[212], t[240], t[808], t[807], x[211], t[246], t[816], x[210], t[247], t[815], x[209], t[248], t[814], x[208], t[249], t[813], t[812], x[223], t[255], t[821], x[222], t[256], t[820], x[221], t[257], t[819], x[220], t[258], t[818], t[817], x[219], t[264], t[826], x[218], t[265], t[825], x[217], t[266], t[824], x[216], t[267], t[823], t[822], t[651], t[1041], x[231], t[273], t[831], t[652], t[1040], x[230], t[274], t[830], t[653], t[1039], x[229], t[275], t[829], t[654], t[1038], t[1037], x[228], t[276], t[828], t[827], t[660], t[1046], x[227], t[282], t[836], t[661], t[1045], x[226], t[283], t[835], t[662], t[1044], x[225], t[284], t[834], t[6], t[674], t[673], t[663], t[1043], t[1042], x[224], t[285], t[833], t[832], x[239], t[75], t[721], t[291], t[841], x[238], t[76], t[720], t[292], t[840], x[237], t[77], t[719], t[293], t[839], x[236], t[78], t[718], t[717], t[294], t[838], t[837], x[235], t[84], t[726], t[300], t[846], x[234], t[85], t[725], t[301], t[845], x[233], t[86], t[724], t[302], t[844], x[232], t[87], t[723], t[722], t[303], t[843], t[842], x[247], t[93], t[731], t[309], t[851], x[246], t[94], t[730], t[310], t[850], x[245], t[95], t[729], t[311], t[849], x[244], t[96], t[728], t[727], t[312], t[848], t[847], x[243], t[102], t[736], t[318], t[856], x[242], t[103], t[735], t[319], t[855], x[241], t[104], t[734], t[320], t[854], x[240], t[105], t[733], t[732], t[321], t[853], t[852], t[57], t[711], x[255], t[111], t[741], t[327], t[861], t[58], t[710], x[254], t[112], t[740], t[328], t[860], t[59], t[709], x[253], t[113], t[739], t[329], t[859], t[60], t[708], t[707], x[252], t[114], t[738], t[737], t[330], t[858], t[857], t[66], t[716], x[251], t[120], t[746], t[336], t[866], t[67], t[715], x[250], t[121], t[745], t[337], t[865], t[68], t[714], x[249], t[122], t[744], t[338], t[864], t[9], t[676], t[675], t[69], t[713], t[712], x[248], t[123], t[743], t[742], t[339], t[863], t[862], t[33], t[692], t[691], t[24], t[686], t[685], t[12], t[678], t[677], t[15], t[680], t[679], x[257], t[54], t[706], t[705], t[48], t[702], t[701], t[51], t[704], t[703], t[42], t[698], t[697], t[39], t[696], t[695], t[45], t[700], t[699], t[36], t[694], t[693], t[27], t[688], t[687], t[21], t[684], t[683], t[18], t[682], t[681], t[30], t[690], t[689], t[3], t[672], t[671], t[627], t[1023], t[626], t[1024], t[625], t[1025], t[624], t[1026], t[1022], t[618], t[1018], t[617], t[1019], t[616], t[1020], t[615], t[1021], t[1017], t[609], t[1013], t[608], t[1014], t[607], t[1015], t[606], t[1016], t[1012], t[600], t[1008], t[599], t[1009], t[598], t[1010], t[597], t[1011], t[1007], t[591], t[1003], t[590], t[1004], t[589], t[1005], t[588], t[1006], t[1002], t[582], t[998], t[581], t[999], t[580], t[1000], t[579], t[1001], t[997], t[573], t[993], t[572], t[994], t[571], t[995], t[570], t[996], t[992], t[564], t[988], t[563], t[989], t[562], t[990], t[561], t[991], t[987], t[555], t[983], t[554], t[984], t[553], t[985], t[552], t[986], t[982], t[546], t[978], t[545], t[979], t[544], t[980], t[543], t[981], t[977], t[537], t[973], t[536], t[974], t[535], t[975], t[534], t[976], t[972], t[528], t[968], t[527], t[969], t[526], t[970], t[525], t[971], t[967], t[519], t[963], t[518], t[964], t[517], t[965], t[516], t[966], t[962], t[510], t[958], t[509], t[959], t[508], t[960], t[507], t[961], t[957], t[501], t[953], t[500], t[954], t[499], t[955], t[498], t[956], t[952], t[492], t[948], t[491], t[949], t[490], t[950], t[489], t[951], t[947], t[483], t[943], t[482], t[944], t[481], t[945], t[480], t[946], t[942], t[474], t[938], t[473], t[939], t[472], t[940], t[471], t[941], t[937], t[465], t[933], t[464], t[934], t[463], t[935], t[462], t[936], t[932], t[456], t[928], t[455], t[929], t[454], t[930], t[453], t[931], t[927], t[447], t[923], t[446], t[924], t[445], t[925], t[444], t[926], t[922], t[438], t[918], t[437], t[919], t[436], t[920], t[435], t[921], t[917], t[429], t[913], t[428], t[914], t[427], t[915], t[426], t[916], t[912], t[420], t[908], t[419], t[909], t[418], t[910], t[417], t[911], t[907], t[411], t[903], t[410], t[904], t[409], t[905], t[408], t[906], t[902], t[402], t[898], t[401], t[899], t[400], t[900], t[399], t[901], t[897], t[393], t[893], t[392], t[894], t[391], t[895], t[390], t[896], t[892], t[384], t[888], t[383], t[889], t[382], t[890], t[381], t[891], t[887], t[375], t[883], t[374], t[884], t[373], t[885], t[372], t[886], t[882], t[366], t[878], t[365], t[879], t[364], t[880], t[363], t[881], t[877], t[357], t[873], t[356], t[874], t[355], t[875], t[354], t[876], t[872], t[348], t[868], t[347], t[869], t[346], t[870], t[345], t[871], t[867], t[0], t[670], t[669]}), .y({t[1466], t[1465], t[1464], t[1463], t[1462], t[1461], t[1460], t[1459], t[1458], t[1457], t[1456], t[1455], t[1454], t[1453], t[1452], t[1451], t[1450], t[1449], t[1448], t[1447], t[1446], t[1445], t[1444], t[1443], t[1442], t[1441], t[1440], t[1439], t[1438], t[1437], t[1436], t[1435], t[1434], t[1433], t[1432], t[1431], t[1430], t[1429], t[1428], t[1427], t[1426], t[1425], t[1424], t[1423], t[1422], t[1421], t[1420], t[1419], t[1418], t[1417], t[1416], t[1415], t[1414], t[1413], t[1412], t[1411], t[1410], t[1409], t[1408], t[1407], t[1406], t[1405], t[1404], t[1403], t[1402], t[1401], t[1400], t[1399], t[1398], t[1397], t[1396], t[1395], t[1394], t[1393], t[1392], t[1391], t[1390], t[1389], t[1388], t[1387], t[1386], t[1385], t[1384], t[1383], t[1382], t[1381], t[1380], t[1379], t[1378], t[1377], t[1376], t[1375], t[1374], t[1373], t[1372], t[1371], t[1370], t[1369], t[1368], t[1367], t[1366], t[1365], t[1364], t[1363], t[1362], t[1361], t[1360], t[1359], t[1358], t[1357], t[1356], t[1355], t[1354], t[1353], t[1352], t[1351], t[1350], t[1349], t[1348], t[1347], t[1346], t[1345], t[1344], t[1343], t[1342], t[1341], t[1340], t[1339], t[1338], t[1337], t[1336], t[1335], t[1334], t[1333], t[1332], t[1331], t[1330], t[1329], t[1328], t[1327], t[1326], t[1325], t[1324], t[1323], t[1322], t[1321], t[1320], t[1319], t[1318], t[1317], t[1316], t[1315], t[1314], t[1313], t[1312], t[1311], t[1310], t[1309], t[1308], t[1307], t[1306], t[1305], t[1304], t[1303], t[1302], t[1301], t[1300], t[1299], t[1298], t[1297], t[1296], t[1295], t[1294], t[1293], t[1292], t[1291], t[1290], t[1289], t[1288], t[1287], t[1286], t[1285], t[1284], t[1283], t[1282], t[1281], t[1280], t[1279], t[1278], t[1277], t[1276], t[1275], t[1274], t[1273], t[1272], t[1271], t[1270], t[1269], t[1268], t[1267], t[1266], t[1265], t[1264], t[1263], t[1262], t[1261], t[1260], t[1259], t[1258], t[1257], t[1256], t[1255], t[1254], t[1253], t[1252], t[1251], t[1250], t[1249], t[1248], t[1247], t[1246], t[1245], t[1244], t[1243], t[1242], t[1241], t[1240], t[1239], t[1238], t[1237], t[1236], t[1235], t[1234], t[1233], t[1232], t[1231], t[1230], t[1229], t[1228], t[1227], t[1226], t[1225], t[1224], t[1223], t[1222], t[1221], t[1220], t[1219], t[1218], t[1217], t[1216], t[1215], t[1214], t[1213], t[1212], t[1211], t[1210], t[1209], t[1208], t[1207], t[1206], t[1205], t[1204], t[1203], t[1202], t[1201], t[1200], t[1199], t[1198], t[1197], t[1196], t[1195], t[1194], t[1193], t[1192], t[1191], t[1190], t[1189], t[1188], t[1187], t[1186], t[1185], t[1184], t[1183], t[1182], t[1181], t[1180], t[1179], t[1178], t[1177], t[1176], t[1175], t[1174], t[1173], t[1172], t[1171], t[1170], t[1169], t[1168], t[1167], t[1166], t[1165], t[1164], t[1163], t[1162], t[1161], t[1160], t[1159], t[1158], t[1157], t[1156], t[1155], t[1154], t[1153], t[1152], t[1151], t[1150], t[1149], t[1148], t[1147], t[1146], t[1145], t[1144], t[1143], t[1142], t[1141], t[1140], t[1139], t[1138], t[1137], t[1136], t[1135], t[1134], t[1133], t[1132], t[1131], t[1130], t[1129], t[1128], t[1127], t[1126], t[1125], t[1124], t[1123], t[1122], t[1121], t[1120], t[1119], t[1118], t[1117], t[1116], t[1115], t[1114], t[1113], t[1112], t[1111], t[1110], t[1109], t[1108], t[1107], t[1106], t[1105], t[1104], t[1103], t[1102], t[1101], t[1100], t[1099], t[1098], t[1097], t[1096], t[1095], t[1094], t[1093], t[1092], t[1091], t[1090], t[1089], t[1088], t[1087], t[1086], t[1085], t[1084], t[1083], t[1082], t[1081], t[1080], t[1079], t[1078], t[1077], t[1076], t[1075], t[1074], t[1073], t[1072], t[1071], t[1070], t[1069], t[1068], t[1067], t[1066], t[1065], t[1064], t[1063], t[1062], t[1061], t[1060], t[1059], t[1058], t[1057], t[1056], t[1055], t[1054], t[1053], t[1052], t[1051], t[1050], t[1049], t[1048], t[1047]}));
  R2_ind R2_ind_inst(.x({t[648], t[649], t[638], t[640], t[647], t[641], t[639], t[637], t[636], t[635], t[634], t[633], t[650], t[646], t[645], t[644], t[643], t[642], x[120], x[121], x[122], x[123], x[124], x[125], x[126], x[127], x[112], x[113], x[114], x[115], x[116], x[117], x[118], x[119], t[611], x[104], t[612], x[105], t[613], x[106], t[614], t[610], t[609], t[608], t[607], t[606], x[107], t[602], x[108], t[603], x[109], t[604], x[110], t[605], t[601], t[600], t[599], t[598], t[597], x[111], t[593], x[96], t[629], t[594], x[97], t[630], t[595], x[98], t[631], t[596], t[592], t[591], t[590], t[589], t[588], x[99], t[632], t[628], t[627], t[626], t[625], t[624], t[584], x[100], t[620], t[585], x[101], t[621], t[586], x[102], t[622], t[587], t[583], t[582], t[581], t[580], t[579], x[103], t[623], t[619], t[618], t[617], t[616], t[615], x[88], x[89], x[90], x[91], x[92], x[93], x[94], x[95], x[80], x[81], x[82], x[83], x[84], x[85], x[86], x[87], x[72], t[557], x[73], t[558], x[74], t[559], x[75], t[560], t[556], t[555], t[554], t[553], t[552], x[76], t[548], x[77], t[549], x[78], t[550], x[79], t[551], t[547], t[546], t[545], t[544], t[543], t[521], x[64], t[539], t[522], x[65], t[540], t[523], x[66], t[541], t[524], t[520], t[519], t[518], t[517], t[516], x[67], t[542], t[538], t[537], t[536], t[535], t[534], t[512], x[68], t[530], t[513], x[69], t[531], t[514], x[70], t[532], t[515], t[511], t[510], t[509], t[508], t[507], x[71], t[533], t[529], t[528], t[527], t[526], t[525], x[56], x[57], x[58], x[59], x[60], x[61], x[62], x[63], x[48], t[485], x[49], t[486], x[50], t[487], x[51], t[488], t[484], t[483], t[482], t[481], t[480], x[52], t[476], x[53], t[477], x[54], t[478], x[55], t[479], t[475], t[474], t[473], t[472], t[471], x[40], t[467], x[41], t[468], x[42], t[469], x[43], t[470], t[466], t[465], t[464], t[463], t[462], x[44], t[458], x[45], t[459], x[46], t[460], x[47], t[461], t[457], t[456], t[455], t[454], t[453], x[32], t[449], x[33], t[450], x[34], t[451], x[35], t[452], t[448], t[447], t[446], t[445], t[444], x[36], t[440], x[37], t[441], x[38], t[442], x[39], t[443], t[439], t[438], t[437], t[436], t[435], t[575], t[503], x[24], t[576], t[504], t[432], x[25], t[577], t[505], t[433], x[26], t[578], t[574], t[573], t[572], t[571], t[570], t[506], t[502], t[501], t[500], t[499], t[498], t[434], x[27], t[566], t[494], t[422], x[28], t[567], t[495], t[423], x[29], t[496], t[568], t[424], x[30], t[431], t[430], t[429], t[428], t[427], t[426], t[497], t[493], t[492], t[491], t[490], t[489], t[569], t[565], t[564], t[563], t[562], t[561], t[425], t[421], t[420], t[419], t[418], t[417], x[31], t[413], x[16], t[414], x[17], t[415], x[18], t[416], t[412], t[411], t[410], t[409], t[408], x[19], t[404], x[20], t[405], x[21], t[406], x[22], t[407], t[403], t[402], t[401], t[400], t[399], x[23], t[395], x[8], t[396], x[9], t[397], x[10], t[398], t[394], t[393], t[392], t[391], t[390], x[11], t[386], x[12], t[387], x[13], t[388], x[14], t[389], t[385], t[384], t[383], t[382], t[381], x[15], t[377], x[0], t[359], t[378], x[1], t[360], t[379], x[2], t[361], t[380], t[376], t[375], t[374], t[373], t[372], x[3], t[362], t[358], t[357], t[356], t[355], t[354], t[368], x[4], t[350], t[369], x[5], t[351], t[370], x[6], t[352], t[371], t[367], t[366], t[365], t[364], t[363], x[7], t[353], t[349], t[348], t[347], t[346], t[345], x[248], x[249], x[250], x[251], x[252], x[253], x[254], x[255], x[240], x[241], x[242], x[243], x[244], x[245], x[246], x[247], x[232], x[233], x[234], x[235], x[236], x[237], x[238], x[239], t[665], x[224], t[666], x[225], t[667], x[226], t[668], t[664], t[663], t[662], t[661], t[660], x[227], t[656], x[228], t[657], x[229], t[658], x[230], t[8], t[7], t[6], t[659], t[655], t[654], t[653], t[652], t[651], x[231], x[216], t[341], x[217], t[342], x[218], t[343], x[219], t[344], t[340], t[339], t[338], t[337], t[336], x[220], t[332], x[221], t[333], x[222], t[334], x[223], t[335], t[331], t[330], t[329], t[328], t[327], x[208], t[323], x[209], t[324], x[210], t[325], x[211], t[326], t[322], t[321], t[320], t[319], t[318], x[212], t[314], x[213], t[315], x[214], t[316], x[215], t[317], t[313], t[312], t[311], t[310], t[309], x[200], t[305], x[201], t[306], x[202], t[307], x[203], t[308], t[304], t[303], t[302], t[301], t[300], x[204], t[296], x[205], t[297], x[206], t[298], x[207], t[299], t[295], t[294], t[293], t[292], t[291], x[192], t[287], x[193], t[288], x[194], t[289], x[195], t[290], t[286], t[285], t[284], t[283], t[282], x[196], t[278], x[197], t[279], x[198], t[280], x[199], t[281], t[277], t[276], t[275], t[274], t[273], x[184], t[269], x[185], t[270], x[186], t[271], x[187], t[272], t[268], t[267], t[266], t[265], t[264], x[188], t[260], x[189], t[261], x[190], t[262], x[191], t[263], t[259], t[258], t[257], t[256], t[255], x[176], t[251], x[177], t[252], x[178], t[253], x[179], t[254], t[250], t[249], t[248], t[247], t[246], x[180], t[242], x[181], t[243], x[182], t[244], x[183], t[245], t[241], t[240], t[239], t[238], t[237], x[168], t[233], x[169], t[234], x[170], t[235], x[171], t[236], t[232], t[231], t[230], t[229], t[228], x[172], t[224], x[173], t[225], x[174], t[226], x[175], t[227], t[223], t[222], t[221], t[220], t[219], x[160], t[215], x[161], t[216], x[162], t[217], x[163], t[218], t[214], t[213], t[212], t[211], t[210], x[164], t[206], x[165], t[207], x[166], t[208], x[167], t[209], t[205], t[204], t[203], t[202], t[201], x[152], t[197], x[153], t[198], x[154], t[199], x[155], t[200], t[196], t[195], t[194], t[193], t[192], x[156], t[188], x[157], t[189], x[158], t[190], x[159], t[191], t[187], t[186], t[185], t[184], t[183], t[125], x[144], t[179], t[126], x[145], t[180], t[127], x[146], t[181], t[128], t[124], t[123], t[122], t[121], t[120], x[147], t[182], t[178], t[177], t[176], t[175], t[174], t[116], x[148], t[170], t[117], x[149], t[171], t[118], x[150], t[172], t[119], t[115], t[114], t[113], t[112], t[111], x[151], t[173], t[169], t[168], t[167], t[166], t[165], t[107], x[136], t[161], t[108], x[137], t[162], t[109], x[138], t[163], t[110], t[106], t[105], t[104], t[103], t[102], x[139], t[164], t[160], t[159], t[158], t[157], t[156], t[98], x[140], t[152], t[99], x[141], t[153], t[100], x[142], t[154], t[101], t[97], t[96], t[95], t[94], t[93], x[143], t[155], t[151], t[150], t[149], t[148], t[147], t[89], x[128], t[143], t[71], t[90], x[129], t[144], t[72], t[91], x[130], t[145], t[73], t[92], t[88], t[87], t[86], t[85], t[84], x[131], t[146], t[142], t[141], t[140], t[139], t[138], t[74], t[70], t[69], t[68], t[67], t[66], t[80], x[132], t[134], t[62], t[81], x[133], t[135], t[63], t[82], x[134], t[136], t[64], t[83], t[79], t[78], t[77], t[76], t[75], x[135], t[137], t[133], t[132], t[131], t[130], t[129], t[65], t[61], t[60], t[59], t[58], t[57], t[35], t[34], t[33], t[26], t[25], t[24], t[14], t[13], t[12], t[17], t[16], t[15], t[11], t[10], t[9], x[257], t[56], t[55], t[54], t[50], t[49], t[48], t[53], t[52], t[51], t[44], t[43], t[42], t[41], t[40], t[39], t[47], t[46], t[45], t[38], t[37], t[36], t[29], t[28], t[27], t[23], t[22], t[21], t[20], t[19], t[18], t[32], t[31], t[30], t[5], t[4], t[3], t[1], t[2], t[1469], t[1468], t[1467], t[0]}), .y({t[1909], t[1908], t[1907], t[1906], t[1905], t[1904], t[1903], t[1902], t[1901], t[1900], t[1899], t[1898], t[1897], t[1896], t[1895], t[1894], t[1893], t[1892], t[1891], t[1890], t[1889], t[1888], t[1887], t[1886], t[1885], t[1884], t[1883], t[1882], t[1881], t[1880], t[1879], t[1878], t[1877], t[1876], t[1875], t[1874], t[1873], t[1872], t[1871], t[1870], t[1869], t[1868], t[1867], t[1866], t[1865], t[1864], t[1863], t[1862], t[1861], t[1860], t[1859], t[1858], t[1857], t[1856], t[1855], t[1854], t[1853], t[1852], t[1851], t[1850], t[1849], t[1848], t[1847], t[1846], t[1845], t[1844], t[1843], t[1842], t[1841], t[1840], t[1839], t[1838], t[1837], t[1836], t[1835], t[1834], t[1833], t[1832], t[1831], t[1830], t[1829], t[1828], t[1827], t[1826], t[1825], t[1824], t[1823], t[1822], t[1821], t[1820], t[1819], t[1818], t[1817], t[1816], t[1815], t[1814], t[1813], t[1812], t[1811], t[1810], t[1809], t[1808], t[1807], t[1806], t[1805], t[1804], t[1803], t[1802], t[1801], t[1800], t[1799], t[1798], t[1797], t[1796], t[1795], t[1794], t[1793], t[1792], t[1791], t[1790], t[1789], t[1788], t[1787], t[1786], t[1785], t[1784], t[1783], t[1782], t[1781], t[1780], t[1779], t[1778], t[1777], t[1776], t[1775], t[1774], t[1773], t[1772], t[1771], t[1770], t[1769], t[1768], t[1767], t[1766], t[1765], t[1764], t[1763], t[1762], t[1761], t[1760], t[1759], t[1758], t[1757], t[1756], t[1755], t[1754], t[1753], t[1752], t[1751], t[1750], t[1749], t[1748], t[1747], t[1746], t[1745], t[1744], t[1743], t[1742], t[1741], t[1740], t[1739], t[1738], t[1737], t[1736], t[1735], t[1734], t[1733], t[1732], t[1731], t[1730], t[1729], t[1728], t[1727], t[1726], t[1725], t[1724], t[1723], t[1722], t[1721], t[1720], t[1719], t[1718], t[1717], t[1716], t[1715], t[1714], t[1713], t[1712], t[1711], t[1710], t[1709], t[1708], t[1707], t[1706], t[1705], t[1704], t[1703], t[1702], t[1701], t[1700], t[1699], t[1698], t[1697], t[1696], t[1695], t[1694], t[1693], t[1692], t[1691], t[1690], t[1689], t[1688], t[1687], t[1686], t[1685], t[1684], t[1683], t[1682], t[1681], t[1680], t[1679], t[1678], t[1677], t[1676], t[1675], t[1674], t[1673], t[1672], t[1671], t[1670], t[1669], t[1668], t[1667], t[1666], t[1665], t[1664], t[1663], t[1662], t[1661], t[1660], t[1659], t[1658], t[1657], t[1656], t[1655], t[1654], t[1653], t[1652], t[1651], t[1650], t[1649], t[1648], t[1647], t[1646], t[1645], t[1644], t[1643], t[1642], t[1641], t[1640], t[1639], t[1638], t[1637], t[1636], t[1635], t[1634], t[1633], t[1632], t[1631], t[1630], t[1629], t[1628], t[1627], t[1626], t[1625], t[1624], t[1623], t[1622], t[1621], t[1620], t[1619], t[1618], t[1617], t[1616], t[1615], t[1614], t[1613], t[1612], t[1611], t[1610], t[1609], t[1608], t[1607], t[1606], t[1605], t[1604], t[1603], t[1602], t[1601], t[1600], t[1599], t[1598], t[1597], t[1596], t[1595], t[1594], t[1593], t[1592], t[1591], t[1590], t[1589], t[1588], t[1587], t[1586], t[1585], t[1584], t[1583], t[1582], t[1581], t[1580], t[1579], t[1578], t[1577], t[1576], t[1575], t[1574], t[1573], t[1572], t[1571], t[1570], t[1569], t[1568], t[1567], t[1566], t[1565], t[1564], t[1563], t[1562], t[1561], t[1560], t[1559], t[1558], t[1557], t[1556], t[1555], t[1554], t[1553], t[1552], t[1551], t[1550], t[1549], t[1548], t[1547], t[1546], t[1545], t[1544], t[1543], t[1542], t[1541], t[1540], t[1539], t[1538], t[1537], t[1536], t[1535], t[1534], t[1533], t[1532], t[1531], t[1530], t[1529], t[1528], t[1527], t[1526], t[1525], t[1524], t[1523], t[1522], t[1521], t[1520], t[1519], t[1518], t[1517], t[1516], t[1515], t[1514], t[1513], t[1512], t[1511], t[1510], t[1509], t[1508], t[1507], t[1506], t[1505], t[1504], t[1503], t[1502], t[1501], t[1500], t[1499], t[1498], t[1497], t[1496], t[1495], t[1494], t[1493], t[1492], t[1491], t[1490], t[1489], t[1488], t[1487], t[1486], t[1485], t[1484], t[1483], t[1482], t[1481], t[1480], t[1479], t[1478], t[1477], t[1476], t[1475], t[1474], t[1473], t[1472], t[1471], t[1470]}));
  Reg1 Reg1_inst(.x({t[1314], t[1315], t[1316], t[1317], t[1318], t[1319], t[1320], t[1321], t[1322], t[1323], t[1324], t[1325], t[1326], t[1327], t[1328], t[1329], t[1330], t[1331], t[1332], t[1333], t[1334], t[1335], t[1336], t[1337], t[1338], t[1339], t[1340], t[1341], t[1342], t[1343], t[1344], t[1345], t[1346], t[1347], t[1348], t[1349], t[1350], t[1351], t[1352], t[1353], t[1354], t[1355], t[1356], t[1357], t[1358], t[1359], t[1360], t[1361], t[1362], t[1363], t[1364], t[1365], t[1366], t[1367], t[1368], t[1369], t[1370], t[1371], t[1372], t[1373], t[1374], t[1375], t[1376], t[1377], t[1378], t[1379], t[1380], t[1381], t[1382], t[1383], t[1384], t[1385], t[1386], t[1387], t[1388], t[1389], t[1390], t[1391], t[1392], t[1393], t[1394], t[1395], t[1396], t[1397], t[1398], t[1399], t[1400], t[1401], t[1402], t[1403], t[1404], t[1405], t[1406], t[1407], t[1408], t[1409], t[1410], t[1411], t[1412], t[1413], t[1414], t[1415], t[1416], t[1417], t[1418], t[1419], t[1420], t[1421], t[1422], t[1423], t[1424], t[1425], t[1426], t[1427], t[1428], t[1429], t[1430], t[1431], t[1432], t[1433], t[1434], t[1435], t[1436], t[1437], t[1438], t[1439], t[1440], t[1441], t[1442], t[1177], t[1176], t[1446], t[1447], t[1448], t[1449], t[1450], t[1444], t[1445], t[1443], x[256], t[1185], t[1184], t[1183], t[1182], t[1181], t[1180], t[1179], t[1178], t[1451], t[1452], t[1453], t[1454], t[1455], t[1456], t[1457], t[1458], t[1461], t[1466], t[1464], t[1459], t[1462], t[1460], t[1463], t[1465], t[1186], t[1187], t[1188], t[1189], t[1190], t[1191], t[1192], t[1193], t[1194], t[1195], t[1196], t[1197], t[1198], t[1199], t[1200], t[1201], t[1202], t[1203], t[1204], t[1205], t[1206], t[1207], t[1208], t[1209], t[1210], t[1211], t[1212], t[1213], t[1214], t[1215], t[1216], t[1217], t[1218], t[1219], t[1220], t[1221], t[1222], t[1223], t[1224], t[1225], t[1226], t[1227], t[1228], t[1229], t[1230], t[1231], t[1232], t[1233], t[1234], t[1235], t[1236], t[1237], t[1238], t[1239], t[1240], t[1241], t[1242], t[1243], t[1244], t[1245], t[1246], t[1247], t[1248], t[1249], t[1250], t[1251], t[1252], t[1253], t[1254], t[1255], t[1256], t[1257], t[1258], t[1259], t[1260], t[1261], t[1262], t[1263], t[1264], t[1265], t[1266], t[1267], t[1268], t[1269], t[1270], t[1271], t[1272], t[1273], t[1274], t[1275], t[1276], t[1277], t[1278], t[1279], t[1280], t[1281], t[1282], t[1283], t[1284], t[1285], t[1286], t[1287], t[1288], t[1289], t[1290], t[1291], t[1292], t[1293], t[1294], t[1295], t[1296], t[1297], t[1298], t[1299], t[1300], t[1301], t[1302], t[1303], t[1304], t[1305], t[1306], t[1307], t[1308], t[1309], t[1310], t[1311], t[1312], t[1313]}), .y({t[663], t[662], t[661], t[660], t[654], t[653], t[652], t[651], t[645], t[644], t[643], t[642], t[636], t[635], t[634], t[633], t[627], t[626], t[625], t[624], t[618], t[617], t[616], t[615], t[609], t[608], t[607], t[606], t[600], t[599], t[598], t[597], t[591], t[590], t[589], t[588], t[582], t[581], t[580], t[579], t[573], t[572], t[571], t[570], t[564], t[563], t[562], t[561], t[555], t[554], t[553], t[552], t[546], t[545], t[544], t[543], t[537], t[536], t[535], t[534], t[528], t[527], t[526], t[525], t[519], t[518], t[517], t[516], t[510], t[509], t[508], t[507], t[501], t[500], t[499], t[498], t[492], t[491], t[490], t[489], t[483], t[482], t[481], t[480], t[474], t[473], t[472], t[471], t[465], t[464], t[463], t[462], t[456], t[455], t[454], t[453], t[447], t[446], t[445], t[444], t[438], t[437], t[436], t[435], t[429], t[428], t[427], t[426], t[420], t[419], t[418], t[417], t[411], t[410], t[409], t[408], t[402], t[401], t[400], t[399], t[393], t[392], t[391], t[390], t[384], t[383], t[382], t[381], t[375], t[374], t[373], t[372], t[366], t[365], t[364], t[363], t[357], t[356], t[355], t[354], t[348], t[347], t[346], t[345], t[339], t[338], t[337], t[336], t[330], t[329], t[328], t[327], t[321], t[320], t[319], t[318], t[312], t[311], t[310], t[309], t[303], t[302], t[301], t[300], t[294], t[293], t[292], t[291], t[285], t[284], t[283], t[282], t[276], t[275], t[274], t[273], t[267], t[266], t[265], t[264], t[258], t[257], t[256], t[255], t[249], t[248], t[247], t[246], t[240], t[239], t[238], t[237], t[231], t[230], t[229], t[228], t[222], t[221], t[220], t[219], t[213], t[212], t[211], t[210], t[204], t[203], t[202], t[201], t[195], t[194], t[193], t[192], t[186], t[185], t[184], t[183], t[177], t[176], t[175], t[174], t[168], t[167], t[166], t[165], t[159], t[158], t[157], t[156], t[150], t[149], t[148], t[147], t[141], t[140], t[139], t[138], t[132], t[131], t[130], t[129], t[123], t[122], t[121], t[120], t[114], t[113], t[112], t[111], t[105], t[104], t[103], t[102], t[96], t[95], t[94], t[93], t[87], t[86], t[85], t[84], t[78], t[77], t[76], t[75], t[69], t[68], t[67], t[66], t[60], t[59], t[58], t[57], t[54], t[51], t[48], t[45], t[42], t[39], t[36], t[33], t[30], t[27], t[24], t[21], t[18], t[15], t[12], t[9], t[6], t[3], t[0]}));
  Reg2 Reg2_inst(.x({t[1889], t[1888], t[1887], t[1886], t[1885], t[1884], t[1883], t[1882], t[1881], t[1880], t[1879], t[1878], t[1877], t[1876], t[1875], t[1874], t[1873], t[1872], t[1871], t[1870], t[1869], t[1868], t[1867], t[1866], t[1865], t[1864], t[1863], t[1862], t[1861], t[1860], t[1859], t[1858], t[1857], t[1856], t[1855], t[1854], t[1853], t[1852], t[1851], t[1850], t[1849], t[1848], t[1847], t[1846], t[1845], t[1844], t[1843], t[1842], t[1841], t[1840], t[1839], t[1838], t[1837], t[1836], t[1835], t[1834], t[1833], t[1832], t[1831], t[1830], t[1829], t[1828], t[1827], t[1826], t[1825], t[1824], t[1823], t[1822], t[1821], t[1820], t[1819], t[1818], t[1817], t[1816], t[1815], t[1814], t[1813], t[1812], t[1811], t[1810], t[1809], t[1808], t[1807], t[1806], t[1805], t[1804], t[1803], t[1802], t[1801], t[1800], t[1799], t[1798], t[1797], t[1796], t[1795], t[1794], t[1793], t[1792], t[1791], t[1790], t[1789], t[1788], t[1787], t[1786], t[1785], t[1784], t[1783], t[1782], t[1781], t[1780], t[1779], t[1778], t[1777], t[1776], t[1775], t[1774], t[1773], t[1772], t[1771], t[1770], t[1769], t[1768], t[1767], t[1766], t[1765], t[1764], t[1763], t[1762], t[1761], t[1760], t[1759], t[1758], t[1757], t[1756], t[1755], t[1754], t[1753], t[1752], t[1751], t[1750], t[1749], t[1748], t[1747], t[1746], t[1745], t[1744], t[1743], t[1742], t[1741], t[1740], t[1739], t[1738], t[1737], t[1736], t[1735], t[1734], t[1733], t[1732], t[1731], t[1730], t[1489], t[1488], t[1487], t[1486], t[1485], t[1484], t[1483], t[1482], t[1481], t[1480], t[1479], t[1478], t[1477], t[1476], t[1475], t[1569], t[1568], t[1567], t[1566], t[1565], t[1564], t[1563], t[1562], t[1561], t[1560], t[1559], t[1558], t[1557], t[1556], t[1555], t[1554], t[1553], t[1552], t[1551], t[1550], t[1549], t[1548], t[1547], t[1546], t[1545], t[1544], t[1543], t[1542], t[1541], t[1540], t[1539], t[1538], t[1537], t[1536], t[1535], t[1494], t[1493], t[1492], t[1491], t[1490], x[256], t[1534], t[1533], t[1532], t[1531], t[1530], t[1529], t[1528], t[1527], t[1526], t[1525], t[1524], t[1523], t[1522], t[1521], t[1520], t[1519], t[1518], t[1517], t[1516], t[1515], t[1514], t[1513], t[1512], t[1511], t[1510], t[1509], t[1508], t[1507], t[1506], t[1505], t[1504], t[1503], t[1502], t[1501], t[1500], t[1499], t[1498], t[1497], t[1496], t[1495], t[1909], t[1908], t[1907], t[1906], t[1905], t[1904], t[1903], t[1902], t[1901], t[1900], t[1899], t[1898], t[1897], t[1896], t[1895], t[1894], t[1893], t[1892], t[1891], t[1890], t[1729], t[1728], t[1727], t[1726], t[1725], t[1724], t[1723], t[1722], t[1721], t[1720], t[1719], t[1718], t[1717], t[1716], t[1715], t[1714], t[1713], t[1712], t[1711], t[1710], t[1709], t[1708], t[1707], t[1706], t[1705], t[1704], t[1703], t[1702], t[1701], t[1700], t[1699], t[1698], t[1697], t[1696], t[1695], t[1694], t[1693], t[1692], t[1691], t[1690], t[1689], t[1688], t[1687], t[1686], t[1685], t[1684], t[1683], t[1682], t[1681], t[1680], t[1679], t[1678], t[1677], t[1676], t[1675], t[1674], t[1673], t[1672], t[1671], t[1670], t[1669], t[1668], t[1667], t[1666], t[1665], t[1664], t[1663], t[1662], t[1661], t[1660], t[1659], t[1658], t[1657], t[1656], t[1655], t[1654], t[1653], t[1652], t[1651], t[1650], t[1649], t[1648], t[1647], t[1646], t[1645], t[1644], t[1643], t[1642], t[1641], t[1640], t[1639], t[1638], t[1637], t[1636], t[1635], t[1634], t[1633], t[1632], t[1631], t[1630], t[1629], t[1628], t[1627], t[1626], t[1625], t[1624], t[1623], t[1622], t[1621], t[1620], t[1619], t[1618], t[1617], t[1616], t[1615], t[1614], t[1613], t[1612], t[1611], t[1610], t[1609], t[1608], t[1607], t[1606], t[1605], t[1604], t[1603], t[1602], t[1601], t[1600], t[1599], t[1598], t[1597], t[1596], t[1595], t[1594], t[1593], t[1592], t[1591], t[1590], t[1589], t[1588], t[1587], t[1586], t[1585], t[1584], t[1583], t[1582], t[1581], t[1580], t[1579], t[1578], t[1577], t[1576], t[1575], t[1574], t[1573], t[1572], t[1571], t[1570]}), .y({t[668], t[667], t[666], t[665], t[664], t[659], t[658], t[657], t[656], t[655], t[650], t[649], t[648], t[647], t[646], t[641], t[640], t[639], t[638], t[637], t[632], t[631], t[630], t[629], t[628], t[623], t[622], t[621], t[620], t[619], t[614], t[613], t[612], t[611], t[610], t[605], t[604], t[603], t[602], t[601], t[596], t[595], t[594], t[593], t[592], t[587], t[586], t[585], t[584], t[583], t[578], t[577], t[576], t[575], t[574], t[569], t[568], t[567], t[566], t[565], t[560], t[559], t[558], t[557], t[556], t[551], t[550], t[549], t[548], t[547], t[542], t[541], t[540], t[539], t[538], t[533], t[532], t[531], t[530], t[529], t[524], t[523], t[522], t[521], t[520], t[515], t[514], t[513], t[512], t[511], t[506], t[505], t[504], t[503], t[502], t[497], t[496], t[495], t[494], t[493], t[488], t[487], t[486], t[485], t[484], t[479], t[478], t[477], t[476], t[475], t[470], t[469], t[468], t[467], t[466], t[461], t[460], t[459], t[458], t[457], t[452], t[451], t[450], t[449], t[448], t[443], t[442], t[441], t[440], t[439], t[434], t[433], t[432], t[431], t[430], t[425], t[424], t[423], t[422], t[421], t[416], t[415], t[414], t[413], t[412], t[407], t[406], t[405], t[404], t[403], t[398], t[397], t[396], t[395], t[394], t[389], t[388], t[387], t[386], t[385], t[380], t[379], t[378], t[377], t[376], t[371], t[370], t[369], t[368], t[367], t[362], t[361], t[360], t[359], t[358], t[353], t[352], t[351], t[350], t[349], t[344], t[343], t[342], t[341], t[340], t[335], t[334], t[333], t[332], t[331], t[326], t[325], t[324], t[323], t[322], t[317], t[316], t[315], t[314], t[313], t[308], t[307], t[306], t[305], t[304], t[299], t[298], t[297], t[296], t[295], t[290], t[289], t[288], t[287], t[286], t[281], t[280], t[279], t[278], t[277], t[272], t[271], t[270], t[269], t[268], t[263], t[262], t[261], t[260], t[259], t[254], t[253], t[252], t[251], t[250], t[245], t[244], t[243], t[242], t[241], t[236], t[235], t[234], t[233], t[232], t[227], t[226], t[225], t[224], t[223], t[218], t[217], t[216], t[215], t[214], t[209], t[208], t[207], t[206], t[205], t[200], t[199], t[198], t[197], t[196], t[191], t[190], t[189], t[188], t[187], t[182], t[181], t[180], t[179], t[178], t[173], t[172], t[171], t[170], t[169], t[164], t[163], t[162], t[161], t[160], t[155], t[154], t[153], t[152], t[151], t[146], t[145], t[144], t[143], t[142], t[137], t[136], t[135], t[134], t[133], t[128], t[127], t[126], t[125], t[124], t[119], t[118], t[117], t[116], t[115], t[110], t[109], t[108], t[107], t[106], t[101], t[100], t[99], t[98], t[97], t[92], t[91], t[90], t[89], t[88], t[83], t[82], t[81], t[80], t[79], t[74], t[73], t[72], t[71], t[70], t[65], t[64], t[63], t[62], t[61], t[56], t[1963], t[1962], t[1961], t[55], t[53], t[1960], t[1959], t[1958], t[52], t[50], t[1957], t[1956], t[1955], t[49], t[47], t[1954], t[1953], t[1952], t[46], t[44], t[1951], t[1950], t[1949], t[43], t[41], t[1948], t[1947], t[1946], t[40], t[38], t[1945], t[1944], t[1943], t[37], t[35], t[1942], t[1941], t[1940], t[34], t[32], t[1939], t[1938], t[1937], t[31], t[29], t[1936], t[1935], t[1934], t[28], t[26], t[1933], t[1932], t[1931], t[25], t[23], t[1930], t[1929], t[1928], t[22], t[20], t[1927], t[1926], t[1925], t[19], t[17], t[1924], t[1923], t[1922], t[16], t[14], t[1921], t[1920], t[1919], t[13], t[11], t[1918], t[1917], t[1916], t[10], t[8], t[1915], t[1914], t[1913], t[7], t[5], t[1912], t[1911], t[1910], t[4], t[2], t[1469], t[1468], t[1467], t[1]}));
  multiplexer #(.WIDTH(129)) multiplexer_inst(.s({t[1470], t[1471], t[1472], t[1473], t[1474], t[1047]}), .d({t[1055], t[1054], t[1053], t[1052], t[1051], t[1050], t[1049], t[1048], t[1063], t[1062], t[1061], t[1060], t[1059], t[1058], t[1057], t[1056], t[1071], t[1070], t[1069], t[1068], t[1067], t[1066], t[1065], t[1064], t[1079], t[1078], t[1077], t[1076], t[1075], t[1074], t[1073], t[1072], t[1087], t[1086], t[1085], t[1084], t[1083], t[1082], t[1081], t[1080], t[1095], t[1094], t[1093], t[1092], t[1091], t[1090], t[1089], t[1088], t[1103], t[1102], t[1101], t[1100], t[1099], t[1098], t[1097], t[1096], t[1111], t[1110], t[1109], t[1108], t[1107], t[1106], t[1105], t[1104], t[1119], t[1118], t[1117], t[1116], t[1115], t[1114], t[1113], t[1112], t[1127], t[1126], t[1125], t[1124], t[1123], t[1122], t[1121], t[1120], t[1135], t[1134], t[1133], t[1132], t[1131], t[1130], t[1129], t[1128], t[1143], t[1142], t[1141], t[1140], t[1139], t[1138], t[1137], t[1136], t[1151], t[1150], t[1149], t[1148], t[1147], t[1146], t[1145], t[1144], t[1159], t[1158], t[1157], t[1156], t[1155], t[1154], t[1153], t[1152], t[1167], t[1166], t[1165], t[1164], t[1163], t[1162], t[1161], t[1160], t[1175], t[1174], t[1173], t[1172], t[1171], t[1170], t[1169], t[1168], t[1470]}), .q({y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], y[8], y[9], y[10], y[11], y[12], y[13], y[14], y[15], y[16], y[17], y[18], y[19], y[20], y[21], y[22], y[23], y[24], y[25], y[26], y[27], y[28], y[29], y[30], y[31], y[32], y[33], y[34], y[35], y[36], y[37], y[38], y[39], y[40], y[41], y[42], y[43], y[44], y[45], y[46], y[47], y[48], y[49], y[50], y[51], y[52], y[53], y[54], y[55], y[56], y[57], y[58], y[59], y[60], y[61], y[62], y[63], y[64], y[65], y[66], y[67], y[68], y[69], y[70], y[71], y[72], y[73], y[74], y[75], y[76], y[77], y[78], y[79], y[80], y[81], y[82], y[83], y[84], y[85], y[86], y[87], y[88], y[89], y[90], y[91], y[92], y[93], y[94], y[95], y[96], y[97], y[98], y[99], y[100], y[101], y[102], y[103], y[104], y[105], y[106], y[107], y[108], y[109], y[110], y[111], y[112], y[113], y[114], y[115], y[116], y[117], y[118], y[119], y[120], y[121], y[122], y[123], y[124], y[125], y[126], y[127], y[128]}));
endmodule

module register_stage(clk, D, Q);
  parameter WIDTH = 8;
  input clk;
  input [WIDTH-1:0] D;
  output [WIDTH-1:0] Q;

  reg [WIDTH-1:0] s_current_state;
  wire [WIDTH-1:0] s_next_state;
  assign s_next_state = D;
  always @ (posedge clk)
  begin
      s_current_state <= s_next_state;
  end
  assign Q = s_current_state;
endmodule

module multiplexer(s, d, q);
  parameter WIDTH = 8;
  input [5:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  muxtree #(.WIDTH(129)) inst_0(.s(s), .d({d[0],d[1],d[2],d[3],d[4],d[5],d[6],d[7],d[8],d[9],d[10],d[11],d[12],d[13],d[14],d[15],d[16],d[17],d[18],d[19],d[20],d[21],d[22],d[23],d[24],d[25],d[26],d[27],d[28],d[29],d[30],d[31],d[32],d[33],d[34],d[35],d[36],d[37],d[38],d[39],d[40],d[41],d[42],d[43],d[44],d[45],d[46],d[47],d[48],d[49],d[50],d[51],d[52],d[53],d[54],d[55],d[56],d[57],d[58],d[59],d[60],d[61],d[62],d[63],d[64],d[65],d[66],d[67],d[68],d[69],d[70],d[71],d[72],d[73],d[74],d[75],d[76],d[77],d[78],d[79],d[80],d[81],d[82],d[83],d[84],d[85],d[86],d[87],d[88],d[89],d[90],d[91],d[92],d[93],d[94],d[95],d[96],d[97],d[98],d[99],d[100],d[101],d[102],d[103],d[104],d[105],d[106],d[107],d[108],d[109],d[110],d[111],d[112],d[113],d[114],d[115],d[116],d[117],d[118],d[119],d[120],d[121],d[122],d[123],d[124],d[125],d[126],d[127],d[128]}), .q({q[0],q[1],q[2],q[3],q[4],q[5],q[6],q[7],q[8],q[9],q[10],q[11],q[12],q[13],q[14],q[15],q[16],q[17],q[18],q[19],q[20],q[21],q[22],q[23],q[24],q[25],q[26],q[27],q[28],q[29],q[30],q[31],q[32],q[33],q[34],q[35],q[36],q[37],q[38],q[39],q[40],q[41],q[42],q[43],q[44],q[45],q[46],q[47],q[48],q[49],q[50],q[51],q[52],q[53],q[54],q[55],q[56],q[57],q[58],q[59],q[60],q[61],q[62],q[63],q[64],q[65],q[66],q[67],q[68],q[69],q[70],q[71],q[72],q[73],q[74],q[75],q[76],q[77],q[78],q[79],q[80],q[81],q[82],q[83],q[84],q[85],q[86],q[87],q[88],q[89],q[90],q[91],q[92],q[93],q[94],q[95],q[96],q[97],q[98],q[99],q[100],q[101],q[102],q[103],q[104],q[105],q[106],q[107],q[108],q[109],q[110],q[111],q[112],q[113],q[114],q[115],q[116],q[117],q[118],q[119],q[120],q[121],q[122],q[123],q[124],q[125],q[126],q[127],q[128]}));
endmodule

module muxtree(s, d, q);
  parameter WIDTH = 8;
  input [5:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  wire [WIDTH-1:0] v0_0;
  wire [WIDTH-1:0] v0_1;
  wire [WIDTH-1:0] v1_0;
  wire [WIDTH-1:0] v1_1;
  wire [WIDTH-1:0] v1_2;
  wire [WIDTH-1:0] v1_3;
  wire [WIDTH-1:0] v2_0;
  wire [WIDTH-1:0] v2_1;
  wire [WIDTH-1:0] v2_2;
  wire [WIDTH-1:0] v2_3;
  wire [WIDTH-1:0] v2_4;
  wire [WIDTH-1:0] v2_5;
  wire [WIDTH-1:0] v2_6;
  wire [WIDTH-1:0] v2_7;
  wire [WIDTH-1:0] v3_0;
  wire [WIDTH-1:0] v3_1;
  wire [WIDTH-1:0] v3_2;
  wire [WIDTH-1:0] v3_3;
  wire [WIDTH-1:0] v3_4;
  wire [WIDTH-1:0] v3_5;
  wire [WIDTH-1:0] v3_6;
  wire [WIDTH-1:0] v3_7;
  wire [WIDTH-1:0] v3_8;
  wire [WIDTH-1:0] v3_9;
  wire [WIDTH-1:0] v3_10;
  wire [WIDTH-1:0] v3_11;
  wire [WIDTH-1:0] v3_12;
  wire [WIDTH-1:0] v3_13;
  wire [WIDTH-1:0] v3_14;
  wire [WIDTH-1:0] v3_15;
  wire [WIDTH-1:0] v4_0;
  wire [WIDTH-1:0] v4_1;
  wire [WIDTH-1:0] v4_2;
  wire [WIDTH-1:0] v4_3;
  wire [WIDTH-1:0] v4_4;
  wire [WIDTH-1:0] v4_5;
  wire [WIDTH-1:0] v4_6;
  wire [WIDTH-1:0] v4_7;
  wire [WIDTH-1:0] v4_8;
  wire [WIDTH-1:0] v4_9;
  wire [WIDTH-1:0] v4_10;
  wire [WIDTH-1:0] v4_11;
  wire [WIDTH-1:0] v4_12;
  wire [WIDTH-1:0] v4_13;
  wire [WIDTH-1:0] v4_14;
  wire [WIDTH-1:0] v4_15;
  wire [WIDTH-1:0] v4_16;
  wire [WIDTH-1:0] v4_17;
  wire [WIDTH-1:0] v4_18;
  wire [WIDTH-1:0] v4_19;
  wire [WIDTH-1:0] v4_20;
  wire [WIDTH-1:0] v4_21;
  wire [WIDTH-1:0] v4_22;
  wire [WIDTH-1:0] v4_23;
  wire [WIDTH-1:0] v4_24;
  wire [WIDTH-1:0] v4_25;
  wire [WIDTH-1:0] v4_26;
  wire [WIDTH-1:0] v4_27;
  wire [WIDTH-1:0] v4_28;
  wire [WIDTH-1:0] v4_29;
  wire [WIDTH-1:0] v4_30;
  wire [WIDTH-1:0] v4_31;

  assign q = s[0] ? v0_1 : {WIDTH{1'b0}};

  assign v0_0 = s[1] ? v1_1 : {WIDTH{1'b0}};
  assign v0_1 = s[1] ? v1_3 : {WIDTH{1'b0}};

  assign v1_0 = s[2] ? {WIDTH{1'b0}} : v2_0;
  assign v1_1 = s[2] ? {WIDTH{1'b0}} : v2_2;
  assign v1_2 = s[2] ? {WIDTH{1'b0}} : v2_4;
  assign v1_3 = s[2] ? {WIDTH{1'b0}} : v2_6;

  assign v2_0 = s[3] ? {WIDTH{1'b0}} : v3_0;
  assign v2_1 = s[3] ? {WIDTH{1'b0}} : v3_2;
  assign v2_2 = s[3] ? {WIDTH{1'b0}} : v3_4;
  assign v2_3 = s[3] ? {WIDTH{1'b0}} : v3_6;
  assign v2_4 = s[3] ? {WIDTH{1'b0}} : v3_8;
  assign v2_5 = s[3] ? {WIDTH{1'b0}} : v3_10;
  assign v2_6 = s[3] ? {WIDTH{1'b0}} : v3_12;
  assign v2_7 = s[3] ? {WIDTH{1'b0}} : v3_14;

  assign v3_0 = s[4] ? {WIDTH{1'b0}} : v4_0;
  assign v3_1 = s[4] ? {WIDTH{1'b0}} : v4_2;
  assign v3_2 = s[4] ? {WIDTH{1'b0}} : v4_4;
  assign v3_3 = s[4] ? {WIDTH{1'b0}} : v4_6;
  assign v3_4 = s[4] ? {WIDTH{1'b0}} : v4_8;
  assign v3_5 = s[4] ? {WIDTH{1'b0}} : v4_10;
  assign v3_6 = s[4] ? {WIDTH{1'b0}} : v4_12;
  assign v3_7 = s[4] ? {WIDTH{1'b0}} : v4_14;
  assign v3_8 = s[4] ? {WIDTH{1'b0}} : v4_16;
  assign v3_9 = s[4] ? {WIDTH{1'b0}} : v4_18;
  assign v3_10 = s[4] ? {WIDTH{1'b0}} : v4_20;
  assign v3_11 = s[4] ? {WIDTH{1'b0}} : v4_22;
  assign v3_12 = s[4] ? {WIDTH{1'b0}} : v4_24;
  assign v3_13 = s[4] ? {WIDTH{1'b0}} : v4_26;
  assign v3_14 = s[4] ? {WIDTH{1'b0}} : v4_28;
  assign v3_15 = s[4] ? {WIDTH{1'b0}} : v4_30;

  assign v4_0 = {WIDTH{1'b0}};
  assign v4_1 = {WIDTH{1'b0}};
  assign v4_2 = {WIDTH{1'b0}};
  assign v4_3 = {WIDTH{1'b0}};
  assign v4_4 = {WIDTH{1'b0}};
  assign v4_5 = {WIDTH{1'b0}};
  assign v4_6 = {WIDTH{1'b0}};
  assign v4_7 = {WIDTH{1'b0}};
  assign v4_8 = {WIDTH{1'b0}};
  assign v4_9 = {WIDTH{1'b0}};
  assign v4_10 = {WIDTH{1'b0}};
  assign v4_11 = {WIDTH{1'b0}};
  assign v4_12 = {WIDTH{1'b0}};
  assign v4_13 = {WIDTH{1'b0}};
  assign v4_14 = {WIDTH{1'b0}};
  assign v4_15 = {WIDTH{1'b0}};
  assign v4_16 = {WIDTH{1'b0}};
  assign v4_17 = {WIDTH{1'b0}};
  assign v4_18 = {WIDTH{1'b0}};
  assign v4_19 = {WIDTH{1'b0}};
  assign v4_20 = {WIDTH{1'b0}};
  assign v4_21 = {WIDTH{1'b0}};
  assign v4_22 = {WIDTH{1'b0}};
  assign v4_23 = {WIDTH{1'b0}};
  assign v4_24 = s[5] ? d : {WIDTH{1'b0}};
  assign v4_25 = {WIDTH{1'b0}};
  assign v4_26 = {WIDTH{1'b0}};
  assign v4_27 = {WIDTH{1'b0}};
  assign v4_28 = {WIDTH{1'b0}};
  assign v4_29 = {WIDTH{1'b0}};
  assign v4_30 = {WIDTH{1'b0}};
  assign v4_31 = {WIDTH{1'b0}};

endmodule

