/* modified netlist. Source: module AES in file ../CaseStudies/07_AES128_byte_serial_encryption/FPGA_based/AES_synthesis.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module AES_GHPC_ClockGating_d1 (clk, start, plaintext_s0, key_s0, plaintext_s1, key_s1, Fresh, done, ciphertext_s0, ciphertext_s1, Synch);
    input clk ;
    input start ;
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [39:0] Fresh ;
    output done ;
    output [127:0] ciphertext_s0 ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire \ctrl/CSenRC_405 ;
    wire intFinal ;
    wire nReset_407 ;
    wire enKS ;
    wire intselXOR_425 ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD ;
    wire \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD ;
    wire \ctrl/finalStep1 ;
    wire \ctrl/seq4/GEN[1].SFF/QD ;
    wire \ctrl/seq4/GEN[0].SFF/QD ;
    wire \ctrl/seq6/GEN[4].SFF/QD ;
    wire \ctrl/seq6/GEN[3].SFF/QD ;
    wire \ctrl/seq6/GEN[2].SFF/QD ;
    wire \ctrl/seq6/GEN[1].SFF/QD ;
    wire \ctrl/seq6/GEN[0].SFF/QD ;
    wire \ctrl/CSselMC_835 ;
    wire \ctrl/seq4/GEN[0].SFF/Q_836 ;
    wire \ctrl/seq4/GEN[1].SFF/Q_837 ;
    wire \ctrl/seq6/GEN[1].SFF/Q_838 ;
    wire \ctrl/seq6/GEN[2].SFF/Q_839 ;
    wire \ctrl/seq6/GEN[3].SFF/Q_840 ;
    wire \ctrl/seq6/GEN[0].SFF/Q_841 ;
    wire \ctrl/seq6/GEN[4].SFF/Q_842 ;
    wire \calcRCon/nReset_inv ;
    wire \calcRCon/MSB_s_current_state[0]_XOR_21_o ;
    wire \calcRCon/MSB_s_current_state[2]_XOR_20_o ;
    wire \calcRCon/MSB_s_current_state[3]_XOR_19_o ;
    wire N01 ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N10 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ;
    wire \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N30 ;
    wire N32 ;
    wire \ctrl/CSselMC_rstpot_1330 ;
    wire nReset_rstpot ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N50 ;
    wire nReset_1_1341 ;
    wire \ctrl/CSselMC_1_1342 ;
    wire [7:0] StateInMC ;
    wire [7:0] SboxIn ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] SboxOut ;
    wire [7:0] \stateArray/input_MC ;
    wire [7:0] \KeyArray/inS00ser ;
    wire [7:0] \calcRCon/s_current_state ;
    wire [3:0] \Inst_bSbox/b7 ;
    wire [3:0] \Inst_bSbox/b6 ;
    wire [3:0] \Inst_bSbox/b5 ;
    wire [3:0] \Inst_bSbox/b4 ;
    wire [3:0] \Inst_bSbox/b3 ;
    wire [3:0] \Inst_bSbox/b2 ;
    wire [3:0] \Inst_bSbox/b1 ;
    wire [3:0] \Inst_bSbox/b0 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2260 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[7].inS00serInst ( .I0 ({key_s1[127], key_s0[127]}), .I1 ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }), .I2 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2142, \KeyArray/inS00ser [7]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[6].inS00serInst ( .I0 ({key_s1[126], key_s0[126]}), .I1 ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }), .I2 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2144, \KeyArray/inS00ser [6]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[5].inS00serInst ( .I0 ({key_s1[125], key_s0[125]}), .I1 ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }), .I2 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2146, \KeyArray/inS00ser [5]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[4].inS00serInst ( .I0 ({key_s1[124], key_s0[124]}), .I1 ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }), .I2 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2148, \KeyArray/inS00ser [4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[3].inS00serInst ( .I0 ({key_s1[123], key_s0[123]}), .I1 ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }), .I2 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2150, \KeyArray/inS00ser [3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[2].inS00serInst ( .I0 ({key_s1[122], key_s0[122]}), .I1 ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }), .I2 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2152, \KeyArray/inS00ser [2]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[1].inS00serInst ( .I0 ({key_s1[121], key_s0[121]}), .I1 ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }), .I2 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2154, \KeyArray/inS00ser [1]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h3CCCAAAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CCCAAAA ) ) \KeyArray/gen00ser[0].inS00serInst ( .I0 ({key_s1[120], key_s0[120]}), .I1 ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }), .I2 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I3 ({1'b0, intselXOR_425}), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_2156, \KeyArray/inS00ser [0]}) ) ;
    LUT5 #( .INIT ( 32'h00800000 ) ) done1 ( .I0 (intFinal), .I1 (nReset_407), .I2 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I3 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I4 (\ctrl/finalStep1 ), .O (done) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<7>1 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .O ({new_AGEMA_signal_1351, StateOutXORroundKey[7]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<6>1 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .O ({new_AGEMA_signal_1354, StateOutXORroundKey[6]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<5>1 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .O ({new_AGEMA_signal_1357, StateOutXORroundKey[5]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<4>1 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .O ({new_AGEMA_signal_1360, StateOutXORroundKey[4]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<3>1 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .O ({new_AGEMA_signal_1363, StateOutXORroundKey[3]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<2>1 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .O ({new_AGEMA_signal_1366, StateOutXORroundKey[2]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<1>1 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .O ({new_AGEMA_signal_1369, StateOutXORroundKey[1]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \StateOutXORroundKey<0>1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .O ({new_AGEMA_signal_1372, StateOutXORroundKey[0]}) ) ;
    LUT3 #( .INIT ( 8'hE0 ) ) \ctrl/intSelXOR1 ( .I0 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I1 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I2 (nReset_407), .O (selXOR) ) ;
    LUT5 #( .INIT ( 32'h00000001 ) ) \ctrl/finalStep11 ( .I0 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I1 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I2 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I3 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I4 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .O (\ctrl/finalStep1 ) ) ;
    LUT3 #( .INIT ( 8'h20 ) ) \ctrl/seq4/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I1 (\ctrl/finalStep1 ), .I2 (nReset_407), .O (\ctrl/seq4/GEN[1].SFF/QD ) ) ;
    LUT3 #( .INIT ( 8'hDF ) ) \ctrl/seq4/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/finalStep1 ), .I2 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .O (\ctrl/seq4/GEN[0].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \ctrl/seq6/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .O (\ctrl/seq6/GEN[4].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/seq6/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .I1 (nReset_407), .O (\ctrl/seq6/GEN[3].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \ctrl/seq6/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .O (\ctrl/seq6/GEN[2].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/seq6/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I1 (nReset_407), .O (\ctrl/seq6/GEN[1].SFF/QD ) ) ;
    LUT3 #( .INIT ( 8'h9F ) ) \ctrl/seq6/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I1 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I2 (nReset_407), .O (\ctrl/seq6/GEN[0].SFF/QD ) ) ;
    LUT2 #( .INIT ( 4'h8 ) ) \ctrl/selMC1 ( .I0 (\ctrl/CSselMC_835 ), .I1 (nReset_407), .O (selMC) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[0]_XOR_21_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [0]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[0]_XOR_21_o ) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[3]_XOR_19_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [3]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[3]_XOR_19_o ) ) ;
    LUT2 #( .INIT ( 4'h6 ) ) \calcRCon/Mxor_MSB_s_current_state[2]_XOR_20_o_xo<0>1 ( .I0 (\calcRCon/s_current_state [2]), .I1 (\calcRCon/s_current_state [7]), .O (\calcRCon/MSB_s_current_state[2]_XOR_20_o ) ) ;
    LUT4 #( .INIT ( 16'h8000 ) ) \calcRCon/final<1>1 ( .I0 (\calcRCon/s_current_state [1]), .I1 (\calcRCon/s_current_state [2]), .I2 (\calcRCon/s_current_state [4]), .I3 (\calcRCon/s_current_state [5]), .O (intFinal) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[0].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[88], ciphertext_s0[88]}), .O ({new_AGEMA_signal_1374, N01}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[0].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[24], ciphertext_s0[24]}), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({ciphertext_s1[56], ciphertext_s0[56]}), .I4 ({ciphertext_s1[31], ciphertext_s0[31]}), .I5 ({new_AGEMA_signal_1374, N01}), .O ({new_AGEMA_signal_1893, StateInMC[0]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[1].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1377, N2}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[1].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[57], ciphertext_s0[57]}), .I3 ({ciphertext_s1[121], ciphertext_s0[121]}), .I4 ({ciphertext_s1[89], ciphertext_s0[89]}), .I5 ({new_AGEMA_signal_1377, N2}), .O ({new_AGEMA_signal_1894, StateInMC[1]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[2].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[90], ciphertext_s0[90]}), .I1 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1380, N4}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[2].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({ciphertext_s1[25], ciphertext_s0[25]}), .I4 ({ciphertext_s1[122], ciphertext_s0[122]}), .I5 ({new_AGEMA_signal_1380, N4}), .O ({new_AGEMA_signal_1895, StateInMC[2]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[3].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[26], ciphertext_s0[26]}), .O ({new_AGEMA_signal_1382, N6}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[3].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[27], ciphertext_s0[27]}), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[59], ciphertext_s0[59]}), .I5 ({new_AGEMA_signal_1382, N6}), .O ({new_AGEMA_signal_1896, StateInMC[3]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \MUX_StateInMC/gen_mux[4].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[92], ciphertext_s0[92]}), .I1 ({ciphertext_s1[60], ciphertext_s0[60]}), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[127], ciphertext_s0[127]}), .O ({new_AGEMA_signal_1385, N8}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[4].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[28], ciphertext_s0[28]}), .I2 ({ciphertext_s1[27], ciphertext_s0[27]}), .I3 ({ciphertext_s1[124], ciphertext_s0[124]}), .I4 ({ciphertext_s1[123], ciphertext_s0[123]}), .I5 ({new_AGEMA_signal_1385, N8}), .O ({new_AGEMA_signal_1897, StateInMC[4]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[5].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[93], ciphertext_s0[93]}), .I1 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1388, N10}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[5].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[28], ciphertext_s0[28]}), .I3 ({ciphertext_s1[124], ciphertext_s0[124]}), .I4 ({ciphertext_s1[125], ciphertext_s0[125]}), .I5 ({new_AGEMA_signal_1388, N10}), .O ({new_AGEMA_signal_1898, StateInMC[5]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[6].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[94], ciphertext_s0[94]}), .I1 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1391, N12}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[6].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({ciphertext_s1[29], ciphertext_s0[29]}), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({new_AGEMA_signal_1391, N12}), .O ({new_AGEMA_signal_1899, StateInMC[6]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MUX_StateInMC/gen_mux[7].mux_inst/Mmux_Q1_SW0 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1394, N14}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \MUX_StateInMC/gen_mux[7].mux_inst/Mmux_Q1 ( .I0 ({1'b0, intFinal}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[127], ciphertext_s0[127]}), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({new_AGEMA_signal_1394, N14}), .O ({new_AGEMA_signal_1900, StateInMC[7]}) ) ;
    LUT4 #( .INIT ( 16'h7FFF ) ) intselXOR_SW0 ( .I0 (\calcRCon/s_current_state [2]), .I1 (\calcRCon/s_current_state [7]), .I2 (\calcRCon/s_current_state [3]), .I3 (\calcRCon/s_current_state [0]), .O (N16) ) ;
    LUT6 #( .INIT ( 64'hFFFFFFFE00000000 ) ) intselXOR ( .I0 (\calcRCon/s_current_state [6]), .I1 (\calcRCon/s_current_state [4]), .I2 (\calcRCon/s_current_state [5]), .I3 (\calcRCon/s_current_state [1]), .I4 (N16), .I5 (selXOR), .O (intselXOR_425) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[56], ciphertext_s0[56]}), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1396, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1396, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[120], ciphertext_s0[120]}), .O ({new_AGEMA_signal_1901, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1397, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1397, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[89], ciphertext_s0[89]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[122], ciphertext_s0[122]}), .O ({new_AGEMA_signal_1902, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1399, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1399, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .I3 ({ciphertext_s1[92], ciphertext_s0[92]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .O ({new_AGEMA_signal_1903, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1401, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1401, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .I3 ({ciphertext_s1[93], ciphertext_s0[93]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[126], ciphertext_s0[126]}), .O ({new_AGEMA_signal_1904, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1402, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1402, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[94], ciphertext_s0[94]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .O ({new_AGEMA_signal_1905, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[120], ciphertext_s0[120]}), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .O ({new_AGEMA_signal_1403, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1403, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[88], ciphertext_s0[88]}), .O ({new_AGEMA_signal_1906, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[26], ciphertext_s0[26]}), .I2 ({ciphertext_s1[89], ciphertext_s0[89]}), .O ({new_AGEMA_signal_1405, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1405, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[57], ciphertext_s0[57]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[90], ciphertext_s0[90]}), .O ({new_AGEMA_signal_1907, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[125], ciphertext_s0[125]}), .I1 ({ciphertext_s1[29], ciphertext_s0[29]}), .I2 ({ciphertext_s1[92], ciphertext_s0[92]}), .O ({new_AGEMA_signal_1406, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1406, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .I3 ({ciphertext_s1[60], ciphertext_s0[60]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .O ({new_AGEMA_signal_1908, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[126], ciphertext_s0[126]}), .I1 ({ciphertext_s1[30], ciphertext_s0[30]}), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .O ({new_AGEMA_signal_1407, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1407, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .I3 ({ciphertext_s1[61], ciphertext_s0[61]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[94], ciphertext_s0[94]}), .O ({new_AGEMA_signal_1909, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[127], ciphertext_s0[127]}), .I1 ({ciphertext_s1[31], ciphertext_s0[31]}), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .O ({new_AGEMA_signal_1408, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1408, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .I3 ({ciphertext_s1[62], ciphertext_s0[62]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .O ({new_AGEMA_signal_1910, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[120], ciphertext_s0[120]}), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1409, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1409, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .I3 ({ciphertext_s1[31], ciphertext_s0[31]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[56], ciphertext_s0[56]}), .O ({new_AGEMA_signal_1911, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .O ({new_AGEMA_signal_1411, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1411, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[25], ciphertext_s0[25]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[58], ciphertext_s0[58]}), .O ({new_AGEMA_signal_1912, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[93], ciphertext_s0[93]}), .I1 ({ciphertext_s1[125], ciphertext_s0[125]}), .I2 ({ciphertext_s1[60], ciphertext_s0[60]}), .O ({new_AGEMA_signal_1412, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1412, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[29], ciphertext_s0[29]}), .I3 ({ciphertext_s1[28], ciphertext_s0[28]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1913, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[94], ciphertext_s0[94]}), .I1 ({ciphertext_s1[126], ciphertext_s0[126]}), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .O ({new_AGEMA_signal_1413, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1413, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[29], ciphertext_s0[29]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1914, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({ciphertext_s1[95], ciphertext_s0[95]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .O ({new_AGEMA_signal_1414, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFAFAD2785050D278 ) , .MASK ( 6'b010001 ), .INIT2 ( 64'hFAFAD2785050D278 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q12 ( .I0 ({1'b0, selMC}), .I1 ({new_AGEMA_signal_1414, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 }), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[30], ciphertext_s0[30]}), .I4 ({1'b0, intFinal}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .O ({new_AGEMA_signal_1915, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I1 ({1'b0, \calcRCon/s_current_state [0]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1415, N18}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I1 ({1'b0, \calcRCon/s_current_state [1]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1416, N20}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I1 ({1'b0, \calcRCon/s_current_state [2]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1417, N22}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I1 ({1'b0, \calcRCon/s_current_state [3]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1418, N24}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I1 ({1'b0, \calcRCon/s_current_state [4]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1419, N26}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I1 ({1'b0, \calcRCon/s_current_state [5]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1420, N28}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I1 ({1'b0, \calcRCon/s_current_state [6]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1421, N30}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h95 ) , .MASK ( 3'b110 ), .INIT2 ( 8'hAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I1 ({1'b0, \calcRCon/s_current_state [7]}), .I2 ({1'b0, \ctrl/CSenRC_405 }), .O ({new_AGEMA_signal_1422, N32}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<5>1 ( .I0 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I1 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1424, SboxIn[5]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<4>1 ( .I0 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I1 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I2 ({ciphertext_s1[124], ciphertext_s0[124]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1426, SboxIn[4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<3>1 ( .I0 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I1 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1428, SboxIn[3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<2>1 ( .I0 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I1 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1430, SboxIn[2]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<1>1 ( .I0 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I1 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1432, SboxIn[1]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<0>1 ( .I0 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I1 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({1'b0, \ctrl/CSselMC_1_1342 }), .I4 ({1'b0, nReset_1_1341}), .O ({new_AGEMA_signal_1434, SboxIn[0]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<7>1 ( .I0 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I1 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({1'b0, \ctrl/CSselMC_835 }), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_1436, SboxIn[7]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAA3C3C3C ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAA3C3C3C ) ) \SboxIn<6>1 ( .I0 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I1 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I2 ({ciphertext_s1[126], ciphertext_s0[126]}), .I3 ({1'b0, \ctrl/CSselMC_835 }), .I4 ({1'b0, nReset_407}), .O ({new_AGEMA_signal_1438, SboxIn[6]}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2156, \KeyArray/inS00ser [0]}), .O ({new_AGEMA_signal_2237, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2154, \KeyArray/inS00ser [1]}), .O ({new_AGEMA_signal_2238, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2152, \KeyArray/inS00ser [2]}), .O ({new_AGEMA_signal_2239, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2150, \KeyArray/inS00ser [3]}), .O ({new_AGEMA_signal_2240, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2148, \KeyArray/inS00ser [4]}), .O ({new_AGEMA_signal_2241, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2146, \KeyArray/inS00ser [5]}), .O ({new_AGEMA_signal_2242, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2144, \KeyArray/inS00ser [6]}), .O ({new_AGEMA_signal_2243, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBF80 ) , .MASK ( 4'b0110 ), .INIT2 ( 16'hBF80 ) ) \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, nReset_407}), .I3 ({new_AGEMA_signal_2142, \KeyArray/inS00ser [7]}), .O ({new_AGEMA_signal_2244, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[57], ciphertext_s0[57]}), .I5 ({ciphertext_s1[25], ciphertext_s0[25]}), .O ({new_AGEMA_signal_1440, N34}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[89], ciphertext_s0[89]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1440, N34}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[121], ciphertext_s0[121]}), .O ({new_AGEMA_signal_1916, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[122], ciphertext_s0[122]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[59], ciphertext_s0[59]}), .I5 ({ciphertext_s1[27], ciphertext_s0[27]}), .O ({new_AGEMA_signal_1443, N36}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[91], ciphertext_s0[91]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1443, N36}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[123], ciphertext_s0[123]}), .O ({new_AGEMA_signal_1917, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[127], ciphertext_s0[127]}), .I2 ({ciphertext_s1[91], ciphertext_s0[91]}), .I3 ({ciphertext_s1[95], ciphertext_s0[95]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[28], ciphertext_s0[28]}), .O ({new_AGEMA_signal_1446, N38}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[92], ciphertext_s0[92]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1446, N38}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[124], ciphertext_s0[124]}), .O ({new_AGEMA_signal_1918, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[88], ciphertext_s0[88]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[56], ciphertext_s0[56]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[25], ciphertext_s0[25]}), .O ({new_AGEMA_signal_1447, N40}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[57], ciphertext_s0[57]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1447, N40}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[89], ciphertext_s0[89]}), .O ({new_AGEMA_signal_1919, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[90], ciphertext_s0[90]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[58], ciphertext_s0[58]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[27], ciphertext_s0[27]}), .O ({new_AGEMA_signal_1448, N42}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[59], ciphertext_s0[59]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1448, N42}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[91], ciphertext_s0[91]}), .O ({new_AGEMA_signal_1920, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[91], ciphertext_s0[91]}), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[63], ciphertext_s0[63]}), .I5 ({ciphertext_s1[28], ciphertext_s0[28]}), .O ({new_AGEMA_signal_1449, N44}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[60], ciphertext_s0[60]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1449, N44}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[92], ciphertext_s0[92]}), .O ({new_AGEMA_signal_1921, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[121], ciphertext_s0[121]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[24], ciphertext_s0[24]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1450, N46}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[25], ciphertext_s0[25]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1450, N46}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[57], ciphertext_s0[57]}), .O ({new_AGEMA_signal_1922, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[123], ciphertext_s0[123]}), .I1 ({ciphertext_s1[91], ciphertext_s0[91]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[26], ciphertext_s0[26]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1451, N48}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[27], ciphertext_s0[27]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1451, N48}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[59], ciphertext_s0[59]}), .O ({new_AGEMA_signal_1923, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13_SW0 ( .I0 ({ciphertext_s1[124], ciphertext_s0[124]}), .I1 ({ciphertext_s1[92], ciphertext_s0[92]}), .I2 ({ciphertext_s1[59], ciphertext_s0[59]}), .I3 ({ciphertext_s1[63], ciphertext_s0[63]}), .I4 ({ciphertext_s1[27], ciphertext_s0[27]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .O ({new_AGEMA_signal_1452, N50}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE6EAAAAA262AAAAA ) , .MASK ( 6'b010110 ), .INIT2 ( 64'hE6EAAAAA262AAAAA ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q13 ( .I0 ({ciphertext_s1[28], ciphertext_s0[28]}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({1'b0, intFinal}), .I3 ({new_AGEMA_signal_1452, N50}), .I4 ({1'b0, nReset_407}), .I5 ({ciphertext_s1[60], ciphertext_s0[60]}), .O ({new_AGEMA_signal_1924, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[88], plaintext_s0[88]}), .I2 ({ciphertext_s1[80], ciphertext_s0[80]}), .O ({new_AGEMA_signal_1455, \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[89], plaintext_s0[89]}), .I2 ({ciphertext_s1[81], ciphertext_s0[81]}), .O ({new_AGEMA_signal_1458, \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[90], plaintext_s0[90]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .O ({new_AGEMA_signal_1461, \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[91], plaintext_s0[91]}), .I2 ({ciphertext_s1[83], ciphertext_s0[83]}), .O ({new_AGEMA_signal_1464, \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[92], plaintext_s0[92]}), .I2 ({ciphertext_s1[84], ciphertext_s0[84]}), .O ({new_AGEMA_signal_1467, \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[93], plaintext_s0[93]}), .I2 ({ciphertext_s1[85], ciphertext_s0[85]}), .O ({new_AGEMA_signal_1470, \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[94], plaintext_s0[94]}), .I2 ({ciphertext_s1[86], ciphertext_s0[86]}), .O ({new_AGEMA_signal_1473, \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[95], plaintext_s0[95]}), .I2 ({ciphertext_s1[87], ciphertext_s0[87]}), .O ({new_AGEMA_signal_1476, \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[80], plaintext_s0[80]}), .I2 ({ciphertext_s1[72], ciphertext_s0[72]}), .O ({new_AGEMA_signal_1479, \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[81], plaintext_s0[81]}), .I2 ({ciphertext_s1[73], ciphertext_s0[73]}), .O ({new_AGEMA_signal_1482, \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[82], plaintext_s0[82]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .O ({new_AGEMA_signal_1485, \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[83], plaintext_s0[83]}), .I2 ({ciphertext_s1[75], ciphertext_s0[75]}), .O ({new_AGEMA_signal_1488, \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[84], plaintext_s0[84]}), .I2 ({ciphertext_s1[76], ciphertext_s0[76]}), .O ({new_AGEMA_signal_1491, \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[85], plaintext_s0[85]}), .I2 ({ciphertext_s1[77], ciphertext_s0[77]}), .O ({new_AGEMA_signal_1494, \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[86], plaintext_s0[86]}), .I2 ({ciphertext_s1[78], ciphertext_s0[78]}), .O ({new_AGEMA_signal_1497, \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[87], plaintext_s0[87]}), .I2 ({ciphertext_s1[79], ciphertext_s0[79]}), .O ({new_AGEMA_signal_1500, \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[72], plaintext_s0[72]}), .I2 ({ciphertext_s1[64], ciphertext_s0[64]}), .O ({new_AGEMA_signal_1503, \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[73], plaintext_s0[73]}), .I2 ({ciphertext_s1[65], ciphertext_s0[65]}), .O ({new_AGEMA_signal_1506, \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[74], plaintext_s0[74]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .O ({new_AGEMA_signal_1509, \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[75], plaintext_s0[75]}), .I2 ({ciphertext_s1[67], ciphertext_s0[67]}), .O ({new_AGEMA_signal_1512, \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[76], plaintext_s0[76]}), .I2 ({ciphertext_s1[68], ciphertext_s0[68]}), .O ({new_AGEMA_signal_1515, \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[77], plaintext_s0[77]}), .I2 ({ciphertext_s1[69], ciphertext_s0[69]}), .O ({new_AGEMA_signal_1518, \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[78], plaintext_s0[78]}), .I2 ({ciphertext_s1[70], ciphertext_s0[70]}), .O ({new_AGEMA_signal_1521, \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hE4 ) , .MASK ( 3'b001 ), .INIT2 ( 8'hE4 ) ) \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({plaintext_s1[79], plaintext_s0[79]}), .I2 ({ciphertext_s1[71], ciphertext_s0[71]}), .O ({new_AGEMA_signal_1524, \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[120], ciphertext_s0[120]}), .I3 ({ciphertext_s1[112], ciphertext_s0[112]}), .I4 ({plaintext_s1[120], plaintext_s0[120]}), .O ({new_AGEMA_signal_1927, \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[121], ciphertext_s0[121]}), .I3 ({ciphertext_s1[113], ciphertext_s0[113]}), .I4 ({plaintext_s1[121], plaintext_s0[121]}), .O ({new_AGEMA_signal_1930, \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[114], ciphertext_s0[114]}), .I4 ({plaintext_s1[122], plaintext_s0[122]}), .O ({new_AGEMA_signal_1933, \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[123], ciphertext_s0[123]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({plaintext_s1[123], plaintext_s0[123]}), .O ({new_AGEMA_signal_1936, \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[124], ciphertext_s0[124]}), .I3 ({ciphertext_s1[116], ciphertext_s0[116]}), .I4 ({plaintext_s1[124], plaintext_s0[124]}), .O ({new_AGEMA_signal_1939, \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[125], ciphertext_s0[125]}), .I3 ({ciphertext_s1[117], ciphertext_s0[117]}), .I4 ({plaintext_s1[125], plaintext_s0[125]}), .O ({new_AGEMA_signal_1942, \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[126], ciphertext_s0[126]}), .I3 ({ciphertext_s1[118], ciphertext_s0[118]}), .I4 ({plaintext_s1[126], plaintext_s0[126]}), .O ({new_AGEMA_signal_1945, \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[127], ciphertext_s0[127]}), .I3 ({ciphertext_s1[119], ciphertext_s0[119]}), .I4 ({plaintext_s1[127], plaintext_s0[127]}), .O ({new_AGEMA_signal_1948, \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[112], ciphertext_s0[112]}), .I3 ({ciphertext_s1[104], ciphertext_s0[104]}), .I4 ({plaintext_s1[112], plaintext_s0[112]}), .O ({new_AGEMA_signal_1951, \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[113], ciphertext_s0[113]}), .I3 ({ciphertext_s1[105], ciphertext_s0[105]}), .I4 ({plaintext_s1[113], plaintext_s0[113]}), .O ({new_AGEMA_signal_1954, \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[106], ciphertext_s0[106]}), .I4 ({plaintext_s1[114], plaintext_s0[114]}), .O ({new_AGEMA_signal_1957, \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[115], ciphertext_s0[115]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({plaintext_s1[115], plaintext_s0[115]}), .O ({new_AGEMA_signal_1960, \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[116], ciphertext_s0[116]}), .I3 ({ciphertext_s1[108], ciphertext_s0[108]}), .I4 ({plaintext_s1[116], plaintext_s0[116]}), .O ({new_AGEMA_signal_1963, \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[117], ciphertext_s0[117]}), .I3 ({ciphertext_s1[109], ciphertext_s0[109]}), .I4 ({plaintext_s1[117], plaintext_s0[117]}), .O ({new_AGEMA_signal_1966, \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[118], ciphertext_s0[118]}), .I3 ({ciphertext_s1[110], ciphertext_s0[110]}), .I4 ({plaintext_s1[118], plaintext_s0[118]}), .O ({new_AGEMA_signal_1969, \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[119], ciphertext_s0[119]}), .I3 ({ciphertext_s1[111], ciphertext_s0[111]}), .I4 ({plaintext_s1[119], plaintext_s0[119]}), .O ({new_AGEMA_signal_1972, \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[104], ciphertext_s0[104]}), .I3 ({ciphertext_s1[96], ciphertext_s0[96]}), .I4 ({plaintext_s1[104], plaintext_s0[104]}), .O ({new_AGEMA_signal_1975, \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[105], ciphertext_s0[105]}), .I3 ({ciphertext_s1[97], ciphertext_s0[97]}), .I4 ({plaintext_s1[105], plaintext_s0[105]}), .O ({new_AGEMA_signal_1978, \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[98], ciphertext_s0[98]}), .I4 ({plaintext_s1[106], plaintext_s0[106]}), .O ({new_AGEMA_signal_1981, \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[107], ciphertext_s0[107]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({plaintext_s1[107], plaintext_s0[107]}), .O ({new_AGEMA_signal_1984, \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[108], ciphertext_s0[108]}), .I3 ({ciphertext_s1[100], ciphertext_s0[100]}), .I4 ({plaintext_s1[108], plaintext_s0[108]}), .O ({new_AGEMA_signal_1987, \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[109], ciphertext_s0[109]}), .I3 ({ciphertext_s1[101], ciphertext_s0[101]}), .I4 ({plaintext_s1[109], plaintext_s0[109]}), .O ({new_AGEMA_signal_1990, \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[110], ciphertext_s0[110]}), .I3 ({ciphertext_s1[102], ciphertext_s0[102]}), .I4 ({plaintext_s1[110], plaintext_s0[110]}), .O ({new_AGEMA_signal_1993, \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[111], ciphertext_s0[111]}), .I3 ({ciphertext_s1[103], ciphertext_s0[103]}), .I4 ({plaintext_s1[111], plaintext_s0[111]}), .O ({new_AGEMA_signal_1996, \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[40], ciphertext_s0[40]}), .I3 ({ciphertext_s1[48], ciphertext_s0[48]}), .I4 ({plaintext_s1[56], plaintext_s0[56]}), .O ({new_AGEMA_signal_2000, \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[41], ciphertext_s0[41]}), .I3 ({ciphertext_s1[49], ciphertext_s0[49]}), .I4 ({plaintext_s1[57], plaintext_s0[57]}), .O ({new_AGEMA_signal_2004, \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[50], ciphertext_s0[50]}), .I4 ({plaintext_s1[58], plaintext_s0[58]}), .O ({new_AGEMA_signal_2008, \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[43], ciphertext_s0[43]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({plaintext_s1[59], plaintext_s0[59]}), .O ({new_AGEMA_signal_2012, \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[44], ciphertext_s0[44]}), .I3 ({ciphertext_s1[52], ciphertext_s0[52]}), .I4 ({plaintext_s1[60], plaintext_s0[60]}), .O ({new_AGEMA_signal_2016, \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[45], ciphertext_s0[45]}), .I3 ({ciphertext_s1[53], ciphertext_s0[53]}), .I4 ({plaintext_s1[61], plaintext_s0[61]}), .O ({new_AGEMA_signal_2020, \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[46], ciphertext_s0[46]}), .I3 ({ciphertext_s1[54], ciphertext_s0[54]}), .I4 ({plaintext_s1[62], plaintext_s0[62]}), .O ({new_AGEMA_signal_2024, \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[47], ciphertext_s0[47]}), .I3 ({ciphertext_s1[55], ciphertext_s0[55]}), .I4 ({plaintext_s1[63], plaintext_s0[63]}), .O ({new_AGEMA_signal_2028, \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[32], ciphertext_s0[32]}), .I3 ({ciphertext_s1[40], ciphertext_s0[40]}), .I4 ({plaintext_s1[48], plaintext_s0[48]}), .O ({new_AGEMA_signal_2031, \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[33], ciphertext_s0[33]}), .I3 ({ciphertext_s1[41], ciphertext_s0[41]}), .I4 ({plaintext_s1[49], plaintext_s0[49]}), .O ({new_AGEMA_signal_2034, \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[42], ciphertext_s0[42]}), .I4 ({plaintext_s1[50], plaintext_s0[50]}), .O ({new_AGEMA_signal_2037, \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[35], ciphertext_s0[35]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({plaintext_s1[51], plaintext_s0[51]}), .O ({new_AGEMA_signal_2040, \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[36], ciphertext_s0[36]}), .I3 ({ciphertext_s1[44], ciphertext_s0[44]}), .I4 ({plaintext_s1[52], plaintext_s0[52]}), .O ({new_AGEMA_signal_2043, \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[37], ciphertext_s0[37]}), .I3 ({ciphertext_s1[45], ciphertext_s0[45]}), .I4 ({plaintext_s1[53], plaintext_s0[53]}), .O ({new_AGEMA_signal_2046, \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[38], ciphertext_s0[38]}), .I3 ({ciphertext_s1[46], ciphertext_s0[46]}), .I4 ({plaintext_s1[54], plaintext_s0[54]}), .O ({new_AGEMA_signal_2049, \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[39], ciphertext_s0[39]}), .I3 ({ciphertext_s1[47], ciphertext_s0[47]}), .I4 ({plaintext_s1[55], plaintext_s0[55]}), .O ({new_AGEMA_signal_2052, \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[56], ciphertext_s0[56]}), .I3 ({ciphertext_s1[32], ciphertext_s0[32]}), .I4 ({plaintext_s1[40], plaintext_s0[40]}), .O ({new_AGEMA_signal_2054, \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[57], ciphertext_s0[57]}), .I3 ({ciphertext_s1[33], ciphertext_s0[33]}), .I4 ({plaintext_s1[41], plaintext_s0[41]}), .O ({new_AGEMA_signal_2056, \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[34], ciphertext_s0[34]}), .I4 ({plaintext_s1[42], plaintext_s0[42]}), .O ({new_AGEMA_signal_2058, \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[59], ciphertext_s0[59]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({plaintext_s1[43], plaintext_s0[43]}), .O ({new_AGEMA_signal_2060, \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[60], ciphertext_s0[60]}), .I3 ({ciphertext_s1[36], ciphertext_s0[36]}), .I4 ({plaintext_s1[44], plaintext_s0[44]}), .O ({new_AGEMA_signal_2062, \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[61], ciphertext_s0[61]}), .I3 ({ciphertext_s1[37], ciphertext_s0[37]}), .I4 ({plaintext_s1[45], plaintext_s0[45]}), .O ({new_AGEMA_signal_2064, \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[62], ciphertext_s0[62]}), .I3 ({ciphertext_s1[38], ciphertext_s0[38]}), .I4 ({plaintext_s1[46], plaintext_s0[46]}), .O ({new_AGEMA_signal_2066, \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[63], ciphertext_s0[63]}), .I3 ({ciphertext_s1[39], ciphertext_s0[39]}), .I4 ({plaintext_s1[47], plaintext_s0[47]}), .O ({new_AGEMA_signal_2068, \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[0], ciphertext_s0[0]}), .I3 ({ciphertext_s1[16], ciphertext_s0[16]}), .I4 ({plaintext_s1[24], plaintext_s0[24]}), .O ({new_AGEMA_signal_2072, \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[1], ciphertext_s0[1]}), .I3 ({ciphertext_s1[17], ciphertext_s0[17]}), .I4 ({plaintext_s1[25], plaintext_s0[25]}), .O ({new_AGEMA_signal_2076, \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[18], ciphertext_s0[18]}), .I4 ({plaintext_s1[26], plaintext_s0[26]}), .O ({new_AGEMA_signal_2080, \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[3], ciphertext_s0[3]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({plaintext_s1[27], plaintext_s0[27]}), .O ({new_AGEMA_signal_2084, \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[4], ciphertext_s0[4]}), .I3 ({ciphertext_s1[20], ciphertext_s0[20]}), .I4 ({plaintext_s1[28], plaintext_s0[28]}), .O ({new_AGEMA_signal_2088, \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[5], ciphertext_s0[5]}), .I3 ({ciphertext_s1[21], ciphertext_s0[21]}), .I4 ({plaintext_s1[29], plaintext_s0[29]}), .O ({new_AGEMA_signal_2092, \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[6], ciphertext_s0[6]}), .I3 ({ciphertext_s1[22], ciphertext_s0[22]}), .I4 ({plaintext_s1[30], plaintext_s0[30]}), .O ({new_AGEMA_signal_2096, \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[7], ciphertext_s0[7]}), .I3 ({ciphertext_s1[23], ciphertext_s0[23]}), .I4 ({plaintext_s1[31], plaintext_s0[31]}), .O ({new_AGEMA_signal_2100, \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[24], ciphertext_s0[24]}), .I3 ({ciphertext_s1[8], ciphertext_s0[8]}), .I4 ({plaintext_s1[16], plaintext_s0[16]}), .O ({new_AGEMA_signal_2103, \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[25], ciphertext_s0[25]}), .I3 ({ciphertext_s1[9], ciphertext_s0[9]}), .I4 ({plaintext_s1[17], plaintext_s0[17]}), .O ({new_AGEMA_signal_2106, \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[10], ciphertext_s0[10]}), .I4 ({plaintext_s1[18], plaintext_s0[18]}), .O ({new_AGEMA_signal_2109, \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[27], ciphertext_s0[27]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({plaintext_s1[19], plaintext_s0[19]}), .O ({new_AGEMA_signal_2112, \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[28], ciphertext_s0[28]}), .I3 ({ciphertext_s1[12], ciphertext_s0[12]}), .I4 ({plaintext_s1[20], plaintext_s0[20]}), .O ({new_AGEMA_signal_2115, \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[29], ciphertext_s0[29]}), .I3 ({ciphertext_s1[13], ciphertext_s0[13]}), .I4 ({plaintext_s1[21], plaintext_s0[21]}), .O ({new_AGEMA_signal_2118, \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[30], ciphertext_s0[30]}), .I3 ({ciphertext_s1[14], ciphertext_s0[14]}), .I4 ({plaintext_s1[22], plaintext_s0[22]}), .O ({new_AGEMA_signal_2121, \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[31], ciphertext_s0[31]}), .I3 ({ciphertext_s1[15], ciphertext_s0[15]}), .I4 ({plaintext_s1[23], plaintext_s0[23]}), .O ({new_AGEMA_signal_2124, \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[16], ciphertext_s0[16]}), .I3 ({ciphertext_s1[0], ciphertext_s0[0]}), .I4 ({plaintext_s1[8], plaintext_s0[8]}), .O ({new_AGEMA_signal_2126, \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[17], ciphertext_s0[17]}), .I3 ({ciphertext_s1[1], ciphertext_s0[1]}), .I4 ({plaintext_s1[9], plaintext_s0[9]}), .O ({new_AGEMA_signal_2128, \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[2], ciphertext_s0[2]}), .I4 ({plaintext_s1[10], plaintext_s0[10]}), .O ({new_AGEMA_signal_2130, \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[19], ciphertext_s0[19]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({plaintext_s1[11], plaintext_s0[11]}), .O ({new_AGEMA_signal_2132, \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[20], ciphertext_s0[20]}), .I3 ({ciphertext_s1[4], ciphertext_s0[4]}), .I4 ({plaintext_s1[12], plaintext_s0[12]}), .O ({new_AGEMA_signal_2134, \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[21], ciphertext_s0[21]}), .I3 ({ciphertext_s1[5], ciphertext_s0[5]}), .I4 ({plaintext_s1[13], plaintext_s0[13]}), .O ({new_AGEMA_signal_2136, \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[22], ciphertext_s0[22]}), .I3 ({ciphertext_s1[6], ciphertext_s0[6]}), .I4 ({plaintext_s1[14], plaintext_s0[14]}), .O ({new_AGEMA_signal_2138, \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[23], ciphertext_s0[23]}), .I3 ({ciphertext_s1[7], ciphertext_s0[7]}), .I4 ({plaintext_s1[15], plaintext_s0[15]}), .O ({new_AGEMA_signal_2140, \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }), .I3 ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }), .I4 ({key_s1[112], key_s0[112]}), .O ({new_AGEMA_signal_1528, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }), .I3 ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }), .I4 ({key_s1[113], key_s0[113]}), .O ({new_AGEMA_signal_1532, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }), .I3 ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }), .I4 ({key_s1[114], key_s0[114]}), .O ({new_AGEMA_signal_1536, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }), .I3 ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }), .I4 ({key_s1[115], key_s0[115]}), .O ({new_AGEMA_signal_1540, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }), .I3 ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }), .I4 ({key_s1[116], key_s0[116]}), .O ({new_AGEMA_signal_1544, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }), .I3 ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }), .I4 ({key_s1[117], key_s0[117]}), .O ({new_AGEMA_signal_1548, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }), .I3 ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }), .I4 ({key_s1[118], key_s0[118]}), .O ({new_AGEMA_signal_1552, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }), .I3 ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }), .I4 ({key_s1[119], key_s0[119]}), .O ({new_AGEMA_signal_1556, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }), .I3 ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }), .I4 ({key_s1[104], key_s0[104]}), .O ({new_AGEMA_signal_1560, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }), .I3 ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }), .I4 ({key_s1[105], key_s0[105]}), .O ({new_AGEMA_signal_1564, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }), .I3 ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }), .I4 ({key_s1[106], key_s0[106]}), .O ({new_AGEMA_signal_1568, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }), .I3 ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }), .I4 ({key_s1[107], key_s0[107]}), .O ({new_AGEMA_signal_1572, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }), .I3 ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }), .I4 ({key_s1[108], key_s0[108]}), .O ({new_AGEMA_signal_1576, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }), .I3 ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }), .I4 ({key_s1[109], key_s0[109]}), .O ({new_AGEMA_signal_1580, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }), .I3 ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }), .I4 ({key_s1[110], key_s0[110]}), .O ({new_AGEMA_signal_1584, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }), .I3 ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }), .I4 ({key_s1[111], key_s0[111]}), .O ({new_AGEMA_signal_1588, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I3 ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }), .I4 ({key_s1[96], key_s0[96]}), .O ({new_AGEMA_signal_1591, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I3 ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }), .I4 ({key_s1[97], key_s0[97]}), .O ({new_AGEMA_signal_1594, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I3 ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }), .I4 ({key_s1[98], key_s0[98]}), .O ({new_AGEMA_signal_1597, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I3 ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }), .I4 ({key_s1[99], key_s0[99]}), .O ({new_AGEMA_signal_1600, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I3 ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }), .I4 ({key_s1[100], key_s0[100]}), .O ({new_AGEMA_signal_1603, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I3 ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }), .I4 ({key_s1[101], key_s0[101]}), .O ({new_AGEMA_signal_1606, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I3 ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }), .I4 ({key_s1[102], key_s0[102]}), .O ({new_AGEMA_signal_1609, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I3 ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }), .I4 ({key_s1[103], key_s0[103]}), .O ({new_AGEMA_signal_1612, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }), .I3 ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }), .I4 ({key_s1[88], key_s0[88]}), .O ({new_AGEMA_signal_1615, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }), .I3 ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }), .I4 ({key_s1[89], key_s0[89]}), .O ({new_AGEMA_signal_1618, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }), .I3 ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }), .I4 ({key_s1[90], key_s0[90]}), .O ({new_AGEMA_signal_1621, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }), .I3 ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }), .I4 ({key_s1[91], key_s0[91]}), .O ({new_AGEMA_signal_1624, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }), .I3 ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }), .I4 ({key_s1[92], key_s0[92]}), .O ({new_AGEMA_signal_1627, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }), .I3 ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }), .I4 ({key_s1[93], key_s0[93]}), .O ({new_AGEMA_signal_1630, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }), .I3 ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }), .I4 ({key_s1[94], key_s0[94]}), .O ({new_AGEMA_signal_1633, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }), .I3 ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }), .I4 ({key_s1[95], key_s0[95]}), .O ({new_AGEMA_signal_1636, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }), .I3 ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }), .I4 ({key_s1[80], key_s0[80]}), .O ({new_AGEMA_signal_1639, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }), .I3 ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }), .I4 ({key_s1[81], key_s0[81]}), .O ({new_AGEMA_signal_1642, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }), .I3 ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }), .I4 ({key_s1[82], key_s0[82]}), .O ({new_AGEMA_signal_1645, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }), .I3 ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }), .I4 ({key_s1[83], key_s0[83]}), .O ({new_AGEMA_signal_1648, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }), .I3 ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }), .I4 ({key_s1[84], key_s0[84]}), .O ({new_AGEMA_signal_1651, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }), .I3 ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }), .I4 ({key_s1[85], key_s0[85]}), .O ({new_AGEMA_signal_1654, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }), .I3 ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }), .I4 ({key_s1[86], key_s0[86]}), .O ({new_AGEMA_signal_1657, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }), .I3 ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }), .I4 ({key_s1[87], key_s0[87]}), .O ({new_AGEMA_signal_1660, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }), .I3 ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }), .I4 ({key_s1[72], key_s0[72]}), .O ({new_AGEMA_signal_1663, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }), .I3 ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }), .I4 ({key_s1[73], key_s0[73]}), .O ({new_AGEMA_signal_1666, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }), .I3 ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }), .I4 ({key_s1[74], key_s0[74]}), .O ({new_AGEMA_signal_1669, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }), .I3 ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }), .I4 ({key_s1[75], key_s0[75]}), .O ({new_AGEMA_signal_1672, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }), .I3 ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }), .I4 ({key_s1[76], key_s0[76]}), .O ({new_AGEMA_signal_1675, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }), .I3 ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }), .I4 ({key_s1[77], key_s0[77]}), .O ({new_AGEMA_signal_1678, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }), .I3 ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }), .I4 ({key_s1[78], key_s0[78]}), .O ({new_AGEMA_signal_1681, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }), .I3 ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }), .I4 ({key_s1[79], key_s0[79]}), .O ({new_AGEMA_signal_1684, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }), .I3 ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }), .I4 ({key_s1[64], key_s0[64]}), .O ({new_AGEMA_signal_1687, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }), .I3 ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }), .I4 ({key_s1[65], key_s0[65]}), .O ({new_AGEMA_signal_1690, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }), .I3 ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }), .I4 ({key_s1[66], key_s0[66]}), .O ({new_AGEMA_signal_1693, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }), .I3 ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }), .I4 ({key_s1[67], key_s0[67]}), .O ({new_AGEMA_signal_1696, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }), .I3 ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }), .I4 ({key_s1[68], key_s0[68]}), .O ({new_AGEMA_signal_1699, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }), .I3 ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }), .I4 ({key_s1[69], key_s0[69]}), .O ({new_AGEMA_signal_1702, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }), .I3 ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }), .I4 ({key_s1[70], key_s0[70]}), .O ({new_AGEMA_signal_1705, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }), .I3 ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }), .I4 ({key_s1[71], key_s0[71]}), .O ({new_AGEMA_signal_1708, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }), .I3 ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }), .I4 ({key_s1[56], key_s0[56]}), .O ({new_AGEMA_signal_1711, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }), .I3 ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }), .I4 ({key_s1[57], key_s0[57]}), .O ({new_AGEMA_signal_1714, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }), .I3 ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }), .I4 ({key_s1[58], key_s0[58]}), .O ({new_AGEMA_signal_1717, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }), .I3 ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }), .I4 ({key_s1[59], key_s0[59]}), .O ({new_AGEMA_signal_1720, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }), .I3 ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }), .I4 ({key_s1[60], key_s0[60]}), .O ({new_AGEMA_signal_1723, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }), .I3 ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }), .I4 ({key_s1[61], key_s0[61]}), .O ({new_AGEMA_signal_1726, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }), .I3 ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }), .I4 ({key_s1[62], key_s0[62]}), .O ({new_AGEMA_signal_1729, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }), .I3 ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }), .I4 ({key_s1[63], key_s0[63]}), .O ({new_AGEMA_signal_1732, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }), .I3 ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }), .I4 ({key_s1[48], key_s0[48]}), .O ({new_AGEMA_signal_1735, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }), .I3 ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }), .I4 ({key_s1[49], key_s0[49]}), .O ({new_AGEMA_signal_1738, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }), .I3 ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }), .I4 ({key_s1[50], key_s0[50]}), .O ({new_AGEMA_signal_1741, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }), .I3 ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }), .I4 ({key_s1[51], key_s0[51]}), .O ({new_AGEMA_signal_1744, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }), .I3 ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }), .I4 ({key_s1[52], key_s0[52]}), .O ({new_AGEMA_signal_1747, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }), .I3 ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }), .I4 ({key_s1[53], key_s0[53]}), .O ({new_AGEMA_signal_1750, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }), .I3 ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }), .I4 ({key_s1[54], key_s0[54]}), .O ({new_AGEMA_signal_1753, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }), .I3 ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }), .I4 ({key_s1[55], key_s0[55]}), .O ({new_AGEMA_signal_1756, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }), .I3 ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }), .I4 ({key_s1[40], key_s0[40]}), .O ({new_AGEMA_signal_1759, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }), .I3 ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }), .I4 ({key_s1[41], key_s0[41]}), .O ({new_AGEMA_signal_1762, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }), .I3 ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }), .I4 ({key_s1[42], key_s0[42]}), .O ({new_AGEMA_signal_1765, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }), .I3 ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }), .I4 ({key_s1[43], key_s0[43]}), .O ({new_AGEMA_signal_1768, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }), .I3 ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }), .I4 ({key_s1[44], key_s0[44]}), .O ({new_AGEMA_signal_1771, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }), .I3 ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }), .I4 ({key_s1[45], key_s0[45]}), .O ({new_AGEMA_signal_1774, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }), .I3 ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }), .I4 ({key_s1[46], key_s0[46]}), .O ({new_AGEMA_signal_1777, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }), .I3 ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }), .I4 ({key_s1[47], key_s0[47]}), .O ({new_AGEMA_signal_1780, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }), .I3 ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }), .I4 ({key_s1[32], key_s0[32]}), .O ({new_AGEMA_signal_1783, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }), .I3 ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }), .I4 ({key_s1[33], key_s0[33]}), .O ({new_AGEMA_signal_1786, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }), .I3 ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }), .I4 ({key_s1[34], key_s0[34]}), .O ({new_AGEMA_signal_1789, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }), .I3 ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }), .I4 ({key_s1[35], key_s0[35]}), .O ({new_AGEMA_signal_1792, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }), .I3 ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }), .I4 ({key_s1[36], key_s0[36]}), .O ({new_AGEMA_signal_1795, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }), .I3 ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }), .I4 ({key_s1[37], key_s0[37]}), .O ({new_AGEMA_signal_1798, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }), .I3 ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }), .I4 ({key_s1[38], key_s0[38]}), .O ({new_AGEMA_signal_1801, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }), .I3 ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }), .I4 ({key_s1[39], key_s0[39]}), .O ({new_AGEMA_signal_1804, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }), .I3 ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }), .I4 ({key_s1[16], key_s0[16]}), .O ({new_AGEMA_signal_1807, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }), .I3 ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }), .I4 ({key_s1[17], key_s0[17]}), .O ({new_AGEMA_signal_1810, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }), .I3 ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }), .I4 ({key_s1[18], key_s0[18]}), .O ({new_AGEMA_signal_1813, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }), .I3 ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }), .I4 ({key_s1[19], key_s0[19]}), .O ({new_AGEMA_signal_1816, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }), .I3 ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }), .I4 ({key_s1[20], key_s0[20]}), .O ({new_AGEMA_signal_1819, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }), .I3 ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }), .I4 ({key_s1[21], key_s0[21]}), .O ({new_AGEMA_signal_1822, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }), .I3 ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }), .I4 ({key_s1[22], key_s0[22]}), .O ({new_AGEMA_signal_1825, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }), .I3 ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }), .I4 ({key_s1[23], key_s0[23]}), .O ({new_AGEMA_signal_1828, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }), .I3 ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }), .I4 ({key_s1[8], key_s0[8]}), .O ({new_AGEMA_signal_1830, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }), .I3 ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }), .I4 ({key_s1[9], key_s0[9]}), .O ({new_AGEMA_signal_1832, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }), .I3 ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }), .I4 ({key_s1[10], key_s0[10]}), .O ({new_AGEMA_signal_1834, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }), .I3 ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }), .I4 ({key_s1[11], key_s0[11]}), .O ({new_AGEMA_signal_1836, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }), .I3 ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }), .I4 ({key_s1[12], key_s0[12]}), .O ({new_AGEMA_signal_1838, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }), .I3 ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }), .I4 ({key_s1[13], key_s0[13]}), .O ({new_AGEMA_signal_1840, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }), .I3 ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }), .I4 ({key_s1[14], key_s0[14]}), .O ({new_AGEMA_signal_1842, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }), .I3 ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }), .I4 ({key_s1[15], key_s0[15]}), .O ({new_AGEMA_signal_1844, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }), .I3 ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }), .I4 ({key_s1[0], key_s0[0]}), .O ({new_AGEMA_signal_1846, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }), .I3 ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }), .I4 ({key_s1[1], key_s0[1]}), .O ({new_AGEMA_signal_1848, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }), .I3 ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }), .I4 ({key_s1[2], key_s0[2]}), .O ({new_AGEMA_signal_1850, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }), .I3 ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }), .I4 ({key_s1[3], key_s0[3]}), .O ({new_AGEMA_signal_1852, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }), .I3 ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }), .I4 ({key_s1[4], key_s0[4]}), .O ({new_AGEMA_signal_1854, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }), .I3 ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }), .I4 ({key_s1[5], key_s0[5]}), .O ({new_AGEMA_signal_1856, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }), .I3 ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }), .I4 ({key_s1[6], key_s0[6]}), .O ({new_AGEMA_signal_1858, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/CSselMC_835 }), .I2 ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }), .I3 ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }), .I4 ({key_s1[7], key_s0[7]}), .O ({new_AGEMA_signal_1860, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[96], ciphertext_s0[96]}), .I3 ({new_AGEMA_signal_1901, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_897 }), .I4 ({plaintext_s1[96], plaintext_s0[96]}), .O ({new_AGEMA_signal_2166, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[97], ciphertext_s0[97]}), .I3 ({new_AGEMA_signal_1916, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[97], plaintext_s0[97]}), .O ({new_AGEMA_signal_2168, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({new_AGEMA_signal_1902, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_900 }), .I4 ({plaintext_s1[98], plaintext_s0[98]}), .O ({new_AGEMA_signal_2170, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[99], ciphertext_s0[99]}), .I3 ({new_AGEMA_signal_1917, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[99], plaintext_s0[99]}), .O ({new_AGEMA_signal_2172, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[100], ciphertext_s0[100]}), .I3 ({new_AGEMA_signal_1918, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[100], plaintext_s0[100]}), .O ({new_AGEMA_signal_2174, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[101], ciphertext_s0[101]}), .I3 ({new_AGEMA_signal_1903, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_904 }), .I4 ({plaintext_s1[101], plaintext_s0[101]}), .O ({new_AGEMA_signal_2176, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[102], ciphertext_s0[102]}), .I3 ({new_AGEMA_signal_1904, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_906 }), .I4 ({plaintext_s1[102], plaintext_s0[102]}), .O ({new_AGEMA_signal_2178, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[103], ciphertext_s0[103]}), .I3 ({new_AGEMA_signal_1905, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_908 }), .I4 ({plaintext_s1[103], plaintext_s0[103]}), .O ({new_AGEMA_signal_2180, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[88], ciphertext_s0[88]}), .I3 ({new_AGEMA_signal_1906, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_910 }), .I4 ({plaintext_s1[64], plaintext_s0[64]}), .O ({new_AGEMA_signal_2182, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[89], ciphertext_s0[89]}), .I3 ({new_AGEMA_signal_1919, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[65], plaintext_s0[65]}), .O ({new_AGEMA_signal_2184, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({new_AGEMA_signal_1907, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_913 }), .I4 ({plaintext_s1[66], plaintext_s0[66]}), .O ({new_AGEMA_signal_2186, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[91], ciphertext_s0[91]}), .I3 ({new_AGEMA_signal_1920, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[67], plaintext_s0[67]}), .O ({new_AGEMA_signal_2188, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[92], ciphertext_s0[92]}), .I3 ({new_AGEMA_signal_1921, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[68], plaintext_s0[68]}), .O ({new_AGEMA_signal_2190, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[93], ciphertext_s0[93]}), .I3 ({new_AGEMA_signal_1908, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_917 }), .I4 ({plaintext_s1[69], plaintext_s0[69]}), .O ({new_AGEMA_signal_2192, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[94], ciphertext_s0[94]}), .I3 ({new_AGEMA_signal_1909, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_919 }), .I4 ({plaintext_s1[70], plaintext_s0[70]}), .O ({new_AGEMA_signal_2194, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[95], ciphertext_s0[95]}), .I3 ({new_AGEMA_signal_1910, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_921 }), .I4 ({plaintext_s1[71], plaintext_s0[71]}), .O ({new_AGEMA_signal_2196, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[48], ciphertext_s0[48]}), .I3 ({new_AGEMA_signal_1911, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11_923 }), .I4 ({plaintext_s1[32], plaintext_s0[32]}), .O ({new_AGEMA_signal_2198, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[49], ciphertext_s0[49]}), .I3 ({new_AGEMA_signal_1922, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[33], plaintext_s0[33]}), .O ({new_AGEMA_signal_2200, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({new_AGEMA_signal_1912, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11_926 }), .I4 ({plaintext_s1[34], plaintext_s0[34]}), .O ({new_AGEMA_signal_2202, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[51], ciphertext_s0[51]}), .I3 ({new_AGEMA_signal_1923, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[35], plaintext_s0[35]}), .O ({new_AGEMA_signal_2204, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q14 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[52], ciphertext_s0[52]}), .I3 ({new_AGEMA_signal_1924, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q12 }), .I4 ({plaintext_s1[36], plaintext_s0[36]}), .O ({new_AGEMA_signal_2206, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[53], ciphertext_s0[53]}), .I3 ({new_AGEMA_signal_1913, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11_930 }), .I4 ({plaintext_s1[37], plaintext_s0[37]}), .O ({new_AGEMA_signal_2208, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[54], ciphertext_s0[54]}), .I3 ({new_AGEMA_signal_1914, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11_932 }), .I4 ({plaintext_s1[38], plaintext_s0[38]}), .O ({new_AGEMA_signal_2210, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hF7D5A280 ) , .MASK ( 5'b00011 ), .INIT2 ( 32'hF7D5A280 ) ) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q13 ( .I0 ({1'b0, nReset_407}), .I1 ({1'b0, \ctrl/finalStep1 }), .I2 ({ciphertext_s1[55], ciphertext_s0[55]}), .I3 ({new_AGEMA_signal_1915, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11_934 }), .I4 ({plaintext_s1[39], plaintext_s0[39]}), .O ({new_AGEMA_signal_2212, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6 #( .INIT ( 64'h0000000000000002 ) ) \ctrl/selSR1 ( .I0 (nReset_407), .I1 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .I2 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I3 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I4 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I5 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .O (selSR) ) ;
    LUT5 #( .INIT ( 32'hFFFF8880 ) ) \ctrl/CSselMC_rstpot ( .I0 (nReset_407), .I1 (\ctrl/CSselMC_835 ), .I2 (\ctrl/seq4/GEN[0].SFF/Q_836 ), .I3 (\ctrl/seq4/GEN[1].SFF/Q_837 ), .I4 (\ctrl/finalStep1 ), .O (\ctrl/CSselMC_rstpot_1330 ) ) ;
    LUT6 #( .INIT ( 64'hFFFFFFFFFFFEFFFF ) ) enKS1 ( .I0 (\ctrl/seq6/GEN[2].SFF/Q_839 ), .I1 (\ctrl/seq6/GEN[4].SFF/Q_842 ), .I2 (\ctrl/seq6/GEN[3].SFF/Q_840 ), .I3 (\ctrl/seq6/GEN[1].SFF/Q_838 ), .I4 (nReset_407), .I5 (\ctrl/seq6/GEN[0].SFF/Q_841 ), .O (enKS) ) ;
    INV \ctrl/nReset_inv1_INV_0 ( .I (nReset_407), .O (\calcRCon/nReset_inv ) ) ;
    INV nReset_rstpot1_INV_0 ( .I (start), .O (nReset_rstpot) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (start), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \Inst_bSbox/b7_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[0]), .O ({new_AGEMA_signal_1861, \Inst_bSbox/b7 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \Inst_bSbox/b7_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[1]), .O ({new_AGEMA_signal_1862, \Inst_bSbox/b7 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \Inst_bSbox/b7_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[2]), .O ({new_AGEMA_signal_1863, \Inst_bSbox/b7 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \Inst_bSbox/b7_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[3]), .O ({new_AGEMA_signal_1864, \Inst_bSbox/b7 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \Inst_bSbox/b6_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[4]), .O ({new_AGEMA_signal_1865, \Inst_bSbox/b6 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \Inst_bSbox/b6_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[5]), .O ({new_AGEMA_signal_1866, \Inst_bSbox/b6 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \Inst_bSbox/b6_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[6]), .O ({new_AGEMA_signal_1867, \Inst_bSbox/b6 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \Inst_bSbox/b6_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[7]), .O ({new_AGEMA_signal_1868, \Inst_bSbox/b6 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \Inst_bSbox/b5_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[8]), .O ({new_AGEMA_signal_1869, \Inst_bSbox/b5 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \Inst_bSbox/b5_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[9]), .O ({new_AGEMA_signal_1870, \Inst_bSbox/b5 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \Inst_bSbox/b5_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[10]), .O ({new_AGEMA_signal_1871, \Inst_bSbox/b5 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \Inst_bSbox/b5_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[11]), .O ({new_AGEMA_signal_1872, \Inst_bSbox/b5 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \Inst_bSbox/b4_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[12]), .O ({new_AGEMA_signal_1873, \Inst_bSbox/b4 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \Inst_bSbox/b4_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[13]), .O ({new_AGEMA_signal_1874, \Inst_bSbox/b4 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \Inst_bSbox/b4_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[14]), .O ({new_AGEMA_signal_1875, \Inst_bSbox/b4 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \Inst_bSbox/b4_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[15]), .O ({new_AGEMA_signal_1876, \Inst_bSbox/b4 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \Inst_bSbox/b3_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[16]), .O ({new_AGEMA_signal_1877, \Inst_bSbox/b3 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \Inst_bSbox/b3_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[17]), .O ({new_AGEMA_signal_1878, \Inst_bSbox/b3 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \Inst_bSbox/b3_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[18]), .O ({new_AGEMA_signal_1879, \Inst_bSbox/b3 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \Inst_bSbox/b3_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[19]), .O ({new_AGEMA_signal_1880, \Inst_bSbox/b3 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \Inst_bSbox/b2_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[20]), .O ({new_AGEMA_signal_1881, \Inst_bSbox/b2 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \Inst_bSbox/b2_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[21]), .O ({new_AGEMA_signal_1882, \Inst_bSbox/b2 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \Inst_bSbox/b2_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[22]), .O ({new_AGEMA_signal_1883, \Inst_bSbox/b2 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \Inst_bSbox/b2_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[23]), .O ({new_AGEMA_signal_1884, \Inst_bSbox/b2 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \Inst_bSbox/b1_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[24]), .O ({new_AGEMA_signal_1885, \Inst_bSbox/b1 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \Inst_bSbox/b1_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[25]), .O ({new_AGEMA_signal_1886, \Inst_bSbox/b1 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \Inst_bSbox/b1_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[26]), .O ({new_AGEMA_signal_1887, \Inst_bSbox/b1 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \Inst_bSbox/b1_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[27]), .O ({new_AGEMA_signal_1888, \Inst_bSbox/b1 [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \Inst_bSbox/b0_3 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[28]), .O ({new_AGEMA_signal_1889, \Inst_bSbox/b0 [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \Inst_bSbox/b0_2 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[29]), .O ({new_AGEMA_signal_1890, \Inst_bSbox/b0 [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \Inst_bSbox/b0_1 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[30]), .O ({new_AGEMA_signal_1891, \Inst_bSbox/b0 [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \Inst_bSbox/b0_0 ( .I0 ({new_AGEMA_signal_1434, SboxIn[0]}), .I1 ({new_AGEMA_signal_1432, SboxIn[1]}), .I2 ({new_AGEMA_signal_1430, SboxIn[2]}), .I3 ({new_AGEMA_signal_1428, SboxIn[3]}), .I4 ({new_AGEMA_signal_1426, SboxIn[4]}), .I5 ({new_AGEMA_signal_1424, SboxIn[5]}), .clk (clk), .r (Fresh[31]), .O ({new_AGEMA_signal_1892, \Inst_bSbox/b0 [0]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[7].Inst1 ( .I0 ({new_AGEMA_signal_1900, StateInMC[7]}), .I1 ({new_AGEMA_signal_2157, SboxOut[7]}), .I2 ({new_AGEMA_signal_1351, StateOutXORroundKey[7]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2213, \stateArray/input_MC [7]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[6].Inst1 ( .I0 ({new_AGEMA_signal_1899, StateInMC[6]}), .I1 ({new_AGEMA_signal_2158, SboxOut[6]}), .I2 ({new_AGEMA_signal_1354, StateOutXORroundKey[6]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2214, \stateArray/input_MC [6]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[5].Inst1 ( .I0 ({new_AGEMA_signal_1898, StateInMC[5]}), .I1 ({new_AGEMA_signal_2159, SboxOut[5]}), .I2 ({new_AGEMA_signal_1357, StateOutXORroundKey[5]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2215, \stateArray/input_MC [5]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[4].Inst1 ( .I0 ({new_AGEMA_signal_1897, StateInMC[4]}), .I1 ({new_AGEMA_signal_2160, SboxOut[4]}), .I2 ({new_AGEMA_signal_1360, StateOutXORroundKey[4]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2216, \stateArray/input_MC [4]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[3].Inst1 ( .I0 ({new_AGEMA_signal_1896, StateInMC[3]}), .I1 ({new_AGEMA_signal_2161, SboxOut[3]}), .I2 ({new_AGEMA_signal_1363, StateOutXORroundKey[3]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2217, \stateArray/input_MC [3]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[2].Inst1 ( .I0 ({new_AGEMA_signal_1895, StateInMC[2]}), .I1 ({new_AGEMA_signal_2162, SboxOut[2]}), .I2 ({new_AGEMA_signal_1366, StateOutXORroundKey[2]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2218, \stateArray/input_MC [2]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[1].Inst1 ( .I0 ({new_AGEMA_signal_1894, StateInMC[1]}), .I1 ({new_AGEMA_signal_2163, SboxOut[1]}), .I2 ({new_AGEMA_signal_1369, StateOutXORroundKey[1]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2219, \stateArray/input_MC [1]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hAAAAF0CC ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hAAAAF0CC ) ) \stateArray/gen33ser[0].Inst1 ( .I0 ({new_AGEMA_signal_1893, StateInMC[0]}), .I1 ({new_AGEMA_signal_2164, SboxOut[0]}), .I2 ({new_AGEMA_signal_1372, StateOutXORroundKey[0]}), .I3 ({1'b0, intFinal}), .I4 ({1'b0, selMC}), .O ({new_AGEMA_signal_2220, \stateArray/input_MC [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b7_4 ( .I0 ({new_AGEMA_signal_1864, \Inst_bSbox/b7 [0]}), .I1 ({new_AGEMA_signal_1863, \Inst_bSbox/b7 [1]}), .I2 ({new_AGEMA_signal_1862, \Inst_bSbox/b7 [2]}), .I3 ({new_AGEMA_signal_1861, \Inst_bSbox/b7 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[32]), .O ({new_AGEMA_signal_2157, SboxOut[7]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b6_4 ( .I0 ({new_AGEMA_signal_1868, \Inst_bSbox/b6 [0]}), .I1 ({new_AGEMA_signal_1867, \Inst_bSbox/b6 [1]}), .I2 ({new_AGEMA_signal_1866, \Inst_bSbox/b6 [2]}), .I3 ({new_AGEMA_signal_1865, \Inst_bSbox/b6 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[33]), .O ({new_AGEMA_signal_2158, SboxOut[6]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b5_4 ( .I0 ({new_AGEMA_signal_1872, \Inst_bSbox/b5 [0]}), .I1 ({new_AGEMA_signal_1871, \Inst_bSbox/b5 [1]}), .I2 ({new_AGEMA_signal_1870, \Inst_bSbox/b5 [2]}), .I3 ({new_AGEMA_signal_1869, \Inst_bSbox/b5 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[34]), .O ({new_AGEMA_signal_2159, SboxOut[5]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b4_4 ( .I0 ({new_AGEMA_signal_1876, \Inst_bSbox/b4 [0]}), .I1 ({new_AGEMA_signal_1875, \Inst_bSbox/b4 [1]}), .I2 ({new_AGEMA_signal_1874, \Inst_bSbox/b4 [2]}), .I3 ({new_AGEMA_signal_1873, \Inst_bSbox/b4 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[35]), .O ({new_AGEMA_signal_2160, SboxOut[4]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b3_4 ( .I0 ({new_AGEMA_signal_1880, \Inst_bSbox/b3 [0]}), .I1 ({new_AGEMA_signal_1879, \Inst_bSbox/b3 [1]}), .I2 ({new_AGEMA_signal_1878, \Inst_bSbox/b3 [2]}), .I3 ({new_AGEMA_signal_1877, \Inst_bSbox/b3 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[36]), .O ({new_AGEMA_signal_2161, SboxOut[3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b2_4 ( .I0 ({new_AGEMA_signal_1884, \Inst_bSbox/b2 [0]}), .I1 ({new_AGEMA_signal_1883, \Inst_bSbox/b2 [1]}), .I2 ({new_AGEMA_signal_1882, \Inst_bSbox/b2 [2]}), .I3 ({new_AGEMA_signal_1881, \Inst_bSbox/b2 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[37]), .O ({new_AGEMA_signal_2162, SboxOut[2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b1_4 ( .I0 ({new_AGEMA_signal_1888, \Inst_bSbox/b1 [0]}), .I1 ({new_AGEMA_signal_1887, \Inst_bSbox/b1 [1]}), .I2 ({new_AGEMA_signal_1886, \Inst_bSbox/b1 [2]}), .I3 ({new_AGEMA_signal_1885, \Inst_bSbox/b1 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[38]), .O ({new_AGEMA_signal_2163, SboxOut[1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \Inst_bSbox/b0_4 ( .I0 ({new_AGEMA_signal_1892, \Inst_bSbox/b0 [0]}), .I1 ({new_AGEMA_signal_1891, \Inst_bSbox/b0 [1]}), .I2 ({new_AGEMA_signal_1890, \Inst_bSbox/b0 [2]}), .I3 ({new_AGEMA_signal_1889, \Inst_bSbox/b0 [3]}), .I4 ({new_AGEMA_signal_1438, SboxIn[6]}), .I5 ({new_AGEMA_signal_1436, SboxIn[7]}), .clk (clk), .r (Fresh[39]), .O ({new_AGEMA_signal_2164, SboxOut[0]}) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[0], plaintext_s0[0]}), .I1 ({ciphertext_s1[8], ciphertext_s0[8]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2220, \stateArray/input_MC [0]}), .O ({new_AGEMA_signal_2246, \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[1], plaintext_s0[1]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2219, \stateArray/input_MC [1]}), .O ({new_AGEMA_signal_2248, \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[2], plaintext_s0[2]}), .I1 ({ciphertext_s1[10], ciphertext_s0[10]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2218, \stateArray/input_MC [2]}), .O ({new_AGEMA_signal_2250, \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[3], plaintext_s0[3]}), .I1 ({ciphertext_s1[11], ciphertext_s0[11]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2217, \stateArray/input_MC [3]}), .O ({new_AGEMA_signal_2252, \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[4], plaintext_s0[4]}), .I1 ({ciphertext_s1[12], ciphertext_s0[12]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2216, \stateArray/input_MC [4]}), .O ({new_AGEMA_signal_2254, \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[5], plaintext_s0[5]}), .I1 ({ciphertext_s1[13], ciphertext_s0[13]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2215, \stateArray/input_MC [5]}), .O ({new_AGEMA_signal_2256, \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[6], plaintext_s0[6]}), .I1 ({ciphertext_s1[14], ciphertext_s0[14]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2214, \stateArray/input_MC [6]}), .O ({new_AGEMA_signal_2258, \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hCAFACA0A ) , .MASK ( 5'b01100 ), .INIT2 ( 32'hCAFACA0A ) ) \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q11 ( .I0 ({plaintext_s1[7], plaintext_s0[7]}), .I1 ({ciphertext_s1[15], ciphertext_s0[15]}), .I2 ({1'b0, nReset_407}), .I3 ({1'b0, \ctrl/finalStep1 }), .I4 ({new_AGEMA_signal_2213, \stateArray/input_MC [7]}), .O ({new_AGEMA_signal_2260, \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[24], key_s0[24]}), .I1 ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1415, N18}), .I5 ({new_AGEMA_signal_2164, SboxOut[0]}), .O ({new_AGEMA_signal_2222, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[25], key_s0[25]}), .I1 ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1416, N20}), .I5 ({new_AGEMA_signal_2163, SboxOut[1]}), .O ({new_AGEMA_signal_2224, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[26], key_s0[26]}), .I1 ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1417, N22}), .I5 ({new_AGEMA_signal_2162, SboxOut[2]}), .O ({new_AGEMA_signal_2226, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[27], key_s0[27]}), .I1 ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1418, N24}), .I5 ({new_AGEMA_signal_2161, SboxOut[3]}), .O ({new_AGEMA_signal_2228, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[28], key_s0[28]}), .I1 ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1419, N26}), .I5 ({new_AGEMA_signal_2160, SboxOut[4]}), .O ({new_AGEMA_signal_2230, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[29], key_s0[29]}), .I1 ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1420, N28}), .I5 ({new_AGEMA_signal_2159, SboxOut[5]}), .O ({new_AGEMA_signal_2232, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[30], key_s0[30]}), .I1 ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1421, N30}), .I5 ({new_AGEMA_signal_2158, SboxOut[6]}), .O ({new_AGEMA_signal_2234, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFCAA0CAA0CAAFCAA ) , .MASK ( 6'b001100 ), .INIT2 ( 64'h0CAAFCAAFCAA0CAA ) ) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/MUXInst/Mmux_Q1 ( .I0 ({key_s1[31], key_s0[31]}), .I1 ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }), .I2 ({1'b0, \ctrl/CSselMC_835 }), .I3 ({1'b0, nReset_407}), .I4 ({new_AGEMA_signal_1422, N32}), .I5 ({new_AGEMA_signal_2157, SboxOut[7]}), .O ({new_AGEMA_signal_2236, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }) ) ;

    /* register cells */
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1927, \stateArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1930, \stateArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1933, \stateArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1936, \stateArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1939, \stateArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1942, \stateArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1945, \stateArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1948, \stateArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1951, \stateArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1954, \stateArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1957, \stateArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1960, \stateArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1963, \stateArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1966, \stateArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1969, \stateArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1972, \stateArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1975, \stateArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1978, \stateArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1981, \stateArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1984, \stateArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1987, \stateArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1990, \stateArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1993, \stateArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1996, \stateArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2166, \stateArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2168, \stateArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2170, \stateArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2172, \stateArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2174, \stateArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2176, \stateArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2178, \stateArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2180, \stateArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1455, \stateArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1458, \stateArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1461, \stateArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1464, \stateArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1467, \stateArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1470, \stateArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1473, \stateArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1476, \stateArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1479, \stateArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1482, \stateArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1485, \stateArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1488, \stateArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1491, \stateArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1494, \stateArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1497, \stateArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1500, \stateArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1503, \stateArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1506, \stateArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1509, \stateArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1512, \stateArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1515, \stateArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1518, \stateArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1521, \stateArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1524, \stateArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2182, \stateArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2184, \stateArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2186, \stateArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2188, \stateArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2190, \stateArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2192, \stateArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2194, \stateArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2196, \stateArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2000, \stateArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2004, \stateArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2008, \stateArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2012, \stateArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2016, \stateArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2020, \stateArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2024, \stateArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2028, \stateArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2031, \stateArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2034, \stateArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2037, \stateArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2040, \stateArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2043, \stateArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2046, \stateArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2049, \stateArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2052, \stateArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2054, \stateArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2056, \stateArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2058, \stateArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2060, \stateArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2062, \stateArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2064, \stateArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2066, \stateArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2068, \stateArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2198, \stateArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2200, \stateArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2202, \stateArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2204, \stateArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2206, \stateArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2208, \stateArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2210, \stateArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2212, \stateArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2072, \stateArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2076, \stateArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2080, \stateArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2084, \stateArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2088, \stateArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2092, \stateArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2096, \stateArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2100, \stateArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2103, \stateArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2106, \stateArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2109, \stateArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2112, \stateArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2115, \stateArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2118, \stateArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2121, \stateArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2124, \stateArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2126, \stateArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2128, \stateArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2130, \stateArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2132, \stateArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2134, \stateArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2136, \stateArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2138, \stateArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2140, \stateArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2246, \stateArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2248, \stateArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2250, \stateArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2252, \stateArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2254, \stateArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2256, \stateArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2258, \stateArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2260, \stateArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2237, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1371, \KeyArray/S00reg/gen_ff[1].gff/GEN[0].SFF/Q_401 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2238, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1368, \KeyArray/S00reg/gen_ff[1].gff/GEN[1].SFF/Q_400 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2239, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1365, \KeyArray/S00reg/gen_ff[1].gff/GEN[2].SFF/Q_399 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2240, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1362, \KeyArray/S00reg/gen_ff[1].gff/GEN[3].SFF/Q_398 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2241, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1359, \KeyArray/S00reg/gen_ff[1].gff/GEN[4].SFF/Q_397 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2242, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1356, \KeyArray/S00reg/gen_ff[1].gff/GEN[5].SFF/Q_396 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2243, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1353, \KeyArray/S00reg/gen_ff[1].gff/GEN[6].SFF/Q_395 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2244, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1350, \KeyArray/S00reg/gen_ff[1].gff/GEN[7].SFF/Q_394 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1528, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1805, \KeyArray/S01reg/gen_ff[1].gff/GEN[0].SFF/Q_691 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1532, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1808, \KeyArray/S01reg/gen_ff[1].gff/GEN[1].SFF/Q_692 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1536, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1811, \KeyArray/S01reg/gen_ff[1].gff/GEN[2].SFF/Q_693 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1540, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1814, \KeyArray/S01reg/gen_ff[1].gff/GEN[3].SFF/Q_694 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1544, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1817, \KeyArray/S01reg/gen_ff[1].gff/GEN[4].SFF/Q_695 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1548, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1820, \KeyArray/S01reg/gen_ff[1].gff/GEN[5].SFF/Q_696 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1552, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1823, \KeyArray/S01reg/gen_ff[1].gff/GEN[6].SFF/Q_697 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1556, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1826, \KeyArray/S01reg/gen_ff[1].gff/GEN[7].SFF/Q_698 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1560, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1526, \KeyArray/S02reg/gen_ff[1].gff/GEN[0].SFF/Q_683 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1564, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1530, \KeyArray/S02reg/gen_ff[1].gff/GEN[1].SFF/Q_684 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1568, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1534, \KeyArray/S02reg/gen_ff[1].gff/GEN[2].SFF/Q_685 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1572, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1538, \KeyArray/S02reg/gen_ff[1].gff/GEN[3].SFF/Q_686 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1576, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1542, \KeyArray/S02reg/gen_ff[1].gff/GEN[4].SFF/Q_687 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1580, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1546, \KeyArray/S02reg/gen_ff[1].gff/GEN[5].SFF/Q_688 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1584, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1550, \KeyArray/S02reg/gen_ff[1].gff/GEN[6].SFF/Q_689 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1588, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1554, \KeyArray/S02reg/gen_ff[1].gff/GEN[7].SFF/Q_690 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1591, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1558, \KeyArray/S03reg/gen_ff[1].gff/GEN[0].SFF/Q_675 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1594, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1562, \KeyArray/S03reg/gen_ff[1].gff/GEN[1].SFF/Q_676 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1597, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1566, \KeyArray/S03reg/gen_ff[1].gff/GEN[2].SFF/Q_677 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1600, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1570, \KeyArray/S03reg/gen_ff[1].gff/GEN[3].SFF/Q_678 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1603, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1574, \KeyArray/S03reg/gen_ff[1].gff/GEN[4].SFF/Q_679 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1606, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1578, \KeyArray/S03reg/gen_ff[1].gff/GEN[5].SFF/Q_680 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1609, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1582, \KeyArray/S03reg/gen_ff[1].gff/GEN[6].SFF/Q_681 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1612, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1586, \KeyArray/S03reg/gen_ff[1].gff/GEN[7].SFF/Q_682 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1615, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1589, \KeyArray/S10reg/gen_ff[1].gff/GEN[0].SFF/Q_667 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1618, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1592, \KeyArray/S10reg/gen_ff[1].gff/GEN[1].SFF/Q_668 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1621, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1595, \KeyArray/S10reg/gen_ff[1].gff/GEN[2].SFF/Q_669 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1624, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1598, \KeyArray/S10reg/gen_ff[1].gff/GEN[3].SFF/Q_670 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1627, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1601, \KeyArray/S10reg/gen_ff[1].gff/GEN[4].SFF/Q_671 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1630, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1604, \KeyArray/S10reg/gen_ff[1].gff/GEN[5].SFF/Q_672 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1633, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1607, \KeyArray/S10reg/gen_ff[1].gff/GEN[6].SFF/Q_673 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1636, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1610, \KeyArray/S10reg/gen_ff[1].gff/GEN[7].SFF/Q_674 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1639, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1525, \KeyArray/S11reg/gen_ff[1].gff/GEN[0].SFF/Q_659 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1642, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1529, \KeyArray/S11reg/gen_ff[1].gff/GEN[1].SFF/Q_660 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1645, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1533, \KeyArray/S11reg/gen_ff[1].gff/GEN[2].SFF/Q_661 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1648, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1537, \KeyArray/S11reg/gen_ff[1].gff/GEN[3].SFF/Q_662 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1651, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1541, \KeyArray/S11reg/gen_ff[1].gff/GEN[4].SFF/Q_663 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1654, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1545, \KeyArray/S11reg/gen_ff[1].gff/GEN[5].SFF/Q_664 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1657, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1549, \KeyArray/S11reg/gen_ff[1].gff/GEN[6].SFF/Q_665 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1660, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1553, \KeyArray/S11reg/gen_ff[1].gff/GEN[7].SFF/Q_666 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1663, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1557, \KeyArray/S12reg/gen_ff[1].gff/GEN[0].SFF/Q_651 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1666, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1561, \KeyArray/S12reg/gen_ff[1].gff/GEN[1].SFF/Q_652 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1669, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1565, \KeyArray/S12reg/gen_ff[1].gff/GEN[2].SFF/Q_653 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1672, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1569, \KeyArray/S12reg/gen_ff[1].gff/GEN[3].SFF/Q_654 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1675, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1573, \KeyArray/S12reg/gen_ff[1].gff/GEN[4].SFF/Q_655 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1678, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1577, \KeyArray/S12reg/gen_ff[1].gff/GEN[5].SFF/Q_656 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1681, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1581, \KeyArray/S12reg/gen_ff[1].gff/GEN[6].SFF/Q_657 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1684, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1585, \KeyArray/S12reg/gen_ff[1].gff/GEN[7].SFF/Q_658 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1687, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1433, \KeyArray/S13reg/gen_ff[1].gff/GEN[0].SFF/Q_393 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1690, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1431, \KeyArray/S13reg/gen_ff[1].gff/GEN[1].SFF/Q_392 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1693, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1429, \KeyArray/S13reg/gen_ff[1].gff/GEN[2].SFF/Q_391 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1696, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1427, \KeyArray/S13reg/gen_ff[1].gff/GEN[3].SFF/Q_390 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1699, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1425, \KeyArray/S13reg/gen_ff[1].gff/GEN[4].SFF/Q_389 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1702, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1423, \KeyArray/S13reg/gen_ff[1].gff/GEN[5].SFF/Q_388 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1705, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1437, \KeyArray/S13reg/gen_ff[1].gff/GEN[6].SFF/Q_387 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1708, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1435, \KeyArray/S13reg/gen_ff[1].gff/GEN[7].SFF/Q_386 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1711, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1613, \KeyArray/S20reg/gen_ff[1].gff/GEN[0].SFF/Q_643 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1714, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1616, \KeyArray/S20reg/gen_ff[1].gff/GEN[1].SFF/Q_644 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1717, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1619, \KeyArray/S20reg/gen_ff[1].gff/GEN[2].SFF/Q_645 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1720, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1622, \KeyArray/S20reg/gen_ff[1].gff/GEN[3].SFF/Q_646 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1723, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1625, \KeyArray/S20reg/gen_ff[1].gff/GEN[4].SFF/Q_647 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1726, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1628, \KeyArray/S20reg/gen_ff[1].gff/GEN[5].SFF/Q_648 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1729, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1631, \KeyArray/S20reg/gen_ff[1].gff/GEN[6].SFF/Q_649 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1732, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1634, \KeyArray/S20reg/gen_ff[1].gff/GEN[7].SFF/Q_650 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1735, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1637, \KeyArray/S21reg/gen_ff[1].gff/GEN[0].SFF/Q_635 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1738, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1640, \KeyArray/S21reg/gen_ff[1].gff/GEN[1].SFF/Q_636 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1741, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1643, \KeyArray/S21reg/gen_ff[1].gff/GEN[2].SFF/Q_637 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1744, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1646, \KeyArray/S21reg/gen_ff[1].gff/GEN[3].SFF/Q_638 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1747, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1649, \KeyArray/S21reg/gen_ff[1].gff/GEN[4].SFF/Q_639 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1750, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1652, \KeyArray/S21reg/gen_ff[1].gff/GEN[5].SFF/Q_640 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1753, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1655, \KeyArray/S21reg/gen_ff[1].gff/GEN[6].SFF/Q_641 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1756, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1658, \KeyArray/S21reg/gen_ff[1].gff/GEN[7].SFF/Q_642 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1759, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1661, \KeyArray/S22reg/gen_ff[1].gff/GEN[0].SFF/Q_627 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1762, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1664, \KeyArray/S22reg/gen_ff[1].gff/GEN[1].SFF/Q_628 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1765, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1667, \KeyArray/S22reg/gen_ff[1].gff/GEN[2].SFF/Q_629 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1768, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1670, \KeyArray/S22reg/gen_ff[1].gff/GEN[3].SFF/Q_630 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1771, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1673, \KeyArray/S22reg/gen_ff[1].gff/GEN[4].SFF/Q_631 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1774, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1676, \KeyArray/S22reg/gen_ff[1].gff/GEN[5].SFF/Q_632 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1777, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1679, \KeyArray/S22reg/gen_ff[1].gff/GEN[6].SFF/Q_633 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1780, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1682, \KeyArray/S22reg/gen_ff[1].gff/GEN[7].SFF/Q_634 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1783, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1685, \KeyArray/S23reg/gen_ff[1].gff/GEN[0].SFF/Q_619 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1786, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1688, \KeyArray/S23reg/gen_ff[1].gff/GEN[1].SFF/Q_620 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1789, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1691, \KeyArray/S23reg/gen_ff[1].gff/GEN[2].SFF/Q_621 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1792, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1694, \KeyArray/S23reg/gen_ff[1].gff/GEN[3].SFF/Q_622 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1795, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1697, \KeyArray/S23reg/gen_ff[1].gff/GEN[4].SFF/Q_623 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1798, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1700, \KeyArray/S23reg/gen_ff[1].gff/GEN[5].SFF/Q_624 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1801, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1703, \KeyArray/S23reg/gen_ff[1].gff/GEN[6].SFF/Q_625 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1804, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1706, \KeyArray/S23reg/gen_ff[1].gff/GEN[7].SFF/Q_626 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_2222, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1709, \KeyArray/S30reg/gen_ff[1].gff/GEN[0].SFF/Q_611 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_2224, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1712, \KeyArray/S30reg/gen_ff[1].gff/GEN[1].SFF/Q_612 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_2226, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1715, \KeyArray/S30reg/gen_ff[1].gff/GEN[2].SFF/Q_613 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_2228, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1718, \KeyArray/S30reg/gen_ff[1].gff/GEN[3].SFF/Q_614 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_2230, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1721, \KeyArray/S30reg/gen_ff[1].gff/GEN[4].SFF/Q_615 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_2232, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1724, \KeyArray/S30reg/gen_ff[1].gff/GEN[5].SFF/Q_616 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_2234, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1727, \KeyArray/S30reg/gen_ff[1].gff/GEN[6].SFF/Q_617 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_2236, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1730, \KeyArray/S30reg/gen_ff[1].gff/GEN[7].SFF/Q_618 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1807, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1733, \KeyArray/S31reg/gen_ff[1].gff/GEN[0].SFF/Q_603 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1810, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1736, \KeyArray/S31reg/gen_ff[1].gff/GEN[1].SFF/Q_604 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1813, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1739, \KeyArray/S31reg/gen_ff[1].gff/GEN[2].SFF/Q_605 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1816, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1742, \KeyArray/S31reg/gen_ff[1].gff/GEN[3].SFF/Q_606 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1819, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1745, \KeyArray/S31reg/gen_ff[1].gff/GEN[4].SFF/Q_607 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1822, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1748, \KeyArray/S31reg/gen_ff[1].gff/GEN[5].SFF/Q_608 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1825, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1751, \KeyArray/S31reg/gen_ff[1].gff/GEN[6].SFF/Q_609 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1828, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1754, \KeyArray/S31reg/gen_ff[1].gff/GEN[7].SFF/Q_610 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1830, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1757, \KeyArray/S32reg/gen_ff[1].gff/GEN[0].SFF/Q_595 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1832, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1760, \KeyArray/S32reg/gen_ff[1].gff/GEN[1].SFF/Q_596 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1834, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1763, \KeyArray/S32reg/gen_ff[1].gff/GEN[2].SFF/Q_597 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1836, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1766, \KeyArray/S32reg/gen_ff[1].gff/GEN[3].SFF/Q_598 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1838, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1769, \KeyArray/S32reg/gen_ff[1].gff/GEN[4].SFF/Q_599 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1840, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1772, \KeyArray/S32reg/gen_ff[1].gff/GEN[5].SFF/Q_600 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1842, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1775, \KeyArray/S32reg/gen_ff[1].gff/GEN[6].SFF/Q_601 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1844, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1778, \KeyArray/S32reg/gen_ff[1].gff/GEN[7].SFF/Q_602 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q ( .D ({new_AGEMA_signal_1846, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1781, \KeyArray/S33reg/gen_ff[1].gff/GEN[0].SFF/Q_587 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q ( .D ({new_AGEMA_signal_1848, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1784, \KeyArray/S33reg/gen_ff[1].gff/GEN[1].SFF/Q_588 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q ( .D ({new_AGEMA_signal_1850, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1787, \KeyArray/S33reg/gen_ff[1].gff/GEN[2].SFF/Q_589 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q ( .D ({new_AGEMA_signal_1852, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1790, \KeyArray/S33reg/gen_ff[1].gff/GEN[3].SFF/Q_590 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q ( .D ({new_AGEMA_signal_1854, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1793, \KeyArray/S33reg/gen_ff[1].gff/GEN[4].SFF/Q_591 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q ( .D ({new_AGEMA_signal_1856, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1796, \KeyArray/S33reg/gen_ff[1].gff/GEN[5].SFF/Q_592 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q ( .D ({new_AGEMA_signal_1858, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1799, \KeyArray/S33reg/gen_ff[1].gff/GEN[6].SFF/Q_593 }) ) ;
    FDE_masked #(.low_latency(0), .pipeline(0)) \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q ( .D ({new_AGEMA_signal_1860, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/QD }), .clk (clk_gated), .CE (enKS), .Q ({new_AGEMA_signal_1802, \KeyArray/S33reg/gen_ff[1].gff/GEN[7].SFF/Q_594 }) ) ;
    FD \ctrl/seq4/GEN[1].SFF/Q ( .D (\ctrl/seq4/GEN[1].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq4/GEN[1].SFF/Q_837 ) ) ;
    FD \ctrl/seq4/GEN[0].SFF/Q ( .D (\ctrl/seq4/GEN[0].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq4/GEN[0].SFF/Q_836 ) ) ;
    FD \ctrl/seq6/GEN[4].SFF/Q ( .D (\ctrl/seq6/GEN[4].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[4].SFF/Q_842 ) ) ;
    FD \ctrl/seq6/GEN[3].SFF/Q ( .D (\ctrl/seq6/GEN[3].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[3].SFF/Q_840 ) ) ;
    FD \ctrl/seq6/GEN[2].SFF/Q ( .D (\ctrl/seq6/GEN[2].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[2].SFF/Q_839 ) ) ;
    FD \ctrl/seq6/GEN[1].SFF/Q ( .D (\ctrl/seq6/GEN[1].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[1].SFF/Q_838 ) ) ;
    FD \ctrl/seq6/GEN[0].SFF/Q ( .D (\ctrl/seq6/GEN[0].SFF/QD ), .C (clk_gated), .Q (\ctrl/seq6/GEN[0].SFF/Q_841 ) ) ;
    FDR \ctrl/CSenRC ( .D (\ctrl/finalStep1 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSenRC_405 ) ) ;
    FDSE \calcRCon/s_current_state_7 ( .D (\calcRCon/s_current_state [6]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [7]) ) ;
    FDRE \calcRCon/s_current_state_6 ( .D (\calcRCon/s_current_state [5]), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [6]) ) ;
    FDRE \calcRCon/s_current_state_5 ( .D (\calcRCon/s_current_state [4]), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [5]) ) ;
    FDRE \calcRCon/s_current_state_4 ( .D (\calcRCon/MSB_s_current_state[3]_XOR_19_o ), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [4]) ) ;
    FDSE \calcRCon/s_current_state_3 ( .D (\calcRCon/MSB_s_current_state[2]_XOR_20_o ), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [3]) ) ;
    FDSE \calcRCon/s_current_state_2 ( .D (\calcRCon/s_current_state [1]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [2]) ) ;
    FDRE \calcRCon/s_current_state_1 ( .D (\calcRCon/MSB_s_current_state[0]_XOR_21_o ), .C (clk_gated), .CE (selSR), .R (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [1]) ) ;
    FDSE \calcRCon/s_current_state_0 ( .D (\calcRCon/s_current_state [7]), .C (clk_gated), .CE (selSR), .S (\calcRCon/nReset_inv ), .Q (\calcRCon/s_current_state [0]) ) ;
    FDR \ctrl/CSselMC ( .D (\ctrl/CSselMC_rstpot_1330 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSselMC_835 ) ) ;
    FD nReset ( .D (nReset_rstpot), .C (clk_gated), .Q (nReset_407) ) ;
    FD nReset_1 ( .D (nReset_rstpot), .C (clk_gated), .Q (nReset_1_1341) ) ;
    FDR \ctrl/CSselMC_1 ( .D (\ctrl/CSselMC_rstpot_1330 ), .C (clk_gated), .R (\calcRCon/nReset_inv ), .Q (\ctrl/CSselMC_1_1342 ) ) ;
endmodule
