/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC1_Pipeline_d4 (SI_s0, clk, SI_s1, SI_s2, SI_s3, SI_s4, Fresh, SO_s0, SO_s1, SO_s2, SO_s3, SO_s4);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [7:0] SI_s4 ;
    input [13019:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    output [7:0] SO_s4 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_17702 ;
    wire new_AGEMA_signal_17703 ;
    wire new_AGEMA_signal_17704 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17708 ;
    wire new_AGEMA_signal_17709 ;
    wire new_AGEMA_signal_17710 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17714 ;
    wire new_AGEMA_signal_17715 ;
    wire new_AGEMA_signal_17716 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17720 ;
    wire new_AGEMA_signal_17721 ;
    wire new_AGEMA_signal_17722 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17726 ;
    wire new_AGEMA_signal_17727 ;
    wire new_AGEMA_signal_17728 ;
    wire new_AGEMA_signal_17729 ;
    wire new_AGEMA_signal_17730 ;
    wire new_AGEMA_signal_17731 ;
    wire new_AGEMA_signal_17732 ;
    wire new_AGEMA_signal_17733 ;
    wire new_AGEMA_signal_17734 ;
    wire new_AGEMA_signal_17735 ;
    wire new_AGEMA_signal_17736 ;
    wire new_AGEMA_signal_17737 ;
    wire new_AGEMA_signal_17738 ;
    wire new_AGEMA_signal_17739 ;
    wire new_AGEMA_signal_17740 ;
    wire new_AGEMA_signal_17741 ;
    wire new_AGEMA_signal_17742 ;
    wire new_AGEMA_signal_17743 ;
    wire new_AGEMA_signal_17744 ;
    wire new_AGEMA_signal_17745 ;
    wire new_AGEMA_signal_17746 ;
    wire new_AGEMA_signal_17747 ;
    wire new_AGEMA_signal_17748 ;
    wire new_AGEMA_signal_17749 ;
    wire new_AGEMA_signal_17750 ;
    wire new_AGEMA_signal_17751 ;
    wire new_AGEMA_signal_17752 ;
    wire new_AGEMA_signal_17753 ;
    wire new_AGEMA_signal_17754 ;
    wire new_AGEMA_signal_17755 ;
    wire new_AGEMA_signal_17756 ;
    wire new_AGEMA_signal_17757 ;
    wire new_AGEMA_signal_17758 ;
    wire new_AGEMA_signal_17759 ;
    wire new_AGEMA_signal_17760 ;
    wire new_AGEMA_signal_17761 ;
    wire new_AGEMA_signal_17762 ;
    wire new_AGEMA_signal_17763 ;
    wire new_AGEMA_signal_17764 ;
    wire new_AGEMA_signal_17765 ;
    wire new_AGEMA_signal_17766 ;
    wire new_AGEMA_signal_17767 ;
    wire new_AGEMA_signal_17768 ;
    wire new_AGEMA_signal_17769 ;
    wire new_AGEMA_signal_17770 ;
    wire new_AGEMA_signal_17771 ;
    wire new_AGEMA_signal_17772 ;
    wire new_AGEMA_signal_17773 ;
    wire new_AGEMA_signal_17774 ;
    wire new_AGEMA_signal_17775 ;
    wire new_AGEMA_signal_17776 ;
    wire new_AGEMA_signal_17777 ;
    wire new_AGEMA_signal_17778 ;
    wire new_AGEMA_signal_17779 ;
    wire new_AGEMA_signal_17780 ;
    wire new_AGEMA_signal_17781 ;
    wire new_AGEMA_signal_17782 ;
    wire new_AGEMA_signal_17783 ;
    wire new_AGEMA_signal_17784 ;
    wire new_AGEMA_signal_17785 ;
    wire new_AGEMA_signal_17786 ;
    wire new_AGEMA_signal_17787 ;
    wire new_AGEMA_signal_17788 ;
    wire new_AGEMA_signal_17789 ;
    wire new_AGEMA_signal_17790 ;
    wire new_AGEMA_signal_17791 ;
    wire new_AGEMA_signal_17792 ;
    wire new_AGEMA_signal_17793 ;
    wire new_AGEMA_signal_17794 ;
    wire new_AGEMA_signal_17795 ;
    wire new_AGEMA_signal_17796 ;
    wire new_AGEMA_signal_17797 ;
    wire new_AGEMA_signal_17798 ;
    wire new_AGEMA_signal_17799 ;
    wire new_AGEMA_signal_17800 ;
    wire new_AGEMA_signal_17801 ;
    wire new_AGEMA_signal_17802 ;
    wire new_AGEMA_signal_17803 ;
    wire new_AGEMA_signal_17804 ;
    wire new_AGEMA_signal_17805 ;
    wire new_AGEMA_signal_17806 ;
    wire new_AGEMA_signal_17807 ;
    wire new_AGEMA_signal_17808 ;
    wire new_AGEMA_signal_17809 ;
    wire new_AGEMA_signal_17810 ;
    wire new_AGEMA_signal_17811 ;
    wire new_AGEMA_signal_17812 ;
    wire new_AGEMA_signal_17813 ;
    wire new_AGEMA_signal_17814 ;
    wire new_AGEMA_signal_17815 ;
    wire new_AGEMA_signal_17816 ;
    wire new_AGEMA_signal_17817 ;
    wire new_AGEMA_signal_17818 ;
    wire new_AGEMA_signal_17819 ;
    wire new_AGEMA_signal_17820 ;
    wire new_AGEMA_signal_17821 ;
    wire new_AGEMA_signal_17822 ;
    wire new_AGEMA_signal_17823 ;
    wire new_AGEMA_signal_17824 ;
    wire new_AGEMA_signal_17825 ;
    wire new_AGEMA_signal_17826 ;
    wire new_AGEMA_signal_17827 ;
    wire new_AGEMA_signal_17828 ;
    wire new_AGEMA_signal_17829 ;
    wire new_AGEMA_signal_17830 ;
    wire new_AGEMA_signal_17831 ;
    wire new_AGEMA_signal_17832 ;
    wire new_AGEMA_signal_17833 ;
    wire new_AGEMA_signal_17834 ;
    wire new_AGEMA_signal_17835 ;
    wire new_AGEMA_signal_17836 ;
    wire new_AGEMA_signal_17837 ;
    wire new_AGEMA_signal_17838 ;
    wire new_AGEMA_signal_17839 ;
    wire new_AGEMA_signal_17840 ;
    wire new_AGEMA_signal_17841 ;
    wire new_AGEMA_signal_17842 ;
    wire new_AGEMA_signal_17843 ;
    wire new_AGEMA_signal_17844 ;
    wire new_AGEMA_signal_17845 ;
    wire new_AGEMA_signal_17846 ;
    wire new_AGEMA_signal_17847 ;
    wire new_AGEMA_signal_17848 ;
    wire new_AGEMA_signal_17849 ;
    wire new_AGEMA_signal_17850 ;
    wire new_AGEMA_signal_17851 ;
    wire new_AGEMA_signal_17852 ;
    wire new_AGEMA_signal_17853 ;
    wire new_AGEMA_signal_17854 ;
    wire new_AGEMA_signal_17855 ;
    wire new_AGEMA_signal_17856 ;
    wire new_AGEMA_signal_17857 ;
    wire new_AGEMA_signal_17858 ;
    wire new_AGEMA_signal_17859 ;
    wire new_AGEMA_signal_17860 ;
    wire new_AGEMA_signal_17861 ;
    wire new_AGEMA_signal_17862 ;
    wire new_AGEMA_signal_17863 ;
    wire new_AGEMA_signal_17864 ;
    wire new_AGEMA_signal_17865 ;
    wire new_AGEMA_signal_17866 ;
    wire new_AGEMA_signal_17867 ;
    wire new_AGEMA_signal_17868 ;
    wire new_AGEMA_signal_17869 ;
    wire new_AGEMA_signal_17870 ;
    wire new_AGEMA_signal_17871 ;
    wire new_AGEMA_signal_17872 ;
    wire new_AGEMA_signal_17873 ;
    wire new_AGEMA_signal_17874 ;
    wire new_AGEMA_signal_17875 ;
    wire new_AGEMA_signal_17876 ;
    wire new_AGEMA_signal_17877 ;
    wire new_AGEMA_signal_17878 ;
    wire new_AGEMA_signal_17879 ;
    wire new_AGEMA_signal_17880 ;
    wire new_AGEMA_signal_17881 ;
    wire new_AGEMA_signal_17882 ;
    wire new_AGEMA_signal_17883 ;
    wire new_AGEMA_signal_17884 ;
    wire new_AGEMA_signal_17885 ;
    wire new_AGEMA_signal_17886 ;
    wire new_AGEMA_signal_17887 ;
    wire new_AGEMA_signal_17888 ;
    wire new_AGEMA_signal_17889 ;
    wire new_AGEMA_signal_17890 ;
    wire new_AGEMA_signal_17891 ;
    wire new_AGEMA_signal_17892 ;
    wire new_AGEMA_signal_17893 ;
    wire new_AGEMA_signal_17894 ;
    wire new_AGEMA_signal_17895 ;
    wire new_AGEMA_signal_17896 ;
    wire new_AGEMA_signal_17897 ;
    wire new_AGEMA_signal_17898 ;
    wire new_AGEMA_signal_17899 ;
    wire new_AGEMA_signal_17900 ;
    wire new_AGEMA_signal_17901 ;
    wire new_AGEMA_signal_17902 ;
    wire new_AGEMA_signal_17903 ;
    wire new_AGEMA_signal_17904 ;
    wire new_AGEMA_signal_17905 ;
    wire new_AGEMA_signal_17906 ;
    wire new_AGEMA_signal_17907 ;
    wire new_AGEMA_signal_17908 ;
    wire new_AGEMA_signal_17909 ;
    wire new_AGEMA_signal_17910 ;
    wire new_AGEMA_signal_17911 ;
    wire new_AGEMA_signal_17912 ;
    wire new_AGEMA_signal_17913 ;
    wire new_AGEMA_signal_17914 ;
    wire new_AGEMA_signal_17915 ;
    wire new_AGEMA_signal_17916 ;
    wire new_AGEMA_signal_17917 ;
    wire new_AGEMA_signal_17918 ;
    wire new_AGEMA_signal_17919 ;
    wire new_AGEMA_signal_17920 ;
    wire new_AGEMA_signal_17921 ;
    wire new_AGEMA_signal_17922 ;
    wire new_AGEMA_signal_17923 ;
    wire new_AGEMA_signal_17924 ;
    wire new_AGEMA_signal_17925 ;
    wire new_AGEMA_signal_17926 ;
    wire new_AGEMA_signal_17927 ;
    wire new_AGEMA_signal_17928 ;
    wire new_AGEMA_signal_17929 ;
    wire new_AGEMA_signal_17930 ;
    wire new_AGEMA_signal_17931 ;
    wire new_AGEMA_signal_17932 ;
    wire new_AGEMA_signal_17933 ;
    wire new_AGEMA_signal_17934 ;
    wire new_AGEMA_signal_17935 ;
    wire new_AGEMA_signal_17936 ;
    wire new_AGEMA_signal_17937 ;
    wire new_AGEMA_signal_17938 ;
    wire new_AGEMA_signal_17939 ;
    wire new_AGEMA_signal_17940 ;
    wire new_AGEMA_signal_17941 ;
    wire new_AGEMA_signal_17942 ;
    wire new_AGEMA_signal_17943 ;
    wire new_AGEMA_signal_17944 ;
    wire new_AGEMA_signal_17945 ;
    wire new_AGEMA_signal_17946 ;
    wire new_AGEMA_signal_17947 ;
    wire new_AGEMA_signal_17948 ;
    wire new_AGEMA_signal_17949 ;
    wire new_AGEMA_signal_17950 ;
    wire new_AGEMA_signal_17951 ;
    wire new_AGEMA_signal_17952 ;
    wire new_AGEMA_signal_17953 ;
    wire new_AGEMA_signal_17954 ;
    wire new_AGEMA_signal_17955 ;
    wire new_AGEMA_signal_17956 ;
    wire new_AGEMA_signal_17957 ;
    wire new_AGEMA_signal_17958 ;
    wire new_AGEMA_signal_17959 ;
    wire new_AGEMA_signal_17960 ;
    wire new_AGEMA_signal_17961 ;
    wire new_AGEMA_signal_17962 ;
    wire new_AGEMA_signal_17963 ;
    wire new_AGEMA_signal_17964 ;
    wire new_AGEMA_signal_17965 ;
    wire new_AGEMA_signal_17966 ;
    wire new_AGEMA_signal_17967 ;
    wire new_AGEMA_signal_17968 ;
    wire new_AGEMA_signal_17969 ;
    wire new_AGEMA_signal_17970 ;
    wire new_AGEMA_signal_17971 ;
    wire new_AGEMA_signal_17972 ;
    wire new_AGEMA_signal_17973 ;
    wire new_AGEMA_signal_17974 ;
    wire new_AGEMA_signal_17975 ;
    wire new_AGEMA_signal_17976 ;
    wire new_AGEMA_signal_17977 ;
    wire new_AGEMA_signal_17978 ;
    wire new_AGEMA_signal_17979 ;
    wire new_AGEMA_signal_17980 ;
    wire new_AGEMA_signal_17981 ;
    wire new_AGEMA_signal_17982 ;
    wire new_AGEMA_signal_17983 ;
    wire new_AGEMA_signal_17984 ;
    wire new_AGEMA_signal_17985 ;
    wire new_AGEMA_signal_17986 ;
    wire new_AGEMA_signal_17987 ;
    wire new_AGEMA_signal_17988 ;
    wire new_AGEMA_signal_17989 ;
    wire new_AGEMA_signal_17990 ;
    wire new_AGEMA_signal_17991 ;
    wire new_AGEMA_signal_17992 ;
    wire new_AGEMA_signal_17993 ;
    wire new_AGEMA_signal_17994 ;
    wire new_AGEMA_signal_17995 ;
    wire new_AGEMA_signal_17996 ;
    wire new_AGEMA_signal_17997 ;
    wire new_AGEMA_signal_17998 ;
    wire new_AGEMA_signal_17999 ;
    wire new_AGEMA_signal_18000 ;
    wire new_AGEMA_signal_18001 ;
    wire new_AGEMA_signal_18002 ;
    wire new_AGEMA_signal_18003 ;
    wire new_AGEMA_signal_18004 ;
    wire new_AGEMA_signal_18005 ;
    wire new_AGEMA_signal_18006 ;
    wire new_AGEMA_signal_18007 ;
    wire new_AGEMA_signal_18008 ;
    wire new_AGEMA_signal_18009 ;
    wire new_AGEMA_signal_18010 ;
    wire new_AGEMA_signal_18011 ;
    wire new_AGEMA_signal_18012 ;
    wire new_AGEMA_signal_18013 ;
    wire new_AGEMA_signal_18014 ;
    wire new_AGEMA_signal_18015 ;
    wire new_AGEMA_signal_18016 ;
    wire new_AGEMA_signal_18017 ;
    wire new_AGEMA_signal_18018 ;
    wire new_AGEMA_signal_18019 ;
    wire new_AGEMA_signal_18020 ;
    wire new_AGEMA_signal_18021 ;
    wire new_AGEMA_signal_18022 ;
    wire new_AGEMA_signal_18023 ;
    wire new_AGEMA_signal_18024 ;
    wire new_AGEMA_signal_18025 ;
    wire new_AGEMA_signal_18026 ;
    wire new_AGEMA_signal_18027 ;
    wire new_AGEMA_signal_18028 ;
    wire new_AGEMA_signal_18029 ;
    wire new_AGEMA_signal_18030 ;
    wire new_AGEMA_signal_18031 ;
    wire new_AGEMA_signal_18032 ;
    wire new_AGEMA_signal_18033 ;
    wire new_AGEMA_signal_18034 ;
    wire new_AGEMA_signal_18035 ;
    wire new_AGEMA_signal_18036 ;
    wire new_AGEMA_signal_18037 ;
    wire new_AGEMA_signal_18038 ;
    wire new_AGEMA_signal_18039 ;
    wire new_AGEMA_signal_18040 ;
    wire new_AGEMA_signal_18041 ;
    wire new_AGEMA_signal_18042 ;
    wire new_AGEMA_signal_18043 ;
    wire new_AGEMA_signal_18044 ;
    wire new_AGEMA_signal_18045 ;
    wire new_AGEMA_signal_18046 ;
    wire new_AGEMA_signal_18047 ;
    wire new_AGEMA_signal_18048 ;
    wire new_AGEMA_signal_18049 ;
    wire new_AGEMA_signal_18050 ;
    wire new_AGEMA_signal_18051 ;
    wire new_AGEMA_signal_18052 ;
    wire new_AGEMA_signal_18053 ;
    wire new_AGEMA_signal_18054 ;
    wire new_AGEMA_signal_18055 ;
    wire new_AGEMA_signal_18056 ;
    wire new_AGEMA_signal_18057 ;
    wire new_AGEMA_signal_18058 ;
    wire new_AGEMA_signal_18059 ;
    wire new_AGEMA_signal_18060 ;
    wire new_AGEMA_signal_18061 ;
    wire new_AGEMA_signal_18062 ;
    wire new_AGEMA_signal_18063 ;
    wire new_AGEMA_signal_18064 ;
    wire new_AGEMA_signal_18065 ;
    wire new_AGEMA_signal_18066 ;
    wire new_AGEMA_signal_18067 ;
    wire new_AGEMA_signal_18068 ;
    wire new_AGEMA_signal_18069 ;
    wire new_AGEMA_signal_18070 ;
    wire new_AGEMA_signal_18071 ;
    wire new_AGEMA_signal_18072 ;
    wire new_AGEMA_signal_18073 ;
    wire new_AGEMA_signal_18074 ;
    wire new_AGEMA_signal_18075 ;
    wire new_AGEMA_signal_18076 ;
    wire new_AGEMA_signal_18077 ;
    wire new_AGEMA_signal_18078 ;
    wire new_AGEMA_signal_18079 ;
    wire new_AGEMA_signal_18080 ;
    wire new_AGEMA_signal_18081 ;
    wire new_AGEMA_signal_18082 ;
    wire new_AGEMA_signal_18083 ;
    wire new_AGEMA_signal_18084 ;
    wire new_AGEMA_signal_18085 ;
    wire new_AGEMA_signal_18086 ;
    wire new_AGEMA_signal_18087 ;
    wire new_AGEMA_signal_18088 ;
    wire new_AGEMA_signal_18089 ;
    wire new_AGEMA_signal_18090 ;
    wire new_AGEMA_signal_18091 ;
    wire new_AGEMA_signal_18092 ;
    wire new_AGEMA_signal_18093 ;
    wire new_AGEMA_signal_18094 ;
    wire new_AGEMA_signal_18095 ;
    wire new_AGEMA_signal_18096 ;
    wire new_AGEMA_signal_18097 ;
    wire new_AGEMA_signal_18098 ;
    wire new_AGEMA_signal_18099 ;
    wire new_AGEMA_signal_18100 ;
    wire new_AGEMA_signal_18101 ;
    wire new_AGEMA_signal_18102 ;
    wire new_AGEMA_signal_18103 ;
    wire new_AGEMA_signal_18104 ;
    wire new_AGEMA_signal_18105 ;
    wire new_AGEMA_signal_18106 ;
    wire new_AGEMA_signal_18107 ;
    wire new_AGEMA_signal_18108 ;
    wire new_AGEMA_signal_18109 ;
    wire new_AGEMA_signal_18110 ;
    wire new_AGEMA_signal_18111 ;
    wire new_AGEMA_signal_18112 ;
    wire new_AGEMA_signal_18113 ;
    wire new_AGEMA_signal_18114 ;
    wire new_AGEMA_signal_18115 ;
    wire new_AGEMA_signal_18116 ;
    wire new_AGEMA_signal_18117 ;
    wire new_AGEMA_signal_18118 ;
    wire new_AGEMA_signal_18119 ;
    wire new_AGEMA_signal_18120 ;
    wire new_AGEMA_signal_18121 ;
    wire new_AGEMA_signal_18122 ;
    wire new_AGEMA_signal_18123 ;
    wire new_AGEMA_signal_18124 ;
    wire new_AGEMA_signal_18125 ;
    wire new_AGEMA_signal_18126 ;
    wire new_AGEMA_signal_18127 ;
    wire new_AGEMA_signal_18128 ;
    wire new_AGEMA_signal_18129 ;
    wire new_AGEMA_signal_18130 ;
    wire new_AGEMA_signal_18131 ;
    wire new_AGEMA_signal_18132 ;
    wire new_AGEMA_signal_18133 ;
    wire new_AGEMA_signal_18134 ;
    wire new_AGEMA_signal_18135 ;
    wire new_AGEMA_signal_18136 ;
    wire new_AGEMA_signal_18137 ;
    wire new_AGEMA_signal_18138 ;
    wire new_AGEMA_signal_18139 ;
    wire new_AGEMA_signal_18140 ;
    wire new_AGEMA_signal_18141 ;
    wire new_AGEMA_signal_18142 ;
    wire new_AGEMA_signal_18143 ;
    wire new_AGEMA_signal_18144 ;
    wire new_AGEMA_signal_18145 ;
    wire new_AGEMA_signal_18146 ;
    wire new_AGEMA_signal_18147 ;
    wire new_AGEMA_signal_18148 ;
    wire new_AGEMA_signal_18149 ;
    wire new_AGEMA_signal_18150 ;
    wire new_AGEMA_signal_18151 ;
    wire new_AGEMA_signal_18152 ;
    wire new_AGEMA_signal_18153 ;
    wire new_AGEMA_signal_18154 ;
    wire new_AGEMA_signal_18155 ;
    wire new_AGEMA_signal_18156 ;
    wire new_AGEMA_signal_18157 ;
    wire new_AGEMA_signal_18158 ;
    wire new_AGEMA_signal_18159 ;
    wire new_AGEMA_signal_18160 ;
    wire new_AGEMA_signal_18161 ;
    wire new_AGEMA_signal_18162 ;
    wire new_AGEMA_signal_18163 ;
    wire new_AGEMA_signal_18164 ;
    wire new_AGEMA_signal_18165 ;
    wire new_AGEMA_signal_18166 ;
    wire new_AGEMA_signal_18167 ;
    wire new_AGEMA_signal_18168 ;
    wire new_AGEMA_signal_18169 ;
    wire new_AGEMA_signal_18170 ;
    wire new_AGEMA_signal_18171 ;
    wire new_AGEMA_signal_18172 ;
    wire new_AGEMA_signal_18173 ;
    wire new_AGEMA_signal_18174 ;
    wire new_AGEMA_signal_18175 ;
    wire new_AGEMA_signal_18176 ;
    wire new_AGEMA_signal_18177 ;
    wire new_AGEMA_signal_18178 ;
    wire new_AGEMA_signal_18179 ;
    wire new_AGEMA_signal_18180 ;
    wire new_AGEMA_signal_18181 ;
    wire new_AGEMA_signal_18182 ;
    wire new_AGEMA_signal_18183 ;
    wire new_AGEMA_signal_18184 ;
    wire new_AGEMA_signal_18185 ;
    wire new_AGEMA_signal_18186 ;
    wire new_AGEMA_signal_18187 ;
    wire new_AGEMA_signal_18188 ;
    wire new_AGEMA_signal_18189 ;
    wire new_AGEMA_signal_18190 ;
    wire new_AGEMA_signal_18191 ;
    wire new_AGEMA_signal_18192 ;
    wire new_AGEMA_signal_18193 ;
    wire new_AGEMA_signal_18194 ;
    wire new_AGEMA_signal_18195 ;
    wire new_AGEMA_signal_18196 ;
    wire new_AGEMA_signal_18197 ;
    wire new_AGEMA_signal_18198 ;
    wire new_AGEMA_signal_18199 ;
    wire new_AGEMA_signal_18200 ;
    wire new_AGEMA_signal_18201 ;
    wire new_AGEMA_signal_18202 ;
    wire new_AGEMA_signal_18203 ;
    wire new_AGEMA_signal_18204 ;
    wire new_AGEMA_signal_18205 ;
    wire new_AGEMA_signal_18206 ;
    wire new_AGEMA_signal_18207 ;
    wire new_AGEMA_signal_18208 ;
    wire new_AGEMA_signal_18209 ;
    wire new_AGEMA_signal_18210 ;
    wire new_AGEMA_signal_18211 ;
    wire new_AGEMA_signal_18212 ;
    wire new_AGEMA_signal_18213 ;
    wire new_AGEMA_signal_18214 ;
    wire new_AGEMA_signal_18215 ;
    wire new_AGEMA_signal_18216 ;
    wire new_AGEMA_signal_18217 ;
    wire new_AGEMA_signal_18218 ;
    wire new_AGEMA_signal_18219 ;
    wire new_AGEMA_signal_18220 ;
    wire new_AGEMA_signal_18221 ;
    wire new_AGEMA_signal_18222 ;
    wire new_AGEMA_signal_18223 ;
    wire new_AGEMA_signal_18224 ;
    wire new_AGEMA_signal_18225 ;
    wire new_AGEMA_signal_18226 ;
    wire new_AGEMA_signal_18227 ;
    wire new_AGEMA_signal_18228 ;
    wire new_AGEMA_signal_18229 ;
    wire new_AGEMA_signal_18230 ;
    wire new_AGEMA_signal_18231 ;
    wire new_AGEMA_signal_18232 ;
    wire new_AGEMA_signal_18233 ;
    wire new_AGEMA_signal_18234 ;
    wire new_AGEMA_signal_18235 ;
    wire new_AGEMA_signal_18236 ;
    wire new_AGEMA_signal_18237 ;
    wire new_AGEMA_signal_18238 ;
    wire new_AGEMA_signal_18239 ;
    wire new_AGEMA_signal_18240 ;
    wire new_AGEMA_signal_18241 ;
    wire new_AGEMA_signal_18242 ;
    wire new_AGEMA_signal_18243 ;
    wire new_AGEMA_signal_18244 ;
    wire new_AGEMA_signal_18245 ;
    wire new_AGEMA_signal_18246 ;
    wire new_AGEMA_signal_18247 ;
    wire new_AGEMA_signal_18248 ;
    wire new_AGEMA_signal_18249 ;
    wire new_AGEMA_signal_18250 ;
    wire new_AGEMA_signal_18251 ;
    wire new_AGEMA_signal_18252 ;
    wire new_AGEMA_signal_18253 ;
    wire new_AGEMA_signal_18254 ;
    wire new_AGEMA_signal_18255 ;
    wire new_AGEMA_signal_18256 ;
    wire new_AGEMA_signal_18257 ;
    wire new_AGEMA_signal_18258 ;
    wire new_AGEMA_signal_18259 ;
    wire new_AGEMA_signal_18260 ;
    wire new_AGEMA_signal_18261 ;
    wire new_AGEMA_signal_18262 ;
    wire new_AGEMA_signal_18263 ;
    wire new_AGEMA_signal_18264 ;
    wire new_AGEMA_signal_18265 ;
    wire new_AGEMA_signal_18266 ;
    wire new_AGEMA_signal_18267 ;
    wire new_AGEMA_signal_18268 ;
    wire new_AGEMA_signal_18269 ;
    wire new_AGEMA_signal_18270 ;
    wire new_AGEMA_signal_18271 ;
    wire new_AGEMA_signal_18272 ;
    wire new_AGEMA_signal_18273 ;
    wire new_AGEMA_signal_18274 ;
    wire new_AGEMA_signal_18275 ;
    wire new_AGEMA_signal_18276 ;
    wire new_AGEMA_signal_18277 ;
    wire new_AGEMA_signal_18278 ;
    wire new_AGEMA_signal_18279 ;
    wire new_AGEMA_signal_18280 ;
    wire new_AGEMA_signal_18281 ;
    wire new_AGEMA_signal_18282 ;
    wire new_AGEMA_signal_18283 ;
    wire new_AGEMA_signal_18284 ;
    wire new_AGEMA_signal_18285 ;
    wire new_AGEMA_signal_18286 ;
    wire new_AGEMA_signal_18287 ;
    wire new_AGEMA_signal_18288 ;
    wire new_AGEMA_signal_18289 ;
    wire new_AGEMA_signal_18290 ;
    wire new_AGEMA_signal_18291 ;
    wire new_AGEMA_signal_18292 ;
    wire new_AGEMA_signal_18293 ;
    wire new_AGEMA_signal_18294 ;
    wire new_AGEMA_signal_18295 ;
    wire new_AGEMA_signal_18296 ;
    wire new_AGEMA_signal_18297 ;
    wire new_AGEMA_signal_18298 ;
    wire new_AGEMA_signal_18299 ;
    wire new_AGEMA_signal_18300 ;
    wire new_AGEMA_signal_18301 ;
    wire new_AGEMA_signal_18302 ;
    wire new_AGEMA_signal_18303 ;
    wire new_AGEMA_signal_18304 ;
    wire new_AGEMA_signal_18305 ;
    wire new_AGEMA_signal_18306 ;
    wire new_AGEMA_signal_18307 ;
    wire new_AGEMA_signal_18308 ;
    wire new_AGEMA_signal_18309 ;
    wire new_AGEMA_signal_18310 ;
    wire new_AGEMA_signal_18311 ;
    wire new_AGEMA_signal_18312 ;
    wire new_AGEMA_signal_18313 ;
    wire new_AGEMA_signal_18314 ;
    wire new_AGEMA_signal_18315 ;
    wire new_AGEMA_signal_18316 ;
    wire new_AGEMA_signal_18317 ;
    wire new_AGEMA_signal_18318 ;
    wire new_AGEMA_signal_18319 ;
    wire new_AGEMA_signal_18320 ;
    wire new_AGEMA_signal_18321 ;
    wire new_AGEMA_signal_18322 ;
    wire new_AGEMA_signal_18323 ;
    wire new_AGEMA_signal_18324 ;
    wire new_AGEMA_signal_18325 ;
    wire new_AGEMA_signal_18326 ;
    wire new_AGEMA_signal_18327 ;
    wire new_AGEMA_signal_18328 ;
    wire new_AGEMA_signal_18329 ;
    wire new_AGEMA_signal_18330 ;
    wire new_AGEMA_signal_18331 ;
    wire new_AGEMA_signal_18332 ;
    wire new_AGEMA_signal_18333 ;
    wire new_AGEMA_signal_18334 ;
    wire new_AGEMA_signal_18335 ;
    wire new_AGEMA_signal_18336 ;
    wire new_AGEMA_signal_18337 ;
    wire new_AGEMA_signal_18338 ;
    wire new_AGEMA_signal_18339 ;
    wire new_AGEMA_signal_18340 ;
    wire new_AGEMA_signal_18341 ;
    wire new_AGEMA_signal_18342 ;
    wire new_AGEMA_signal_18343 ;
    wire new_AGEMA_signal_18344 ;
    wire new_AGEMA_signal_18345 ;
    wire new_AGEMA_signal_18346 ;
    wire new_AGEMA_signal_18347 ;
    wire new_AGEMA_signal_18348 ;
    wire new_AGEMA_signal_18349 ;
    wire new_AGEMA_signal_18350 ;
    wire new_AGEMA_signal_18351 ;
    wire new_AGEMA_signal_18352 ;
    wire new_AGEMA_signal_18353 ;
    wire new_AGEMA_signal_18354 ;
    wire new_AGEMA_signal_18355 ;
    wire new_AGEMA_signal_18356 ;
    wire new_AGEMA_signal_18357 ;
    wire new_AGEMA_signal_18358 ;
    wire new_AGEMA_signal_18359 ;
    wire new_AGEMA_signal_18360 ;
    wire new_AGEMA_signal_18361 ;
    wire new_AGEMA_signal_18362 ;
    wire new_AGEMA_signal_18363 ;
    wire new_AGEMA_signal_18364 ;
    wire new_AGEMA_signal_18365 ;
    wire new_AGEMA_signal_18366 ;
    wire new_AGEMA_signal_18367 ;
    wire new_AGEMA_signal_18368 ;
    wire new_AGEMA_signal_18369 ;
    wire new_AGEMA_signal_18370 ;
    wire new_AGEMA_signal_18371 ;
    wire new_AGEMA_signal_18372 ;
    wire new_AGEMA_signal_18373 ;
    wire new_AGEMA_signal_18374 ;
    wire new_AGEMA_signal_18375 ;
    wire new_AGEMA_signal_18376 ;
    wire new_AGEMA_signal_18377 ;
    wire new_AGEMA_signal_18378 ;
    wire new_AGEMA_signal_18379 ;
    wire new_AGEMA_signal_18380 ;
    wire new_AGEMA_signal_18381 ;
    wire new_AGEMA_signal_18382 ;
    wire new_AGEMA_signal_18383 ;
    wire new_AGEMA_signal_18384 ;
    wire new_AGEMA_signal_18385 ;
    wire new_AGEMA_signal_18386 ;
    wire new_AGEMA_signal_18387 ;
    wire new_AGEMA_signal_18388 ;
    wire new_AGEMA_signal_18389 ;
    wire new_AGEMA_signal_18390 ;
    wire new_AGEMA_signal_18391 ;
    wire new_AGEMA_signal_18392 ;
    wire new_AGEMA_signal_18393 ;
    wire new_AGEMA_signal_18394 ;
    wire new_AGEMA_signal_18395 ;
    wire new_AGEMA_signal_18396 ;
    wire new_AGEMA_signal_18397 ;
    wire new_AGEMA_signal_18398 ;
    wire new_AGEMA_signal_18399 ;
    wire new_AGEMA_signal_18400 ;
    wire new_AGEMA_signal_18401 ;
    wire new_AGEMA_signal_18402 ;
    wire new_AGEMA_signal_18403 ;
    wire new_AGEMA_signal_18404 ;
    wire new_AGEMA_signal_18405 ;
    wire new_AGEMA_signal_18406 ;
    wire new_AGEMA_signal_18407 ;
    wire new_AGEMA_signal_18408 ;
    wire new_AGEMA_signal_18409 ;
    wire new_AGEMA_signal_18410 ;
    wire new_AGEMA_signal_18411 ;
    wire new_AGEMA_signal_18412 ;
    wire new_AGEMA_signal_18413 ;
    wire new_AGEMA_signal_18414 ;
    wire new_AGEMA_signal_18415 ;
    wire new_AGEMA_signal_18416 ;
    wire new_AGEMA_signal_18417 ;
    wire new_AGEMA_signal_18418 ;
    wire new_AGEMA_signal_18419 ;
    wire new_AGEMA_signal_18420 ;
    wire new_AGEMA_signal_18421 ;
    wire new_AGEMA_signal_18422 ;
    wire new_AGEMA_signal_18423 ;
    wire new_AGEMA_signal_18424 ;
    wire new_AGEMA_signal_18425 ;
    wire new_AGEMA_signal_18426 ;
    wire new_AGEMA_signal_18427 ;
    wire new_AGEMA_signal_18428 ;
    wire new_AGEMA_signal_18429 ;
    wire new_AGEMA_signal_18430 ;
    wire new_AGEMA_signal_18431 ;
    wire new_AGEMA_signal_18432 ;
    wire new_AGEMA_signal_18433 ;
    wire new_AGEMA_signal_18434 ;
    wire new_AGEMA_signal_18435 ;
    wire new_AGEMA_signal_18436 ;
    wire new_AGEMA_signal_18437 ;
    wire new_AGEMA_signal_18438 ;
    wire new_AGEMA_signal_18439 ;
    wire new_AGEMA_signal_18440 ;
    wire new_AGEMA_signal_18441 ;
    wire new_AGEMA_signal_18442 ;
    wire new_AGEMA_signal_18443 ;
    wire new_AGEMA_signal_18444 ;
    wire new_AGEMA_signal_18445 ;
    wire new_AGEMA_signal_18446 ;
    wire new_AGEMA_signal_18447 ;
    wire new_AGEMA_signal_18448 ;
    wire new_AGEMA_signal_18449 ;
    wire new_AGEMA_signal_18450 ;
    wire new_AGEMA_signal_18451 ;
    wire new_AGEMA_signal_18452 ;
    wire new_AGEMA_signal_18453 ;
    wire new_AGEMA_signal_18454 ;
    wire new_AGEMA_signal_18455 ;
    wire new_AGEMA_signal_18456 ;
    wire new_AGEMA_signal_18457 ;
    wire new_AGEMA_signal_18458 ;
    wire new_AGEMA_signal_18459 ;
    wire new_AGEMA_signal_18460 ;
    wire new_AGEMA_signal_18461 ;
    wire new_AGEMA_signal_18462 ;
    wire new_AGEMA_signal_18463 ;
    wire new_AGEMA_signal_18464 ;
    wire new_AGEMA_signal_18465 ;
    wire new_AGEMA_signal_18466 ;
    wire new_AGEMA_signal_18467 ;
    wire new_AGEMA_signal_18468 ;
    wire new_AGEMA_signal_18469 ;
    wire new_AGEMA_signal_18470 ;
    wire new_AGEMA_signal_18471 ;
    wire new_AGEMA_signal_18472 ;
    wire new_AGEMA_signal_18473 ;
    wire new_AGEMA_signal_18474 ;
    wire new_AGEMA_signal_18475 ;
    wire new_AGEMA_signal_18476 ;
    wire new_AGEMA_signal_18477 ;
    wire new_AGEMA_signal_18478 ;
    wire new_AGEMA_signal_18479 ;
    wire new_AGEMA_signal_18480 ;
    wire new_AGEMA_signal_18481 ;
    wire new_AGEMA_signal_18482 ;
    wire new_AGEMA_signal_18483 ;
    wire new_AGEMA_signal_18484 ;
    wire new_AGEMA_signal_18485 ;
    wire new_AGEMA_signal_18486 ;
    wire new_AGEMA_signal_18487 ;
    wire new_AGEMA_signal_18488 ;
    wire new_AGEMA_signal_18489 ;
    wire new_AGEMA_signal_18490 ;
    wire new_AGEMA_signal_18491 ;
    wire new_AGEMA_signal_18492 ;
    wire new_AGEMA_signal_18493 ;
    wire new_AGEMA_signal_18494 ;
    wire new_AGEMA_signal_18495 ;
    wire new_AGEMA_signal_18496 ;
    wire new_AGEMA_signal_18497 ;
    wire new_AGEMA_signal_18498 ;
    wire new_AGEMA_signal_18499 ;
    wire new_AGEMA_signal_18500 ;
    wire new_AGEMA_signal_18501 ;
    wire new_AGEMA_signal_18502 ;
    wire new_AGEMA_signal_18503 ;
    wire new_AGEMA_signal_18504 ;
    wire new_AGEMA_signal_18505 ;
    wire new_AGEMA_signal_18506 ;
    wire new_AGEMA_signal_18507 ;
    wire new_AGEMA_signal_18508 ;
    wire new_AGEMA_signal_18509 ;
    wire new_AGEMA_signal_18510 ;
    wire new_AGEMA_signal_18511 ;
    wire new_AGEMA_signal_18512 ;
    wire new_AGEMA_signal_18513 ;
    wire new_AGEMA_signal_18514 ;
    wire new_AGEMA_signal_18515 ;
    wire new_AGEMA_signal_18516 ;
    wire new_AGEMA_signal_18517 ;
    wire new_AGEMA_signal_18518 ;
    wire new_AGEMA_signal_18519 ;
    wire new_AGEMA_signal_18520 ;
    wire new_AGEMA_signal_18521 ;
    wire new_AGEMA_signal_18522 ;
    wire new_AGEMA_signal_18523 ;
    wire new_AGEMA_signal_18524 ;
    wire new_AGEMA_signal_18525 ;
    wire new_AGEMA_signal_18526 ;
    wire new_AGEMA_signal_18527 ;
    wire new_AGEMA_signal_18528 ;
    wire new_AGEMA_signal_18529 ;
    wire new_AGEMA_signal_18530 ;
    wire new_AGEMA_signal_18531 ;
    wire new_AGEMA_signal_18532 ;
    wire new_AGEMA_signal_18533 ;
    wire new_AGEMA_signal_18534 ;
    wire new_AGEMA_signal_18535 ;
    wire new_AGEMA_signal_18536 ;
    wire new_AGEMA_signal_18537 ;
    wire new_AGEMA_signal_18538 ;
    wire new_AGEMA_signal_18539 ;
    wire new_AGEMA_signal_18540 ;
    wire new_AGEMA_signal_18541 ;
    wire new_AGEMA_signal_18542 ;
    wire new_AGEMA_signal_18543 ;
    wire new_AGEMA_signal_18544 ;
    wire new_AGEMA_signal_18545 ;
    wire new_AGEMA_signal_18546 ;
    wire new_AGEMA_signal_18547 ;
    wire new_AGEMA_signal_18548 ;
    wire new_AGEMA_signal_18549 ;
    wire new_AGEMA_signal_18550 ;
    wire new_AGEMA_signal_18551 ;
    wire new_AGEMA_signal_18552 ;
    wire new_AGEMA_signal_18553 ;
    wire new_AGEMA_signal_18554 ;
    wire new_AGEMA_signal_18555 ;
    wire new_AGEMA_signal_18556 ;
    wire new_AGEMA_signal_18557 ;
    wire new_AGEMA_signal_18558 ;
    wire new_AGEMA_signal_18559 ;
    wire new_AGEMA_signal_18560 ;
    wire new_AGEMA_signal_18561 ;
    wire new_AGEMA_signal_18562 ;
    wire new_AGEMA_signal_18563 ;
    wire new_AGEMA_signal_18564 ;
    wire new_AGEMA_signal_18565 ;
    wire new_AGEMA_signal_18566 ;
    wire new_AGEMA_signal_18567 ;
    wire new_AGEMA_signal_18568 ;
    wire new_AGEMA_signal_18569 ;
    wire new_AGEMA_signal_18570 ;
    wire new_AGEMA_signal_18571 ;
    wire new_AGEMA_signal_18572 ;
    wire new_AGEMA_signal_18573 ;
    wire new_AGEMA_signal_18574 ;
    wire new_AGEMA_signal_18575 ;
    wire new_AGEMA_signal_18576 ;
    wire new_AGEMA_signal_18577 ;
    wire new_AGEMA_signal_18578 ;
    wire new_AGEMA_signal_18579 ;
    wire new_AGEMA_signal_18580 ;
    wire new_AGEMA_signal_18581 ;
    wire new_AGEMA_signal_18582 ;
    wire new_AGEMA_signal_18583 ;
    wire new_AGEMA_signal_18584 ;
    wire new_AGEMA_signal_18585 ;
    wire new_AGEMA_signal_18586 ;
    wire new_AGEMA_signal_18587 ;
    wire new_AGEMA_signal_18588 ;
    wire new_AGEMA_signal_18589 ;
    wire new_AGEMA_signal_18590 ;
    wire new_AGEMA_signal_18591 ;
    wire new_AGEMA_signal_18592 ;
    wire new_AGEMA_signal_18593 ;
    wire new_AGEMA_signal_18594 ;
    wire new_AGEMA_signal_18595 ;
    wire new_AGEMA_signal_18596 ;
    wire new_AGEMA_signal_18597 ;
    wire new_AGEMA_signal_18598 ;
    wire new_AGEMA_signal_18599 ;
    wire new_AGEMA_signal_18600 ;
    wire new_AGEMA_signal_18601 ;
    wire new_AGEMA_signal_18602 ;
    wire new_AGEMA_signal_18603 ;
    wire new_AGEMA_signal_18604 ;
    wire new_AGEMA_signal_18605 ;
    wire new_AGEMA_signal_18606 ;
    wire new_AGEMA_signal_18607 ;
    wire new_AGEMA_signal_18608 ;
    wire new_AGEMA_signal_18609 ;
    wire new_AGEMA_signal_18610 ;
    wire new_AGEMA_signal_18611 ;
    wire new_AGEMA_signal_18612 ;
    wire new_AGEMA_signal_18613 ;
    wire new_AGEMA_signal_18614 ;
    wire new_AGEMA_signal_18615 ;
    wire new_AGEMA_signal_18616 ;
    wire new_AGEMA_signal_18617 ;
    wire new_AGEMA_signal_18618 ;
    wire new_AGEMA_signal_18619 ;
    wire new_AGEMA_signal_18620 ;
    wire new_AGEMA_signal_18621 ;
    wire new_AGEMA_signal_18622 ;
    wire new_AGEMA_signal_18623 ;
    wire new_AGEMA_signal_18624 ;
    wire new_AGEMA_signal_18625 ;
    wire new_AGEMA_signal_18626 ;
    wire new_AGEMA_signal_18627 ;
    wire new_AGEMA_signal_18628 ;
    wire new_AGEMA_signal_18629 ;
    wire new_AGEMA_signal_18630 ;
    wire new_AGEMA_signal_18631 ;
    wire new_AGEMA_signal_18632 ;
    wire new_AGEMA_signal_18633 ;
    wire new_AGEMA_signal_18634 ;
    wire new_AGEMA_signal_18635 ;
    wire new_AGEMA_signal_18636 ;
    wire new_AGEMA_signal_18637 ;
    wire new_AGEMA_signal_18638 ;
    wire new_AGEMA_signal_18639 ;
    wire new_AGEMA_signal_18640 ;
    wire new_AGEMA_signal_18641 ;
    wire new_AGEMA_signal_18642 ;
    wire new_AGEMA_signal_18643 ;
    wire new_AGEMA_signal_18644 ;
    wire new_AGEMA_signal_18645 ;
    wire new_AGEMA_signal_18646 ;
    wire new_AGEMA_signal_18647 ;
    wire new_AGEMA_signal_18648 ;
    wire new_AGEMA_signal_18649 ;
    wire new_AGEMA_signal_18650 ;
    wire new_AGEMA_signal_18651 ;
    wire new_AGEMA_signal_18652 ;
    wire new_AGEMA_signal_18653 ;
    wire new_AGEMA_signal_18654 ;
    wire new_AGEMA_signal_18655 ;
    wire new_AGEMA_signal_18656 ;
    wire new_AGEMA_signal_18657 ;
    wire new_AGEMA_signal_18658 ;
    wire new_AGEMA_signal_18659 ;
    wire new_AGEMA_signal_18660 ;
    wire new_AGEMA_signal_18661 ;
    wire new_AGEMA_signal_18662 ;
    wire new_AGEMA_signal_18663 ;
    wire new_AGEMA_signal_18664 ;
    wire new_AGEMA_signal_18665 ;
    wire new_AGEMA_signal_18666 ;
    wire new_AGEMA_signal_18667 ;
    wire new_AGEMA_signal_18668 ;
    wire new_AGEMA_signal_18669 ;
    wire new_AGEMA_signal_18670 ;
    wire new_AGEMA_signal_18671 ;
    wire new_AGEMA_signal_18672 ;
    wire new_AGEMA_signal_18673 ;
    wire new_AGEMA_signal_18674 ;
    wire new_AGEMA_signal_18675 ;
    wire new_AGEMA_signal_18676 ;
    wire new_AGEMA_signal_18677 ;
    wire new_AGEMA_signal_18678 ;
    wire new_AGEMA_signal_18679 ;
    wire new_AGEMA_signal_18680 ;
    wire new_AGEMA_signal_18681 ;
    wire new_AGEMA_signal_18682 ;
    wire new_AGEMA_signal_18683 ;
    wire new_AGEMA_signal_18684 ;
    wire new_AGEMA_signal_18685 ;
    wire new_AGEMA_signal_18686 ;
    wire new_AGEMA_signal_18687 ;
    wire new_AGEMA_signal_18688 ;
    wire new_AGEMA_signal_18689 ;
    wire new_AGEMA_signal_18690 ;
    wire new_AGEMA_signal_18691 ;
    wire new_AGEMA_signal_18692 ;
    wire new_AGEMA_signal_18693 ;
    wire new_AGEMA_signal_18694 ;
    wire new_AGEMA_signal_18695 ;
    wire new_AGEMA_signal_18696 ;
    wire new_AGEMA_signal_18697 ;
    wire new_AGEMA_signal_18698 ;
    wire new_AGEMA_signal_18699 ;
    wire new_AGEMA_signal_18700 ;
    wire new_AGEMA_signal_18701 ;
    wire new_AGEMA_signal_18702 ;
    wire new_AGEMA_signal_18703 ;
    wire new_AGEMA_signal_18704 ;
    wire new_AGEMA_signal_18705 ;
    wire new_AGEMA_signal_18706 ;
    wire new_AGEMA_signal_18707 ;
    wire new_AGEMA_signal_18708 ;
    wire new_AGEMA_signal_18709 ;
    wire new_AGEMA_signal_18710 ;
    wire new_AGEMA_signal_18711 ;
    wire new_AGEMA_signal_18712 ;
    wire new_AGEMA_signal_18713 ;
    wire new_AGEMA_signal_18714 ;
    wire new_AGEMA_signal_18715 ;
    wire new_AGEMA_signal_18716 ;
    wire new_AGEMA_signal_18717 ;
    wire new_AGEMA_signal_18718 ;
    wire new_AGEMA_signal_18719 ;
    wire new_AGEMA_signal_18720 ;
    wire new_AGEMA_signal_18721 ;
    wire new_AGEMA_signal_18722 ;
    wire new_AGEMA_signal_18723 ;
    wire new_AGEMA_signal_18724 ;
    wire new_AGEMA_signal_18725 ;
    wire new_AGEMA_signal_18726 ;
    wire new_AGEMA_signal_18727 ;
    wire new_AGEMA_signal_18728 ;
    wire new_AGEMA_signal_18729 ;
    wire new_AGEMA_signal_18730 ;
    wire new_AGEMA_signal_18731 ;
    wire new_AGEMA_signal_18732 ;
    wire new_AGEMA_signal_18733 ;
    wire new_AGEMA_signal_18734 ;
    wire new_AGEMA_signal_18735 ;
    wire new_AGEMA_signal_18736 ;
    wire new_AGEMA_signal_18737 ;
    wire new_AGEMA_signal_18738 ;
    wire new_AGEMA_signal_18739 ;
    wire new_AGEMA_signal_18740 ;
    wire new_AGEMA_signal_18741 ;
    wire new_AGEMA_signal_18742 ;
    wire new_AGEMA_signal_18743 ;
    wire new_AGEMA_signal_18744 ;
    wire new_AGEMA_signal_18745 ;
    wire new_AGEMA_signal_18746 ;
    wire new_AGEMA_signal_18747 ;
    wire new_AGEMA_signal_18748 ;
    wire new_AGEMA_signal_18749 ;
    wire new_AGEMA_signal_18750 ;
    wire new_AGEMA_signal_18751 ;
    wire new_AGEMA_signal_18752 ;
    wire new_AGEMA_signal_18753 ;
    wire new_AGEMA_signal_18754 ;
    wire new_AGEMA_signal_18755 ;
    wire new_AGEMA_signal_18756 ;
    wire new_AGEMA_signal_18757 ;
    wire new_AGEMA_signal_18758 ;
    wire new_AGEMA_signal_18759 ;
    wire new_AGEMA_signal_18760 ;
    wire new_AGEMA_signal_18761 ;
    wire new_AGEMA_signal_18762 ;
    wire new_AGEMA_signal_18763 ;
    wire new_AGEMA_signal_18764 ;
    wire new_AGEMA_signal_18765 ;
    wire new_AGEMA_signal_18766 ;
    wire new_AGEMA_signal_18767 ;
    wire new_AGEMA_signal_18768 ;
    wire new_AGEMA_signal_18769 ;
    wire new_AGEMA_signal_18770 ;
    wire new_AGEMA_signal_18771 ;
    wire new_AGEMA_signal_18772 ;
    wire new_AGEMA_signal_18773 ;
    wire new_AGEMA_signal_18774 ;
    wire new_AGEMA_signal_18775 ;
    wire new_AGEMA_signal_18776 ;
    wire new_AGEMA_signal_18777 ;
    wire new_AGEMA_signal_18778 ;
    wire new_AGEMA_signal_18779 ;
    wire new_AGEMA_signal_18780 ;
    wire new_AGEMA_signal_18781 ;
    wire new_AGEMA_signal_18782 ;
    wire new_AGEMA_signal_18783 ;
    wire new_AGEMA_signal_18784 ;
    wire new_AGEMA_signal_18785 ;
    wire new_AGEMA_signal_18786 ;
    wire new_AGEMA_signal_18787 ;
    wire new_AGEMA_signal_18788 ;
    wire new_AGEMA_signal_18789 ;
    wire new_AGEMA_signal_18790 ;
    wire new_AGEMA_signal_18791 ;
    wire new_AGEMA_signal_18792 ;
    wire new_AGEMA_signal_18793 ;
    wire new_AGEMA_signal_18794 ;
    wire new_AGEMA_signal_18795 ;
    wire new_AGEMA_signal_18796 ;
    wire new_AGEMA_signal_18797 ;
    wire new_AGEMA_signal_18798 ;
    wire new_AGEMA_signal_18799 ;
    wire new_AGEMA_signal_18800 ;
    wire new_AGEMA_signal_18801 ;
    wire new_AGEMA_signal_18802 ;
    wire new_AGEMA_signal_18803 ;
    wire new_AGEMA_signal_18804 ;
    wire new_AGEMA_signal_18805 ;
    wire new_AGEMA_signal_18806 ;
    wire new_AGEMA_signal_18807 ;
    wire new_AGEMA_signal_18808 ;
    wire new_AGEMA_signal_18809 ;
    wire new_AGEMA_signal_18810 ;
    wire new_AGEMA_signal_18811 ;
    wire new_AGEMA_signal_18812 ;
    wire new_AGEMA_signal_18813 ;
    wire new_AGEMA_signal_18814 ;
    wire new_AGEMA_signal_18815 ;
    wire new_AGEMA_signal_18816 ;
    wire new_AGEMA_signal_18817 ;
    wire new_AGEMA_signal_18818 ;
    wire new_AGEMA_signal_18819 ;
    wire new_AGEMA_signal_18820 ;
    wire new_AGEMA_signal_18821 ;
    wire new_AGEMA_signal_18822 ;
    wire new_AGEMA_signal_18823 ;
    wire new_AGEMA_signal_18824 ;
    wire new_AGEMA_signal_18825 ;
    wire new_AGEMA_signal_18826 ;
    wire new_AGEMA_signal_18827 ;
    wire new_AGEMA_signal_18828 ;
    wire new_AGEMA_signal_18829 ;
    wire new_AGEMA_signal_18830 ;
    wire new_AGEMA_signal_18831 ;
    wire new_AGEMA_signal_18832 ;
    wire new_AGEMA_signal_18833 ;
    wire new_AGEMA_signal_18834 ;
    wire new_AGEMA_signal_18835 ;
    wire new_AGEMA_signal_18836 ;
    wire new_AGEMA_signal_18837 ;
    wire new_AGEMA_signal_18838 ;
    wire new_AGEMA_signal_18839 ;
    wire new_AGEMA_signal_18840 ;
    wire new_AGEMA_signal_18841 ;
    wire new_AGEMA_signal_18842 ;
    wire new_AGEMA_signal_18843 ;
    wire new_AGEMA_signal_18844 ;
    wire new_AGEMA_signal_18845 ;
    wire new_AGEMA_signal_18846 ;
    wire new_AGEMA_signal_18847 ;
    wire new_AGEMA_signal_18848 ;
    wire new_AGEMA_signal_18849 ;
    wire new_AGEMA_signal_18850 ;
    wire new_AGEMA_signal_18851 ;
    wire new_AGEMA_signal_18852 ;
    wire new_AGEMA_signal_18853 ;
    wire new_AGEMA_signal_18854 ;
    wire new_AGEMA_signal_18855 ;
    wire new_AGEMA_signal_18856 ;
    wire new_AGEMA_signal_18857 ;
    wire new_AGEMA_signal_18858 ;
    wire new_AGEMA_signal_18859 ;
    wire new_AGEMA_signal_18860 ;
    wire new_AGEMA_signal_18861 ;
    wire new_AGEMA_signal_18862 ;
    wire new_AGEMA_signal_18863 ;
    wire new_AGEMA_signal_18864 ;
    wire new_AGEMA_signal_18865 ;
    wire new_AGEMA_signal_18866 ;
    wire new_AGEMA_signal_18867 ;
    wire new_AGEMA_signal_18868 ;
    wire new_AGEMA_signal_18869 ;
    wire new_AGEMA_signal_18870 ;
    wire new_AGEMA_signal_18871 ;
    wire new_AGEMA_signal_18872 ;
    wire new_AGEMA_signal_18873 ;
    wire new_AGEMA_signal_18874 ;
    wire new_AGEMA_signal_18875 ;
    wire new_AGEMA_signal_18876 ;
    wire new_AGEMA_signal_18877 ;
    wire new_AGEMA_signal_18878 ;
    wire new_AGEMA_signal_18879 ;
    wire new_AGEMA_signal_18880 ;
    wire new_AGEMA_signal_18881 ;
    wire new_AGEMA_signal_18882 ;
    wire new_AGEMA_signal_18883 ;
    wire new_AGEMA_signal_18884 ;
    wire new_AGEMA_signal_18885 ;
    wire new_AGEMA_signal_18886 ;
    wire new_AGEMA_signal_18887 ;
    wire new_AGEMA_signal_18888 ;
    wire new_AGEMA_signal_18889 ;
    wire new_AGEMA_signal_18890 ;
    wire new_AGEMA_signal_18891 ;
    wire new_AGEMA_signal_18892 ;
    wire new_AGEMA_signal_18893 ;
    wire new_AGEMA_signal_18894 ;
    wire new_AGEMA_signal_18895 ;
    wire new_AGEMA_signal_18896 ;
    wire new_AGEMA_signal_18897 ;
    wire new_AGEMA_signal_18898 ;
    wire new_AGEMA_signal_18899 ;
    wire new_AGEMA_signal_18900 ;
    wire new_AGEMA_signal_18901 ;
    wire new_AGEMA_signal_18902 ;
    wire new_AGEMA_signal_18903 ;
    wire new_AGEMA_signal_18904 ;
    wire new_AGEMA_signal_18905 ;
    wire new_AGEMA_signal_18906 ;
    wire new_AGEMA_signal_18907 ;
    wire new_AGEMA_signal_18908 ;
    wire new_AGEMA_signal_18909 ;
    wire new_AGEMA_signal_18910 ;
    wire new_AGEMA_signal_18911 ;
    wire new_AGEMA_signal_18912 ;
    wire new_AGEMA_signal_18913 ;
    wire new_AGEMA_signal_18914 ;
    wire new_AGEMA_signal_18915 ;
    wire new_AGEMA_signal_18916 ;
    wire new_AGEMA_signal_18917 ;
    wire new_AGEMA_signal_18918 ;
    wire new_AGEMA_signal_18919 ;
    wire new_AGEMA_signal_18920 ;
    wire new_AGEMA_signal_18921 ;
    wire new_AGEMA_signal_18922 ;
    wire new_AGEMA_signal_18923 ;
    wire new_AGEMA_signal_18924 ;
    wire new_AGEMA_signal_18925 ;
    wire new_AGEMA_signal_18926 ;
    wire new_AGEMA_signal_18927 ;
    wire new_AGEMA_signal_18928 ;
    wire new_AGEMA_signal_18929 ;
    wire new_AGEMA_signal_18930 ;
    wire new_AGEMA_signal_18931 ;
    wire new_AGEMA_signal_18932 ;
    wire new_AGEMA_signal_18933 ;
    wire new_AGEMA_signal_18934 ;
    wire new_AGEMA_signal_18935 ;
    wire new_AGEMA_signal_18936 ;
    wire new_AGEMA_signal_18937 ;
    wire new_AGEMA_signal_18938 ;
    wire new_AGEMA_signal_18939 ;
    wire new_AGEMA_signal_18940 ;
    wire new_AGEMA_signal_18941 ;
    wire new_AGEMA_signal_18942 ;
    wire new_AGEMA_signal_18943 ;
    wire new_AGEMA_signal_18944 ;
    wire new_AGEMA_signal_18945 ;
    wire new_AGEMA_signal_18946 ;
    wire new_AGEMA_signal_18947 ;
    wire new_AGEMA_signal_18948 ;
    wire new_AGEMA_signal_18949 ;
    wire new_AGEMA_signal_18950 ;
    wire new_AGEMA_signal_18951 ;
    wire new_AGEMA_signal_18952 ;
    wire new_AGEMA_signal_18953 ;
    wire new_AGEMA_signal_18954 ;
    wire new_AGEMA_signal_18955 ;
    wire new_AGEMA_signal_18956 ;
    wire new_AGEMA_signal_18957 ;
    wire new_AGEMA_signal_18958 ;
    wire new_AGEMA_signal_18959 ;
    wire new_AGEMA_signal_18960 ;
    wire new_AGEMA_signal_18961 ;
    wire new_AGEMA_signal_18962 ;
    wire new_AGEMA_signal_18963 ;
    wire new_AGEMA_signal_18964 ;
    wire new_AGEMA_signal_18965 ;
    wire new_AGEMA_signal_18966 ;
    wire new_AGEMA_signal_18967 ;
    wire new_AGEMA_signal_18968 ;
    wire new_AGEMA_signal_18969 ;
    wire new_AGEMA_signal_18970 ;
    wire new_AGEMA_signal_18971 ;
    wire new_AGEMA_signal_18972 ;
    wire new_AGEMA_signal_18973 ;
    wire new_AGEMA_signal_18974 ;
    wire new_AGEMA_signal_18975 ;
    wire new_AGEMA_signal_18976 ;
    wire new_AGEMA_signal_18977 ;
    wire new_AGEMA_signal_18978 ;
    wire new_AGEMA_signal_18979 ;
    wire new_AGEMA_signal_18980 ;
    wire new_AGEMA_signal_18981 ;
    wire new_AGEMA_signal_18982 ;
    wire new_AGEMA_signal_18983 ;
    wire new_AGEMA_signal_18984 ;
    wire new_AGEMA_signal_18985 ;
    wire new_AGEMA_signal_18986 ;
    wire new_AGEMA_signal_18987 ;
    wire new_AGEMA_signal_18988 ;
    wire new_AGEMA_signal_18989 ;
    wire new_AGEMA_signal_18990 ;
    wire new_AGEMA_signal_18991 ;
    wire new_AGEMA_signal_18992 ;
    wire new_AGEMA_signal_18993 ;
    wire new_AGEMA_signal_18994 ;
    wire new_AGEMA_signal_18995 ;
    wire new_AGEMA_signal_18996 ;
    wire new_AGEMA_signal_18997 ;
    wire new_AGEMA_signal_18998 ;
    wire new_AGEMA_signal_18999 ;
    wire new_AGEMA_signal_19000 ;
    wire new_AGEMA_signal_19001 ;
    wire new_AGEMA_signal_19002 ;
    wire new_AGEMA_signal_19003 ;
    wire new_AGEMA_signal_19004 ;
    wire new_AGEMA_signal_19005 ;
    wire new_AGEMA_signal_19006 ;
    wire new_AGEMA_signal_19007 ;
    wire new_AGEMA_signal_19008 ;
    wire new_AGEMA_signal_19009 ;
    wire new_AGEMA_signal_19010 ;
    wire new_AGEMA_signal_19011 ;
    wire new_AGEMA_signal_19012 ;
    wire new_AGEMA_signal_19013 ;
    wire new_AGEMA_signal_19014 ;
    wire new_AGEMA_signal_19015 ;
    wire new_AGEMA_signal_19016 ;
    wire new_AGEMA_signal_19017 ;
    wire new_AGEMA_signal_19018 ;
    wire new_AGEMA_signal_19019 ;
    wire new_AGEMA_signal_19020 ;
    wire new_AGEMA_signal_19021 ;
    wire new_AGEMA_signal_19022 ;
    wire new_AGEMA_signal_19023 ;
    wire new_AGEMA_signal_19024 ;
    wire new_AGEMA_signal_19025 ;
    wire new_AGEMA_signal_19026 ;
    wire new_AGEMA_signal_19027 ;
    wire new_AGEMA_signal_19028 ;
    wire new_AGEMA_signal_19029 ;
    wire new_AGEMA_signal_19030 ;
    wire new_AGEMA_signal_19031 ;
    wire new_AGEMA_signal_19032 ;
    wire new_AGEMA_signal_19033 ;
    wire new_AGEMA_signal_19034 ;
    wire new_AGEMA_signal_19035 ;
    wire new_AGEMA_signal_19036 ;
    wire new_AGEMA_signal_19037 ;
    wire new_AGEMA_signal_19038 ;
    wire new_AGEMA_signal_19039 ;
    wire new_AGEMA_signal_19040 ;
    wire new_AGEMA_signal_19041 ;
    wire new_AGEMA_signal_19042 ;
    wire new_AGEMA_signal_19043 ;
    wire new_AGEMA_signal_19044 ;
    wire new_AGEMA_signal_19045 ;
    wire new_AGEMA_signal_19046 ;
    wire new_AGEMA_signal_19047 ;
    wire new_AGEMA_signal_19048 ;
    wire new_AGEMA_signal_19049 ;
    wire new_AGEMA_signal_19050 ;
    wire new_AGEMA_signal_19051 ;
    wire new_AGEMA_signal_19052 ;
    wire new_AGEMA_signal_19053 ;
    wire new_AGEMA_signal_19054 ;
    wire new_AGEMA_signal_19055 ;
    wire new_AGEMA_signal_19056 ;
    wire new_AGEMA_signal_19057 ;
    wire new_AGEMA_signal_19058 ;
    wire new_AGEMA_signal_19059 ;
    wire new_AGEMA_signal_19060 ;
    wire new_AGEMA_signal_19061 ;
    wire new_AGEMA_signal_19062 ;
    wire new_AGEMA_signal_19063 ;
    wire new_AGEMA_signal_19064 ;
    wire new_AGEMA_signal_19065 ;
    wire new_AGEMA_signal_19066 ;
    wire new_AGEMA_signal_19067 ;
    wire new_AGEMA_signal_19068 ;
    wire new_AGEMA_signal_19069 ;
    wire new_AGEMA_signal_19070 ;
    wire new_AGEMA_signal_19071 ;
    wire new_AGEMA_signal_19072 ;
    wire new_AGEMA_signal_19073 ;
    wire new_AGEMA_signal_19074 ;
    wire new_AGEMA_signal_19075 ;
    wire new_AGEMA_signal_19076 ;
    wire new_AGEMA_signal_19077 ;
    wire new_AGEMA_signal_19078 ;
    wire new_AGEMA_signal_19079 ;
    wire new_AGEMA_signal_19080 ;
    wire new_AGEMA_signal_19081 ;
    wire new_AGEMA_signal_19082 ;
    wire new_AGEMA_signal_19083 ;
    wire new_AGEMA_signal_19084 ;
    wire new_AGEMA_signal_19085 ;
    wire new_AGEMA_signal_19086 ;
    wire new_AGEMA_signal_19087 ;
    wire new_AGEMA_signal_19088 ;
    wire new_AGEMA_signal_19089 ;
    wire new_AGEMA_signal_19090 ;
    wire new_AGEMA_signal_19091 ;
    wire new_AGEMA_signal_19092 ;
    wire new_AGEMA_signal_19093 ;
    wire new_AGEMA_signal_19094 ;
    wire new_AGEMA_signal_19095 ;
    wire new_AGEMA_signal_19096 ;
    wire new_AGEMA_signal_19097 ;
    wire new_AGEMA_signal_19098 ;
    wire new_AGEMA_signal_19099 ;
    wire new_AGEMA_signal_19100 ;
    wire new_AGEMA_signal_19101 ;
    wire new_AGEMA_signal_19102 ;
    wire new_AGEMA_signal_19103 ;
    wire new_AGEMA_signal_19104 ;
    wire new_AGEMA_signal_19105 ;
    wire new_AGEMA_signal_19106 ;
    wire new_AGEMA_signal_19107 ;
    wire new_AGEMA_signal_19108 ;
    wire new_AGEMA_signal_19109 ;
    wire new_AGEMA_signal_19110 ;
    wire new_AGEMA_signal_19111 ;
    wire new_AGEMA_signal_19112 ;
    wire new_AGEMA_signal_19113 ;
    wire new_AGEMA_signal_19114 ;
    wire new_AGEMA_signal_19115 ;
    wire new_AGEMA_signal_19116 ;
    wire new_AGEMA_signal_19117 ;
    wire new_AGEMA_signal_19118 ;
    wire new_AGEMA_signal_19119 ;
    wire new_AGEMA_signal_19120 ;
    wire new_AGEMA_signal_19121 ;
    wire new_AGEMA_signal_19122 ;
    wire new_AGEMA_signal_19123 ;
    wire new_AGEMA_signal_19124 ;
    wire new_AGEMA_signal_19125 ;
    wire new_AGEMA_signal_19126 ;
    wire new_AGEMA_signal_19127 ;
    wire new_AGEMA_signal_19128 ;
    wire new_AGEMA_signal_19129 ;
    wire new_AGEMA_signal_19130 ;
    wire new_AGEMA_signal_19131 ;
    wire new_AGEMA_signal_19132 ;
    wire new_AGEMA_signal_19133 ;
    wire new_AGEMA_signal_19134 ;
    wire new_AGEMA_signal_19135 ;
    wire new_AGEMA_signal_19136 ;
    wire new_AGEMA_signal_19137 ;
    wire new_AGEMA_signal_19138 ;
    wire new_AGEMA_signal_19139 ;
    wire new_AGEMA_signal_19140 ;
    wire new_AGEMA_signal_19141 ;
    wire new_AGEMA_signal_19142 ;
    wire new_AGEMA_signal_19143 ;
    wire new_AGEMA_signal_19144 ;
    wire new_AGEMA_signal_19145 ;
    wire new_AGEMA_signal_19146 ;
    wire new_AGEMA_signal_19147 ;
    wire new_AGEMA_signal_19148 ;
    wire new_AGEMA_signal_19149 ;
    wire new_AGEMA_signal_19150 ;
    wire new_AGEMA_signal_19151 ;
    wire new_AGEMA_signal_19152 ;
    wire new_AGEMA_signal_19153 ;
    wire new_AGEMA_signal_19154 ;
    wire new_AGEMA_signal_19155 ;
    wire new_AGEMA_signal_19156 ;
    wire new_AGEMA_signal_19157 ;
    wire new_AGEMA_signal_19158 ;
    wire new_AGEMA_signal_19159 ;
    wire new_AGEMA_signal_19160 ;
    wire new_AGEMA_signal_19161 ;
    wire new_AGEMA_signal_19162 ;
    wire new_AGEMA_signal_19163 ;
    wire new_AGEMA_signal_19164 ;
    wire new_AGEMA_signal_19165 ;
    wire new_AGEMA_signal_19166 ;
    wire new_AGEMA_signal_19167 ;
    wire new_AGEMA_signal_19168 ;
    wire new_AGEMA_signal_19169 ;
    wire new_AGEMA_signal_19170 ;
    wire new_AGEMA_signal_19171 ;
    wire new_AGEMA_signal_19172 ;
    wire new_AGEMA_signal_19173 ;
    wire new_AGEMA_signal_19174 ;
    wire new_AGEMA_signal_19175 ;
    wire new_AGEMA_signal_19176 ;
    wire new_AGEMA_signal_19177 ;
    wire new_AGEMA_signal_19178 ;
    wire new_AGEMA_signal_19179 ;
    wire new_AGEMA_signal_19180 ;
    wire new_AGEMA_signal_19181 ;
    wire new_AGEMA_signal_19182 ;
    wire new_AGEMA_signal_19183 ;
    wire new_AGEMA_signal_19184 ;
    wire new_AGEMA_signal_19185 ;
    wire new_AGEMA_signal_19186 ;
    wire new_AGEMA_signal_19187 ;
    wire new_AGEMA_signal_19188 ;
    wire new_AGEMA_signal_19189 ;
    wire new_AGEMA_signal_19190 ;
    wire new_AGEMA_signal_19191 ;
    wire new_AGEMA_signal_19192 ;
    wire new_AGEMA_signal_19193 ;
    wire new_AGEMA_signal_19194 ;
    wire new_AGEMA_signal_19195 ;
    wire new_AGEMA_signal_19196 ;
    wire new_AGEMA_signal_19197 ;
    wire new_AGEMA_signal_19198 ;
    wire new_AGEMA_signal_19199 ;
    wire new_AGEMA_signal_19200 ;
    wire new_AGEMA_signal_19201 ;
    wire new_AGEMA_signal_19202 ;
    wire new_AGEMA_signal_19203 ;
    wire new_AGEMA_signal_19204 ;
    wire new_AGEMA_signal_19205 ;
    wire new_AGEMA_signal_19206 ;
    wire new_AGEMA_signal_19207 ;
    wire new_AGEMA_signal_19208 ;
    wire new_AGEMA_signal_19209 ;
    wire new_AGEMA_signal_19210 ;
    wire new_AGEMA_signal_19211 ;
    wire new_AGEMA_signal_19212 ;
    wire new_AGEMA_signal_19213 ;
    wire new_AGEMA_signal_19214 ;
    wire new_AGEMA_signal_19215 ;
    wire new_AGEMA_signal_19216 ;
    wire new_AGEMA_signal_19217 ;
    wire new_AGEMA_signal_19218 ;
    wire new_AGEMA_signal_19219 ;
    wire new_AGEMA_signal_19220 ;
    wire new_AGEMA_signal_19221 ;
    wire new_AGEMA_signal_19222 ;
    wire new_AGEMA_signal_19223 ;
    wire new_AGEMA_signal_19224 ;
    wire new_AGEMA_signal_19225 ;
    wire new_AGEMA_signal_19226 ;
    wire new_AGEMA_signal_19227 ;
    wire new_AGEMA_signal_19228 ;
    wire new_AGEMA_signal_19229 ;
    wire new_AGEMA_signal_19230 ;
    wire new_AGEMA_signal_19231 ;
    wire new_AGEMA_signal_19232 ;
    wire new_AGEMA_signal_19233 ;
    wire new_AGEMA_signal_19234 ;
    wire new_AGEMA_signal_19235 ;
    wire new_AGEMA_signal_19236 ;
    wire new_AGEMA_signal_19237 ;
    wire new_AGEMA_signal_19238 ;
    wire new_AGEMA_signal_19239 ;
    wire new_AGEMA_signal_19240 ;
    wire new_AGEMA_signal_19241 ;
    wire new_AGEMA_signal_19242 ;
    wire new_AGEMA_signal_19243 ;
    wire new_AGEMA_signal_19244 ;
    wire new_AGEMA_signal_19245 ;
    wire new_AGEMA_signal_19246 ;
    wire new_AGEMA_signal_19247 ;
    wire new_AGEMA_signal_19248 ;
    wire new_AGEMA_signal_19249 ;
    wire new_AGEMA_signal_19250 ;
    wire new_AGEMA_signal_19251 ;
    wire new_AGEMA_signal_19252 ;
    wire new_AGEMA_signal_19253 ;
    wire new_AGEMA_signal_19254 ;
    wire new_AGEMA_signal_19255 ;
    wire new_AGEMA_signal_19256 ;
    wire new_AGEMA_signal_19257 ;
    wire new_AGEMA_signal_19258 ;
    wire new_AGEMA_signal_19259 ;
    wire new_AGEMA_signal_19260 ;
    wire new_AGEMA_signal_19261 ;
    wire new_AGEMA_signal_19262 ;
    wire new_AGEMA_signal_19263 ;
    wire new_AGEMA_signal_19264 ;
    wire new_AGEMA_signal_19265 ;
    wire new_AGEMA_signal_19266 ;
    wire new_AGEMA_signal_19267 ;
    wire new_AGEMA_signal_19268 ;
    wire new_AGEMA_signal_19269 ;
    wire new_AGEMA_signal_19270 ;
    wire new_AGEMA_signal_19271 ;
    wire new_AGEMA_signal_19272 ;
    wire new_AGEMA_signal_19273 ;
    wire new_AGEMA_signal_19274 ;
    wire new_AGEMA_signal_19275 ;
    wire new_AGEMA_signal_19276 ;
    wire new_AGEMA_signal_19277 ;
    wire new_AGEMA_signal_19278 ;
    wire new_AGEMA_signal_19279 ;
    wire new_AGEMA_signal_19280 ;
    wire new_AGEMA_signal_19281 ;
    wire new_AGEMA_signal_19282 ;
    wire new_AGEMA_signal_19283 ;
    wire new_AGEMA_signal_19284 ;
    wire new_AGEMA_signal_19285 ;
    wire new_AGEMA_signal_19286 ;
    wire new_AGEMA_signal_19287 ;
    wire new_AGEMA_signal_19288 ;
    wire new_AGEMA_signal_19289 ;
    wire new_AGEMA_signal_19290 ;
    wire new_AGEMA_signal_19291 ;
    wire new_AGEMA_signal_19292 ;
    wire new_AGEMA_signal_19293 ;
    wire new_AGEMA_signal_19294 ;
    wire new_AGEMA_signal_19295 ;
    wire new_AGEMA_signal_19296 ;
    wire new_AGEMA_signal_19297 ;
    wire new_AGEMA_signal_19298 ;
    wire new_AGEMA_signal_19299 ;
    wire new_AGEMA_signal_19300 ;
    wire new_AGEMA_signal_19301 ;
    wire new_AGEMA_signal_19302 ;
    wire new_AGEMA_signal_19303 ;
    wire new_AGEMA_signal_19304 ;
    wire new_AGEMA_signal_19305 ;
    wire new_AGEMA_signal_19306 ;
    wire new_AGEMA_signal_19307 ;
    wire new_AGEMA_signal_19308 ;
    wire new_AGEMA_signal_19309 ;
    wire new_AGEMA_signal_19310 ;
    wire new_AGEMA_signal_19311 ;
    wire new_AGEMA_signal_19312 ;
    wire new_AGEMA_signal_19313 ;
    wire new_AGEMA_signal_19314 ;
    wire new_AGEMA_signal_19315 ;
    wire new_AGEMA_signal_19316 ;
    wire new_AGEMA_signal_19317 ;
    wire new_AGEMA_signal_19318 ;
    wire new_AGEMA_signal_19319 ;
    wire new_AGEMA_signal_19320 ;
    wire new_AGEMA_signal_19321 ;
    wire new_AGEMA_signal_19322 ;
    wire new_AGEMA_signal_19323 ;
    wire new_AGEMA_signal_19324 ;
    wire new_AGEMA_signal_19325 ;
    wire new_AGEMA_signal_19326 ;
    wire new_AGEMA_signal_19327 ;
    wire new_AGEMA_signal_19328 ;
    wire new_AGEMA_signal_19329 ;
    wire new_AGEMA_signal_19330 ;
    wire new_AGEMA_signal_19331 ;
    wire new_AGEMA_signal_19332 ;
    wire new_AGEMA_signal_19333 ;
    wire new_AGEMA_signal_19334 ;
    wire new_AGEMA_signal_19335 ;
    wire new_AGEMA_signal_19336 ;
    wire new_AGEMA_signal_19337 ;
    wire new_AGEMA_signal_19338 ;
    wire new_AGEMA_signal_19339 ;
    wire new_AGEMA_signal_19340 ;
    wire new_AGEMA_signal_19341 ;
    wire new_AGEMA_signal_19342 ;
    wire new_AGEMA_signal_19343 ;
    wire new_AGEMA_signal_19344 ;
    wire new_AGEMA_signal_19345 ;
    wire new_AGEMA_signal_19346 ;
    wire new_AGEMA_signal_19347 ;
    wire new_AGEMA_signal_19348 ;
    wire new_AGEMA_signal_19349 ;
    wire new_AGEMA_signal_19350 ;
    wire new_AGEMA_signal_19351 ;
    wire new_AGEMA_signal_19352 ;
    wire new_AGEMA_signal_19353 ;
    wire new_AGEMA_signal_19354 ;
    wire new_AGEMA_signal_19355 ;
    wire new_AGEMA_signal_19356 ;
    wire new_AGEMA_signal_19357 ;
    wire new_AGEMA_signal_19358 ;
    wire new_AGEMA_signal_19359 ;
    wire new_AGEMA_signal_19360 ;
    wire new_AGEMA_signal_19361 ;
    wire new_AGEMA_signal_19362 ;
    wire new_AGEMA_signal_19363 ;
    wire new_AGEMA_signal_19364 ;
    wire new_AGEMA_signal_19365 ;
    wire new_AGEMA_signal_19366 ;
    wire new_AGEMA_signal_19367 ;
    wire new_AGEMA_signal_19368 ;
    wire new_AGEMA_signal_19369 ;
    wire new_AGEMA_signal_19370 ;
    wire new_AGEMA_signal_19371 ;
    wire new_AGEMA_signal_19372 ;
    wire new_AGEMA_signal_19373 ;
    wire new_AGEMA_signal_19374 ;
    wire new_AGEMA_signal_19375 ;
    wire new_AGEMA_signal_19376 ;
    wire new_AGEMA_signal_19377 ;
    wire new_AGEMA_signal_19378 ;
    wire new_AGEMA_signal_19379 ;
    wire new_AGEMA_signal_19380 ;
    wire new_AGEMA_signal_19381 ;
    wire new_AGEMA_signal_19382 ;
    wire new_AGEMA_signal_19383 ;
    wire new_AGEMA_signal_19384 ;
    wire new_AGEMA_signal_19385 ;
    wire new_AGEMA_signal_19386 ;
    wire new_AGEMA_signal_19387 ;
    wire new_AGEMA_signal_19388 ;
    wire new_AGEMA_signal_19389 ;
    wire new_AGEMA_signal_19390 ;
    wire new_AGEMA_signal_19391 ;
    wire new_AGEMA_signal_19392 ;
    wire new_AGEMA_signal_19393 ;
    wire new_AGEMA_signal_19394 ;
    wire new_AGEMA_signal_19395 ;
    wire new_AGEMA_signal_19396 ;
    wire new_AGEMA_signal_19397 ;
    wire new_AGEMA_signal_19398 ;
    wire new_AGEMA_signal_19399 ;
    wire new_AGEMA_signal_19400 ;
    wire new_AGEMA_signal_19401 ;
    wire new_AGEMA_signal_19402 ;
    wire new_AGEMA_signal_19403 ;
    wire new_AGEMA_signal_19404 ;
    wire new_AGEMA_signal_19405 ;
    wire new_AGEMA_signal_19406 ;
    wire new_AGEMA_signal_19407 ;
    wire new_AGEMA_signal_19408 ;
    wire new_AGEMA_signal_19409 ;
    wire new_AGEMA_signal_19410 ;
    wire new_AGEMA_signal_19411 ;
    wire new_AGEMA_signal_19412 ;
    wire new_AGEMA_signal_19413 ;
    wire new_AGEMA_signal_19414 ;
    wire new_AGEMA_signal_19415 ;
    wire new_AGEMA_signal_19416 ;
    wire new_AGEMA_signal_19417 ;
    wire new_AGEMA_signal_19418 ;
    wire new_AGEMA_signal_19419 ;
    wire new_AGEMA_signal_19420 ;
    wire new_AGEMA_signal_19421 ;
    wire new_AGEMA_signal_19422 ;
    wire new_AGEMA_signal_19423 ;
    wire new_AGEMA_signal_19424 ;
    wire new_AGEMA_signal_19425 ;
    wire new_AGEMA_signal_19426 ;
    wire new_AGEMA_signal_19427 ;
    wire new_AGEMA_signal_19428 ;
    wire new_AGEMA_signal_19429 ;
    wire new_AGEMA_signal_19430 ;
    wire new_AGEMA_signal_19431 ;
    wire new_AGEMA_signal_19432 ;
    wire new_AGEMA_signal_19433 ;
    wire new_AGEMA_signal_19434 ;
    wire new_AGEMA_signal_19435 ;
    wire new_AGEMA_signal_19436 ;
    wire new_AGEMA_signal_19437 ;
    wire new_AGEMA_signal_19438 ;
    wire new_AGEMA_signal_19439 ;
    wire new_AGEMA_signal_19440 ;
    wire new_AGEMA_signal_19441 ;
    wire new_AGEMA_signal_19442 ;
    wire new_AGEMA_signal_19443 ;
    wire new_AGEMA_signal_19444 ;
    wire new_AGEMA_signal_19445 ;
    wire new_AGEMA_signal_19446 ;
    wire new_AGEMA_signal_19447 ;
    wire new_AGEMA_signal_19448 ;
    wire new_AGEMA_signal_19449 ;
    wire new_AGEMA_signal_19450 ;
    wire new_AGEMA_signal_19451 ;
    wire new_AGEMA_signal_19452 ;
    wire new_AGEMA_signal_19453 ;
    wire new_AGEMA_signal_19454 ;
    wire new_AGEMA_signal_19455 ;
    wire new_AGEMA_signal_19456 ;
    wire new_AGEMA_signal_19457 ;
    wire new_AGEMA_signal_19458 ;
    wire new_AGEMA_signal_19459 ;
    wire new_AGEMA_signal_19460 ;
    wire new_AGEMA_signal_19461 ;
    wire new_AGEMA_signal_19462 ;
    wire new_AGEMA_signal_19463 ;
    wire new_AGEMA_signal_19464 ;
    wire new_AGEMA_signal_19465 ;
    wire new_AGEMA_signal_19466 ;
    wire new_AGEMA_signal_19467 ;
    wire new_AGEMA_signal_19468 ;
    wire new_AGEMA_signal_19469 ;
    wire new_AGEMA_signal_19470 ;
    wire new_AGEMA_signal_19471 ;
    wire new_AGEMA_signal_19472 ;
    wire new_AGEMA_signal_19473 ;
    wire new_AGEMA_signal_19474 ;
    wire new_AGEMA_signal_19475 ;
    wire new_AGEMA_signal_19476 ;
    wire new_AGEMA_signal_19477 ;
    wire new_AGEMA_signal_19478 ;
    wire new_AGEMA_signal_19479 ;
    wire new_AGEMA_signal_19480 ;
    wire new_AGEMA_signal_19481 ;
    wire new_AGEMA_signal_19482 ;
    wire new_AGEMA_signal_19483 ;
    wire new_AGEMA_signal_19484 ;
    wire new_AGEMA_signal_19485 ;
    wire new_AGEMA_signal_19486 ;
    wire new_AGEMA_signal_19487 ;
    wire new_AGEMA_signal_19488 ;
    wire new_AGEMA_signal_19489 ;
    wire new_AGEMA_signal_19490 ;
    wire new_AGEMA_signal_19491 ;
    wire new_AGEMA_signal_19492 ;
    wire new_AGEMA_signal_19493 ;
    wire new_AGEMA_signal_19494 ;
    wire new_AGEMA_signal_19495 ;
    wire new_AGEMA_signal_19496 ;
    wire new_AGEMA_signal_19497 ;
    wire new_AGEMA_signal_19498 ;
    wire new_AGEMA_signal_19499 ;
    wire new_AGEMA_signal_19500 ;
    wire new_AGEMA_signal_19501 ;
    wire new_AGEMA_signal_19502 ;
    wire new_AGEMA_signal_19503 ;
    wire new_AGEMA_signal_19504 ;
    wire new_AGEMA_signal_19505 ;
    wire new_AGEMA_signal_19506 ;
    wire new_AGEMA_signal_19507 ;
    wire new_AGEMA_signal_19508 ;
    wire new_AGEMA_signal_19509 ;
    wire new_AGEMA_signal_19510 ;
    wire new_AGEMA_signal_19511 ;
    wire new_AGEMA_signal_19512 ;
    wire new_AGEMA_signal_19513 ;
    wire new_AGEMA_signal_19514 ;
    wire new_AGEMA_signal_19515 ;
    wire new_AGEMA_signal_19516 ;
    wire new_AGEMA_signal_19517 ;
    wire new_AGEMA_signal_19518 ;
    wire new_AGEMA_signal_19519 ;
    wire new_AGEMA_signal_19520 ;
    wire new_AGEMA_signal_19521 ;
    wire new_AGEMA_signal_19522 ;
    wire new_AGEMA_signal_19523 ;
    wire new_AGEMA_signal_19524 ;
    wire new_AGEMA_signal_19525 ;
    wire new_AGEMA_signal_19526 ;
    wire new_AGEMA_signal_19527 ;
    wire new_AGEMA_signal_19528 ;
    wire new_AGEMA_signal_19529 ;
    wire new_AGEMA_signal_19530 ;
    wire new_AGEMA_signal_19531 ;
    wire new_AGEMA_signal_19532 ;
    wire new_AGEMA_signal_19533 ;
    wire new_AGEMA_signal_19534 ;
    wire new_AGEMA_signal_19535 ;
    wire new_AGEMA_signal_19536 ;
    wire new_AGEMA_signal_19537 ;
    wire new_AGEMA_signal_19538 ;
    wire new_AGEMA_signal_19539 ;
    wire new_AGEMA_signal_19540 ;
    wire new_AGEMA_signal_19541 ;
    wire new_AGEMA_signal_19542 ;
    wire new_AGEMA_signal_19543 ;
    wire new_AGEMA_signal_19544 ;
    wire new_AGEMA_signal_19545 ;
    wire new_AGEMA_signal_19546 ;
    wire new_AGEMA_signal_19547 ;
    wire new_AGEMA_signal_19548 ;
    wire new_AGEMA_signal_19549 ;
    wire new_AGEMA_signal_19550 ;
    wire new_AGEMA_signal_19551 ;
    wire new_AGEMA_signal_19552 ;
    wire new_AGEMA_signal_19553 ;
    wire new_AGEMA_signal_19554 ;
    wire new_AGEMA_signal_19555 ;
    wire new_AGEMA_signal_19556 ;
    wire new_AGEMA_signal_19557 ;
    wire new_AGEMA_signal_19558 ;
    wire new_AGEMA_signal_19559 ;
    wire new_AGEMA_signal_19560 ;
    wire new_AGEMA_signal_19561 ;
    wire new_AGEMA_signal_19562 ;
    wire new_AGEMA_signal_19563 ;
    wire new_AGEMA_signal_19564 ;
    wire new_AGEMA_signal_19565 ;
    wire new_AGEMA_signal_19566 ;
    wire new_AGEMA_signal_19567 ;
    wire new_AGEMA_signal_19568 ;
    wire new_AGEMA_signal_19569 ;
    wire new_AGEMA_signal_19570 ;
    wire new_AGEMA_signal_19571 ;
    wire new_AGEMA_signal_19572 ;
    wire new_AGEMA_signal_19573 ;
    wire new_AGEMA_signal_19574 ;
    wire new_AGEMA_signal_19575 ;
    wire new_AGEMA_signal_19576 ;
    wire new_AGEMA_signal_19577 ;
    wire new_AGEMA_signal_19578 ;
    wire new_AGEMA_signal_19579 ;
    wire new_AGEMA_signal_19580 ;
    wire new_AGEMA_signal_19581 ;
    wire new_AGEMA_signal_19582 ;
    wire new_AGEMA_signal_19583 ;
    wire new_AGEMA_signal_19584 ;
    wire new_AGEMA_signal_19585 ;
    wire new_AGEMA_signal_19586 ;
    wire new_AGEMA_signal_19587 ;
    wire new_AGEMA_signal_19588 ;
    wire new_AGEMA_signal_19589 ;
    wire new_AGEMA_signal_19590 ;
    wire new_AGEMA_signal_19591 ;
    wire new_AGEMA_signal_19592 ;
    wire new_AGEMA_signal_19593 ;
    wire new_AGEMA_signal_19594 ;
    wire new_AGEMA_signal_19595 ;
    wire new_AGEMA_signal_19596 ;
    wire new_AGEMA_signal_19597 ;
    wire new_AGEMA_signal_19598 ;
    wire new_AGEMA_signal_19599 ;
    wire new_AGEMA_signal_19600 ;
    wire new_AGEMA_signal_19601 ;
    wire new_AGEMA_signal_19602 ;
    wire new_AGEMA_signal_19603 ;
    wire new_AGEMA_signal_19604 ;
    wire new_AGEMA_signal_19605 ;
    wire new_AGEMA_signal_19606 ;
    wire new_AGEMA_signal_19607 ;
    wire new_AGEMA_signal_19608 ;
    wire new_AGEMA_signal_19609 ;
    wire new_AGEMA_signal_19610 ;
    wire new_AGEMA_signal_19611 ;
    wire new_AGEMA_signal_19612 ;
    wire new_AGEMA_signal_19613 ;
    wire new_AGEMA_signal_19614 ;
    wire new_AGEMA_signal_19615 ;
    wire new_AGEMA_signal_19616 ;
    wire new_AGEMA_signal_19617 ;
    wire new_AGEMA_signal_19618 ;
    wire new_AGEMA_signal_19619 ;
    wire new_AGEMA_signal_19620 ;
    wire new_AGEMA_signal_19621 ;
    wire new_AGEMA_signal_19622 ;
    wire new_AGEMA_signal_19623 ;
    wire new_AGEMA_signal_19624 ;
    wire new_AGEMA_signal_19625 ;
    wire new_AGEMA_signal_19626 ;
    wire new_AGEMA_signal_19627 ;
    wire new_AGEMA_signal_19628 ;
    wire new_AGEMA_signal_19629 ;
    wire new_AGEMA_signal_19630 ;
    wire new_AGEMA_signal_19631 ;
    wire new_AGEMA_signal_19632 ;
    wire new_AGEMA_signal_19633 ;
    wire new_AGEMA_signal_19634 ;
    wire new_AGEMA_signal_19635 ;
    wire new_AGEMA_signal_19636 ;
    wire new_AGEMA_signal_19637 ;
    wire new_AGEMA_signal_19638 ;
    wire new_AGEMA_signal_19639 ;
    wire new_AGEMA_signal_19640 ;
    wire new_AGEMA_signal_19641 ;
    wire new_AGEMA_signal_19642 ;
    wire new_AGEMA_signal_19643 ;
    wire new_AGEMA_signal_19644 ;
    wire new_AGEMA_signal_19645 ;
    wire new_AGEMA_signal_19646 ;
    wire new_AGEMA_signal_19647 ;
    wire new_AGEMA_signal_19648 ;
    wire new_AGEMA_signal_19649 ;
    wire new_AGEMA_signal_19650 ;
    wire new_AGEMA_signal_19651 ;
    wire new_AGEMA_signal_19652 ;
    wire new_AGEMA_signal_19653 ;
    wire new_AGEMA_signal_19654 ;
    wire new_AGEMA_signal_19655 ;
    wire new_AGEMA_signal_19656 ;
    wire new_AGEMA_signal_19657 ;
    wire new_AGEMA_signal_19658 ;
    wire new_AGEMA_signal_19659 ;
    wire new_AGEMA_signal_19660 ;
    wire new_AGEMA_signal_19661 ;
    wire new_AGEMA_signal_19662 ;
    wire new_AGEMA_signal_19663 ;
    wire new_AGEMA_signal_19664 ;
    wire new_AGEMA_signal_19665 ;
    wire new_AGEMA_signal_19666 ;
    wire new_AGEMA_signal_19667 ;
    wire new_AGEMA_signal_19668 ;
    wire new_AGEMA_signal_19669 ;
    wire new_AGEMA_signal_19670 ;
    wire new_AGEMA_signal_19671 ;
    wire new_AGEMA_signal_19672 ;
    wire new_AGEMA_signal_19673 ;
    wire new_AGEMA_signal_19674 ;
    wire new_AGEMA_signal_19675 ;
    wire new_AGEMA_signal_19676 ;
    wire new_AGEMA_signal_19677 ;
    wire new_AGEMA_signal_19678 ;
    wire new_AGEMA_signal_19679 ;
    wire new_AGEMA_signal_19680 ;
    wire new_AGEMA_signal_19681 ;
    wire new_AGEMA_signal_19682 ;
    wire new_AGEMA_signal_19683 ;
    wire new_AGEMA_signal_19684 ;
    wire new_AGEMA_signal_19685 ;
    wire new_AGEMA_signal_19686 ;
    wire new_AGEMA_signal_19687 ;
    wire new_AGEMA_signal_19688 ;
    wire new_AGEMA_signal_19689 ;
    wire new_AGEMA_signal_19690 ;
    wire new_AGEMA_signal_19691 ;
    wire new_AGEMA_signal_19692 ;
    wire new_AGEMA_signal_19693 ;
    wire new_AGEMA_signal_19694 ;
    wire new_AGEMA_signal_19695 ;
    wire new_AGEMA_signal_19696 ;
    wire new_AGEMA_signal_19697 ;
    wire new_AGEMA_signal_19698 ;
    wire new_AGEMA_signal_19699 ;
    wire new_AGEMA_signal_19700 ;
    wire new_AGEMA_signal_19701 ;
    wire new_AGEMA_signal_19702 ;
    wire new_AGEMA_signal_19703 ;
    wire new_AGEMA_signal_19704 ;
    wire new_AGEMA_signal_19705 ;
    wire new_AGEMA_signal_19706 ;
    wire new_AGEMA_signal_19707 ;
    wire new_AGEMA_signal_19708 ;
    wire new_AGEMA_signal_19709 ;
    wire new_AGEMA_signal_19710 ;
    wire new_AGEMA_signal_19711 ;
    wire new_AGEMA_signal_19712 ;
    wire new_AGEMA_signal_19713 ;
    wire new_AGEMA_signal_19714 ;
    wire new_AGEMA_signal_19715 ;
    wire new_AGEMA_signal_19716 ;
    wire new_AGEMA_signal_19717 ;
    wire new_AGEMA_signal_19718 ;
    wire new_AGEMA_signal_19719 ;
    wire new_AGEMA_signal_19720 ;
    wire new_AGEMA_signal_19721 ;
    wire new_AGEMA_signal_19722 ;
    wire new_AGEMA_signal_19723 ;
    wire new_AGEMA_signal_19724 ;
    wire new_AGEMA_signal_19725 ;
    wire new_AGEMA_signal_19726 ;
    wire new_AGEMA_signal_19727 ;
    wire new_AGEMA_signal_19728 ;
    wire new_AGEMA_signal_19729 ;
    wire new_AGEMA_signal_19730 ;
    wire new_AGEMA_signal_19731 ;
    wire new_AGEMA_signal_19732 ;
    wire new_AGEMA_signal_19733 ;
    wire new_AGEMA_signal_19734 ;
    wire new_AGEMA_signal_19735 ;
    wire new_AGEMA_signal_19736 ;
    wire new_AGEMA_signal_19737 ;
    wire new_AGEMA_signal_19738 ;
    wire new_AGEMA_signal_19739 ;
    wire new_AGEMA_signal_19740 ;
    wire new_AGEMA_signal_19741 ;
    wire new_AGEMA_signal_19742 ;
    wire new_AGEMA_signal_19743 ;
    wire new_AGEMA_signal_19744 ;
    wire new_AGEMA_signal_19745 ;
    wire new_AGEMA_signal_19746 ;
    wire new_AGEMA_signal_19747 ;
    wire new_AGEMA_signal_19748 ;
    wire new_AGEMA_signal_19749 ;
    wire new_AGEMA_signal_19750 ;
    wire new_AGEMA_signal_19751 ;
    wire new_AGEMA_signal_19752 ;
    wire new_AGEMA_signal_19753 ;
    wire new_AGEMA_signal_19754 ;
    wire new_AGEMA_signal_19755 ;
    wire new_AGEMA_signal_19756 ;
    wire new_AGEMA_signal_19757 ;
    wire new_AGEMA_signal_19758 ;
    wire new_AGEMA_signal_19759 ;
    wire new_AGEMA_signal_19760 ;
    wire new_AGEMA_signal_19761 ;
    wire new_AGEMA_signal_19762 ;
    wire new_AGEMA_signal_19763 ;
    wire new_AGEMA_signal_19764 ;
    wire new_AGEMA_signal_19765 ;
    wire new_AGEMA_signal_19766 ;
    wire new_AGEMA_signal_19767 ;
    wire new_AGEMA_signal_19768 ;
    wire new_AGEMA_signal_19769 ;
    wire new_AGEMA_signal_19770 ;
    wire new_AGEMA_signal_19771 ;
    wire new_AGEMA_signal_19772 ;
    wire new_AGEMA_signal_19773 ;
    wire new_AGEMA_signal_19774 ;
    wire new_AGEMA_signal_19775 ;
    wire new_AGEMA_signal_19776 ;
    wire new_AGEMA_signal_19777 ;
    wire new_AGEMA_signal_19778 ;
    wire new_AGEMA_signal_19779 ;
    wire new_AGEMA_signal_19780 ;
    wire new_AGEMA_signal_19781 ;
    wire new_AGEMA_signal_19782 ;
    wire new_AGEMA_signal_19783 ;
    wire new_AGEMA_signal_19784 ;
    wire new_AGEMA_signal_19785 ;
    wire new_AGEMA_signal_19786 ;
    wire new_AGEMA_signal_19787 ;
    wire new_AGEMA_signal_19788 ;
    wire new_AGEMA_signal_19789 ;
    wire new_AGEMA_signal_19790 ;
    wire new_AGEMA_signal_19791 ;
    wire new_AGEMA_signal_19792 ;
    wire new_AGEMA_signal_19793 ;
    wire new_AGEMA_signal_19794 ;
    wire new_AGEMA_signal_19795 ;
    wire new_AGEMA_signal_19796 ;
    wire new_AGEMA_signal_19797 ;
    wire new_AGEMA_signal_19798 ;
    wire new_AGEMA_signal_19799 ;
    wire new_AGEMA_signal_19800 ;
    wire new_AGEMA_signal_19801 ;
    wire new_AGEMA_signal_19802 ;
    wire new_AGEMA_signal_19803 ;
    wire new_AGEMA_signal_19804 ;
    wire new_AGEMA_signal_19805 ;
    wire new_AGEMA_signal_19806 ;
    wire new_AGEMA_signal_19807 ;
    wire new_AGEMA_signal_19808 ;
    wire new_AGEMA_signal_19809 ;
    wire new_AGEMA_signal_19810 ;
    wire new_AGEMA_signal_19811 ;
    wire new_AGEMA_signal_19812 ;
    wire new_AGEMA_signal_19813 ;
    wire new_AGEMA_signal_19814 ;
    wire new_AGEMA_signal_19815 ;
    wire new_AGEMA_signal_19816 ;
    wire new_AGEMA_signal_19817 ;
    wire new_AGEMA_signal_19818 ;
    wire new_AGEMA_signal_19819 ;
    wire new_AGEMA_signal_19820 ;
    wire new_AGEMA_signal_19821 ;
    wire new_AGEMA_signal_19822 ;
    wire new_AGEMA_signal_19823 ;
    wire new_AGEMA_signal_19824 ;
    wire new_AGEMA_signal_19825 ;
    wire new_AGEMA_signal_19826 ;
    wire new_AGEMA_signal_19827 ;
    wire new_AGEMA_signal_19828 ;
    wire new_AGEMA_signal_19829 ;
    wire new_AGEMA_signal_19830 ;
    wire new_AGEMA_signal_19831 ;
    wire new_AGEMA_signal_19832 ;
    wire new_AGEMA_signal_19833 ;
    wire new_AGEMA_signal_19834 ;
    wire new_AGEMA_signal_19835 ;
    wire new_AGEMA_signal_19836 ;
    wire new_AGEMA_signal_19837 ;
    wire new_AGEMA_signal_19838 ;
    wire new_AGEMA_signal_19839 ;
    wire new_AGEMA_signal_19840 ;
    wire new_AGEMA_signal_19841 ;
    wire new_AGEMA_signal_19842 ;
    wire new_AGEMA_signal_19843 ;
    wire new_AGEMA_signal_19844 ;
    wire new_AGEMA_signal_19845 ;
    wire new_AGEMA_signal_19846 ;
    wire new_AGEMA_signal_19847 ;
    wire new_AGEMA_signal_19848 ;
    wire new_AGEMA_signal_19849 ;
    wire new_AGEMA_signal_19850 ;
    wire new_AGEMA_signal_19851 ;
    wire new_AGEMA_signal_19852 ;
    wire new_AGEMA_signal_19853 ;
    wire new_AGEMA_signal_19854 ;
    wire new_AGEMA_signal_19855 ;
    wire new_AGEMA_signal_19856 ;
    wire new_AGEMA_signal_19857 ;
    wire new_AGEMA_signal_19858 ;
    wire new_AGEMA_signal_19859 ;
    wire new_AGEMA_signal_19860 ;
    wire new_AGEMA_signal_19861 ;
    wire new_AGEMA_signal_19862 ;
    wire new_AGEMA_signal_19863 ;
    wire new_AGEMA_signal_19864 ;
    wire new_AGEMA_signal_19865 ;
    wire new_AGEMA_signal_19866 ;
    wire new_AGEMA_signal_19867 ;
    wire new_AGEMA_signal_19868 ;
    wire new_AGEMA_signal_19869 ;
    wire new_AGEMA_signal_19870 ;
    wire new_AGEMA_signal_19871 ;
    wire new_AGEMA_signal_19872 ;
    wire new_AGEMA_signal_19873 ;
    wire new_AGEMA_signal_19874 ;
    wire new_AGEMA_signal_19875 ;
    wire new_AGEMA_signal_19876 ;
    wire new_AGEMA_signal_19877 ;
    wire new_AGEMA_signal_19878 ;
    wire new_AGEMA_signal_19879 ;
    wire new_AGEMA_signal_19880 ;
    wire new_AGEMA_signal_19881 ;
    wire new_AGEMA_signal_19882 ;
    wire new_AGEMA_signal_19883 ;
    wire new_AGEMA_signal_19884 ;
    wire new_AGEMA_signal_19885 ;
    wire new_AGEMA_signal_19886 ;
    wire new_AGEMA_signal_19887 ;
    wire new_AGEMA_signal_19888 ;
    wire new_AGEMA_signal_19889 ;
    wire new_AGEMA_signal_19890 ;
    wire new_AGEMA_signal_19891 ;
    wire new_AGEMA_signal_19892 ;
    wire new_AGEMA_signal_19893 ;
    wire new_AGEMA_signal_19894 ;
    wire new_AGEMA_signal_19895 ;
    wire new_AGEMA_signal_19896 ;
    wire new_AGEMA_signal_19897 ;
    wire new_AGEMA_signal_19898 ;
    wire new_AGEMA_signal_19899 ;
    wire new_AGEMA_signal_19900 ;
    wire new_AGEMA_signal_19901 ;
    wire new_AGEMA_signal_19902 ;
    wire new_AGEMA_signal_19903 ;
    wire new_AGEMA_signal_19904 ;
    wire new_AGEMA_signal_19905 ;
    wire new_AGEMA_signal_19906 ;
    wire new_AGEMA_signal_19907 ;
    wire new_AGEMA_signal_19908 ;
    wire new_AGEMA_signal_19909 ;
    wire new_AGEMA_signal_19910 ;
    wire new_AGEMA_signal_19911 ;
    wire new_AGEMA_signal_19912 ;
    wire new_AGEMA_signal_19913 ;
    wire new_AGEMA_signal_19914 ;
    wire new_AGEMA_signal_19915 ;
    wire new_AGEMA_signal_19916 ;
    wire new_AGEMA_signal_19917 ;
    wire new_AGEMA_signal_19918 ;
    wire new_AGEMA_signal_19919 ;
    wire new_AGEMA_signal_19920 ;
    wire new_AGEMA_signal_19921 ;
    wire new_AGEMA_signal_19922 ;
    wire new_AGEMA_signal_19923 ;
    wire new_AGEMA_signal_19924 ;
    wire new_AGEMA_signal_19925 ;
    wire new_AGEMA_signal_19926 ;
    wire new_AGEMA_signal_19927 ;
    wire new_AGEMA_signal_19928 ;
    wire new_AGEMA_signal_19929 ;
    wire new_AGEMA_signal_19930 ;
    wire new_AGEMA_signal_19931 ;
    wire new_AGEMA_signal_19932 ;
    wire new_AGEMA_signal_19933 ;
    wire new_AGEMA_signal_19934 ;
    wire new_AGEMA_signal_19935 ;
    wire new_AGEMA_signal_19936 ;
    wire new_AGEMA_signal_19937 ;
    wire new_AGEMA_signal_19938 ;
    wire new_AGEMA_signal_19939 ;
    wire new_AGEMA_signal_19940 ;
    wire new_AGEMA_signal_19941 ;
    wire new_AGEMA_signal_19942 ;
    wire new_AGEMA_signal_19943 ;
    wire new_AGEMA_signal_19944 ;
    wire new_AGEMA_signal_19945 ;
    wire new_AGEMA_signal_19946 ;
    wire new_AGEMA_signal_19947 ;
    wire new_AGEMA_signal_19948 ;
    wire new_AGEMA_signal_19949 ;
    wire new_AGEMA_signal_19950 ;
    wire new_AGEMA_signal_19951 ;
    wire new_AGEMA_signal_19952 ;
    wire new_AGEMA_signal_19953 ;
    wire new_AGEMA_signal_19954 ;
    wire new_AGEMA_signal_19955 ;
    wire new_AGEMA_signal_19956 ;
    wire new_AGEMA_signal_19957 ;
    wire new_AGEMA_signal_19958 ;
    wire new_AGEMA_signal_19959 ;
    wire new_AGEMA_signal_19960 ;
    wire new_AGEMA_signal_19961 ;
    wire new_AGEMA_signal_19962 ;
    wire new_AGEMA_signal_19963 ;
    wire new_AGEMA_signal_19964 ;
    wire new_AGEMA_signal_19965 ;
    wire new_AGEMA_signal_19966 ;
    wire new_AGEMA_signal_19967 ;
    wire new_AGEMA_signal_19968 ;
    wire new_AGEMA_signal_19969 ;
    wire new_AGEMA_signal_19970 ;
    wire new_AGEMA_signal_19971 ;
    wire new_AGEMA_signal_19972 ;
    wire new_AGEMA_signal_19973 ;
    wire new_AGEMA_signal_19974 ;
    wire new_AGEMA_signal_19975 ;
    wire new_AGEMA_signal_19976 ;
    wire new_AGEMA_signal_19977 ;
    wire new_AGEMA_signal_19978 ;
    wire new_AGEMA_signal_19979 ;
    wire new_AGEMA_signal_19980 ;
    wire new_AGEMA_signal_19981 ;
    wire new_AGEMA_signal_19982 ;
    wire new_AGEMA_signal_19983 ;
    wire new_AGEMA_signal_19984 ;
    wire new_AGEMA_signal_19985 ;
    wire new_AGEMA_signal_19986 ;
    wire new_AGEMA_signal_19987 ;
    wire new_AGEMA_signal_19988 ;
    wire new_AGEMA_signal_19989 ;
    wire new_AGEMA_signal_19990 ;
    wire new_AGEMA_signal_19991 ;
    wire new_AGEMA_signal_19992 ;
    wire new_AGEMA_signal_19993 ;
    wire new_AGEMA_signal_19994 ;
    wire new_AGEMA_signal_19995 ;
    wire new_AGEMA_signal_19996 ;
    wire new_AGEMA_signal_19997 ;
    wire new_AGEMA_signal_19998 ;
    wire new_AGEMA_signal_19999 ;
    wire new_AGEMA_signal_20000 ;
    wire new_AGEMA_signal_20001 ;
    wire new_AGEMA_signal_20002 ;
    wire new_AGEMA_signal_20003 ;
    wire new_AGEMA_signal_20004 ;
    wire new_AGEMA_signal_20005 ;
    wire new_AGEMA_signal_20006 ;
    wire new_AGEMA_signal_20007 ;
    wire new_AGEMA_signal_20008 ;
    wire new_AGEMA_signal_20009 ;
    wire new_AGEMA_signal_20010 ;
    wire new_AGEMA_signal_20011 ;
    wire new_AGEMA_signal_20012 ;
    wire new_AGEMA_signal_20013 ;
    wire new_AGEMA_signal_20014 ;
    wire new_AGEMA_signal_20015 ;
    wire new_AGEMA_signal_20016 ;
    wire new_AGEMA_signal_20017 ;
    wire new_AGEMA_signal_20018 ;
    wire new_AGEMA_signal_20019 ;
    wire new_AGEMA_signal_20020 ;
    wire new_AGEMA_signal_20021 ;
    wire new_AGEMA_signal_20022 ;
    wire new_AGEMA_signal_20023 ;
    wire new_AGEMA_signal_20024 ;
    wire new_AGEMA_signal_20025 ;
    wire new_AGEMA_signal_20026 ;
    wire new_AGEMA_signal_20027 ;
    wire new_AGEMA_signal_20028 ;
    wire new_AGEMA_signal_20029 ;
    wire new_AGEMA_signal_20030 ;
    wire new_AGEMA_signal_20031 ;
    wire new_AGEMA_signal_20032 ;
    wire new_AGEMA_signal_20033 ;
    wire new_AGEMA_signal_20034 ;
    wire new_AGEMA_signal_20035 ;
    wire new_AGEMA_signal_20036 ;
    wire new_AGEMA_signal_20037 ;
    wire new_AGEMA_signal_20038 ;
    wire new_AGEMA_signal_20039 ;
    wire new_AGEMA_signal_20040 ;
    wire new_AGEMA_signal_20041 ;
    wire new_AGEMA_signal_20042 ;
    wire new_AGEMA_signal_20043 ;
    wire new_AGEMA_signal_20044 ;
    wire new_AGEMA_signal_20045 ;
    wire new_AGEMA_signal_20046 ;
    wire new_AGEMA_signal_20047 ;
    wire new_AGEMA_signal_20048 ;
    wire new_AGEMA_signal_20049 ;
    wire new_AGEMA_signal_20050 ;
    wire new_AGEMA_signal_20051 ;
    wire new_AGEMA_signal_20052 ;
    wire new_AGEMA_signal_20053 ;
    wire new_AGEMA_signal_20054 ;
    wire new_AGEMA_signal_20055 ;
    wire new_AGEMA_signal_20056 ;
    wire new_AGEMA_signal_20057 ;
    wire new_AGEMA_signal_20058 ;
    wire new_AGEMA_signal_20059 ;
    wire new_AGEMA_signal_20060 ;
    wire new_AGEMA_signal_20061 ;
    wire new_AGEMA_signal_20062 ;
    wire new_AGEMA_signal_20063 ;
    wire new_AGEMA_signal_20064 ;
    wire new_AGEMA_signal_20065 ;
    wire new_AGEMA_signal_20066 ;
    wire new_AGEMA_signal_20067 ;
    wire new_AGEMA_signal_20068 ;
    wire new_AGEMA_signal_20069 ;
    wire new_AGEMA_signal_20070 ;
    wire new_AGEMA_signal_20071 ;
    wire new_AGEMA_signal_20072 ;
    wire new_AGEMA_signal_20073 ;
    wire new_AGEMA_signal_20074 ;
    wire new_AGEMA_signal_20075 ;
    wire new_AGEMA_signal_20076 ;
    wire new_AGEMA_signal_20077 ;
    wire new_AGEMA_signal_20078 ;
    wire new_AGEMA_signal_20079 ;
    wire new_AGEMA_signal_20080 ;
    wire new_AGEMA_signal_20081 ;
    wire new_AGEMA_signal_20082 ;
    wire new_AGEMA_signal_20083 ;
    wire new_AGEMA_signal_20084 ;
    wire new_AGEMA_signal_20085 ;
    wire new_AGEMA_signal_20086 ;
    wire new_AGEMA_signal_20087 ;
    wire new_AGEMA_signal_20088 ;
    wire new_AGEMA_signal_20089 ;
    wire new_AGEMA_signal_20090 ;
    wire new_AGEMA_signal_20091 ;
    wire new_AGEMA_signal_20092 ;
    wire new_AGEMA_signal_20093 ;
    wire new_AGEMA_signal_20094 ;
    wire new_AGEMA_signal_20095 ;
    wire new_AGEMA_signal_20096 ;
    wire new_AGEMA_signal_20097 ;
    wire new_AGEMA_signal_20098 ;
    wire new_AGEMA_signal_20099 ;
    wire new_AGEMA_signal_20100 ;
    wire new_AGEMA_signal_20101 ;
    wire new_AGEMA_signal_20102 ;
    wire new_AGEMA_signal_20103 ;
    wire new_AGEMA_signal_20104 ;
    wire new_AGEMA_signal_20105 ;
    wire new_AGEMA_signal_20106 ;
    wire new_AGEMA_signal_20107 ;
    wire new_AGEMA_signal_20108 ;
    wire new_AGEMA_signal_20109 ;
    wire new_AGEMA_signal_20110 ;
    wire new_AGEMA_signal_20111 ;
    wire new_AGEMA_signal_20112 ;
    wire new_AGEMA_signal_20113 ;
    wire new_AGEMA_signal_20114 ;
    wire new_AGEMA_signal_20115 ;
    wire new_AGEMA_signal_20116 ;
    wire new_AGEMA_signal_20117 ;
    wire new_AGEMA_signal_20118 ;
    wire new_AGEMA_signal_20119 ;
    wire new_AGEMA_signal_20120 ;
    wire new_AGEMA_signal_20121 ;
    wire new_AGEMA_signal_20122 ;
    wire new_AGEMA_signal_20123 ;
    wire new_AGEMA_signal_20124 ;
    wire new_AGEMA_signal_20125 ;
    wire new_AGEMA_signal_20126 ;
    wire new_AGEMA_signal_20127 ;
    wire new_AGEMA_signal_20128 ;
    wire new_AGEMA_signal_20129 ;
    wire new_AGEMA_signal_20130 ;
    wire new_AGEMA_signal_20131 ;
    wire new_AGEMA_signal_20132 ;
    wire new_AGEMA_signal_20133 ;
    wire new_AGEMA_signal_20134 ;
    wire new_AGEMA_signal_20135 ;
    wire new_AGEMA_signal_20136 ;
    wire new_AGEMA_signal_20137 ;
    wire new_AGEMA_signal_20138 ;
    wire new_AGEMA_signal_20139 ;
    wire new_AGEMA_signal_20140 ;
    wire new_AGEMA_signal_20141 ;
    wire new_AGEMA_signal_20142 ;
    wire new_AGEMA_signal_20143 ;
    wire new_AGEMA_signal_20144 ;
    wire new_AGEMA_signal_20145 ;
    wire new_AGEMA_signal_20146 ;
    wire new_AGEMA_signal_20147 ;
    wire new_AGEMA_signal_20148 ;
    wire new_AGEMA_signal_20149 ;
    wire new_AGEMA_signal_20150 ;
    wire new_AGEMA_signal_20151 ;
    wire new_AGEMA_signal_20152 ;
    wire new_AGEMA_signal_20153 ;
    wire new_AGEMA_signal_20154 ;
    wire new_AGEMA_signal_20155 ;
    wire new_AGEMA_signal_20156 ;
    wire new_AGEMA_signal_20157 ;
    wire new_AGEMA_signal_20158 ;
    wire new_AGEMA_signal_20159 ;
    wire new_AGEMA_signal_20160 ;
    wire new_AGEMA_signal_20161 ;
    wire new_AGEMA_signal_20162 ;
    wire new_AGEMA_signal_20163 ;
    wire new_AGEMA_signal_20164 ;
    wire new_AGEMA_signal_20165 ;
    wire new_AGEMA_signal_20166 ;
    wire new_AGEMA_signal_20167 ;
    wire new_AGEMA_signal_20168 ;
    wire new_AGEMA_signal_20169 ;
    wire new_AGEMA_signal_20170 ;
    wire new_AGEMA_signal_20171 ;
    wire new_AGEMA_signal_20172 ;
    wire new_AGEMA_signal_20173 ;
    wire new_AGEMA_signal_20174 ;
    wire new_AGEMA_signal_20175 ;
    wire new_AGEMA_signal_20176 ;
    wire new_AGEMA_signal_20177 ;
    wire new_AGEMA_signal_20178 ;
    wire new_AGEMA_signal_20179 ;
    wire new_AGEMA_signal_20180 ;
    wire new_AGEMA_signal_20181 ;
    wire new_AGEMA_signal_20182 ;
    wire new_AGEMA_signal_20183 ;
    wire new_AGEMA_signal_20184 ;
    wire new_AGEMA_signal_20185 ;
    wire new_AGEMA_signal_20186 ;
    wire new_AGEMA_signal_20187 ;
    wire new_AGEMA_signal_20188 ;
    wire new_AGEMA_signal_20189 ;
    wire new_AGEMA_signal_20190 ;
    wire new_AGEMA_signal_20191 ;
    wire new_AGEMA_signal_20192 ;
    wire new_AGEMA_signal_20193 ;
    wire new_AGEMA_signal_20194 ;
    wire new_AGEMA_signal_20195 ;
    wire new_AGEMA_signal_20196 ;
    wire new_AGEMA_signal_20197 ;
    wire new_AGEMA_signal_20198 ;
    wire new_AGEMA_signal_20199 ;
    wire new_AGEMA_signal_20200 ;
    wire new_AGEMA_signal_20201 ;
    wire new_AGEMA_signal_20202 ;
    wire new_AGEMA_signal_20203 ;
    wire new_AGEMA_signal_20204 ;
    wire new_AGEMA_signal_20205 ;
    wire new_AGEMA_signal_20206 ;
    wire new_AGEMA_signal_20207 ;
    wire new_AGEMA_signal_20208 ;
    wire new_AGEMA_signal_20209 ;
    wire new_AGEMA_signal_20210 ;
    wire new_AGEMA_signal_20211 ;
    wire new_AGEMA_signal_20212 ;
    wire new_AGEMA_signal_20213 ;
    wire new_AGEMA_signal_20214 ;
    wire new_AGEMA_signal_20215 ;
    wire new_AGEMA_signal_20216 ;
    wire new_AGEMA_signal_20217 ;
    wire new_AGEMA_signal_20218 ;
    wire new_AGEMA_signal_20219 ;
    wire new_AGEMA_signal_20220 ;
    wire new_AGEMA_signal_20221 ;
    wire new_AGEMA_signal_20222 ;
    wire new_AGEMA_signal_20223 ;
    wire new_AGEMA_signal_20224 ;
    wire new_AGEMA_signal_20225 ;
    wire new_AGEMA_signal_20226 ;
    wire new_AGEMA_signal_20227 ;
    wire new_AGEMA_signal_20228 ;
    wire new_AGEMA_signal_20229 ;
    wire new_AGEMA_signal_20230 ;
    wire new_AGEMA_signal_20231 ;
    wire new_AGEMA_signal_20232 ;
    wire new_AGEMA_signal_20233 ;
    wire new_AGEMA_signal_20234 ;
    wire new_AGEMA_signal_20235 ;
    wire new_AGEMA_signal_20236 ;
    wire new_AGEMA_signal_20237 ;
    wire new_AGEMA_signal_20238 ;
    wire new_AGEMA_signal_20239 ;
    wire new_AGEMA_signal_20240 ;
    wire new_AGEMA_signal_20241 ;
    wire new_AGEMA_signal_20242 ;
    wire new_AGEMA_signal_20243 ;
    wire new_AGEMA_signal_20244 ;
    wire new_AGEMA_signal_20245 ;
    wire new_AGEMA_signal_20246 ;
    wire new_AGEMA_signal_20247 ;
    wire new_AGEMA_signal_20248 ;
    wire new_AGEMA_signal_20249 ;
    wire new_AGEMA_signal_20250 ;
    wire new_AGEMA_signal_20251 ;
    wire new_AGEMA_signal_20252 ;
    wire new_AGEMA_signal_20253 ;
    wire new_AGEMA_signal_20254 ;
    wire new_AGEMA_signal_20255 ;
    wire new_AGEMA_signal_20256 ;
    wire new_AGEMA_signal_20257 ;
    wire new_AGEMA_signal_20258 ;
    wire new_AGEMA_signal_20259 ;
    wire new_AGEMA_signal_20260 ;
    wire new_AGEMA_signal_20261 ;
    wire new_AGEMA_signal_20262 ;
    wire new_AGEMA_signal_20263 ;
    wire new_AGEMA_signal_20264 ;
    wire new_AGEMA_signal_20265 ;
    wire new_AGEMA_signal_20266 ;
    wire new_AGEMA_signal_20267 ;
    wire new_AGEMA_signal_20268 ;
    wire new_AGEMA_signal_20269 ;
    wire new_AGEMA_signal_20270 ;
    wire new_AGEMA_signal_20271 ;
    wire new_AGEMA_signal_20272 ;
    wire new_AGEMA_signal_20273 ;
    wire new_AGEMA_signal_20274 ;
    wire new_AGEMA_signal_20275 ;
    wire new_AGEMA_signal_20276 ;
    wire new_AGEMA_signal_20277 ;
    wire new_AGEMA_signal_20278 ;
    wire new_AGEMA_signal_20279 ;
    wire new_AGEMA_signal_20280 ;
    wire new_AGEMA_signal_20281 ;
    wire new_AGEMA_signal_20282 ;
    wire new_AGEMA_signal_20283 ;
    wire new_AGEMA_signal_20284 ;
    wire new_AGEMA_signal_20285 ;
    wire new_AGEMA_signal_20286 ;
    wire new_AGEMA_signal_20287 ;
    wire new_AGEMA_signal_20288 ;
    wire new_AGEMA_signal_20289 ;
    wire new_AGEMA_signal_20290 ;
    wire new_AGEMA_signal_20291 ;
    wire new_AGEMA_signal_20292 ;
    wire new_AGEMA_signal_20293 ;
    wire new_AGEMA_signal_20294 ;
    wire new_AGEMA_signal_20295 ;
    wire new_AGEMA_signal_20296 ;
    wire new_AGEMA_signal_20297 ;
    wire new_AGEMA_signal_20298 ;
    wire new_AGEMA_signal_20299 ;
    wire new_AGEMA_signal_20300 ;
    wire new_AGEMA_signal_20301 ;
    wire new_AGEMA_signal_20302 ;
    wire new_AGEMA_signal_20303 ;
    wire new_AGEMA_signal_20304 ;
    wire new_AGEMA_signal_20305 ;
    wire new_AGEMA_signal_20306 ;
    wire new_AGEMA_signal_20307 ;
    wire new_AGEMA_signal_20308 ;
    wire new_AGEMA_signal_20309 ;
    wire new_AGEMA_signal_20310 ;
    wire new_AGEMA_signal_20311 ;
    wire new_AGEMA_signal_20312 ;
    wire new_AGEMA_signal_20313 ;
    wire new_AGEMA_signal_20314 ;
    wire new_AGEMA_signal_20315 ;
    wire new_AGEMA_signal_20316 ;
    wire new_AGEMA_signal_20317 ;
    wire new_AGEMA_signal_20318 ;
    wire new_AGEMA_signal_20319 ;
    wire new_AGEMA_signal_20320 ;
    wire new_AGEMA_signal_20321 ;
    wire new_AGEMA_signal_20322 ;
    wire new_AGEMA_signal_20323 ;
    wire new_AGEMA_signal_20324 ;
    wire new_AGEMA_signal_20325 ;
    wire new_AGEMA_signal_20326 ;
    wire new_AGEMA_signal_20327 ;
    wire new_AGEMA_signal_20328 ;
    wire new_AGEMA_signal_20329 ;
    wire new_AGEMA_signal_20330 ;
    wire new_AGEMA_signal_20331 ;
    wire new_AGEMA_signal_20332 ;
    wire new_AGEMA_signal_20333 ;
    wire new_AGEMA_signal_20334 ;
    wire new_AGEMA_signal_20335 ;
    wire new_AGEMA_signal_20336 ;
    wire new_AGEMA_signal_20337 ;
    wire new_AGEMA_signal_20338 ;
    wire new_AGEMA_signal_20339 ;
    wire new_AGEMA_signal_20340 ;
    wire new_AGEMA_signal_20341 ;
    wire new_AGEMA_signal_20342 ;
    wire new_AGEMA_signal_20343 ;
    wire new_AGEMA_signal_20344 ;
    wire new_AGEMA_signal_20345 ;
    wire new_AGEMA_signal_20346 ;
    wire new_AGEMA_signal_20347 ;
    wire new_AGEMA_signal_20348 ;
    wire new_AGEMA_signal_20349 ;
    wire new_AGEMA_signal_20350 ;
    wire new_AGEMA_signal_20351 ;
    wire new_AGEMA_signal_20352 ;
    wire new_AGEMA_signal_20353 ;
    wire new_AGEMA_signal_20354 ;
    wire new_AGEMA_signal_20355 ;
    wire new_AGEMA_signal_20356 ;
    wire new_AGEMA_signal_20357 ;
    wire new_AGEMA_signal_20358 ;
    wire new_AGEMA_signal_20359 ;
    wire new_AGEMA_signal_20360 ;
    wire new_AGEMA_signal_20361 ;
    wire new_AGEMA_signal_20362 ;
    wire new_AGEMA_signal_20363 ;
    wire new_AGEMA_signal_20364 ;
    wire new_AGEMA_signal_20365 ;
    wire new_AGEMA_signal_20366 ;
    wire new_AGEMA_signal_20367 ;
    wire new_AGEMA_signal_20368 ;
    wire new_AGEMA_signal_20369 ;
    wire new_AGEMA_signal_20370 ;
    wire new_AGEMA_signal_20371 ;
    wire new_AGEMA_signal_20372 ;
    wire new_AGEMA_signal_20373 ;
    wire new_AGEMA_signal_20374 ;
    wire new_AGEMA_signal_20375 ;
    wire new_AGEMA_signal_20376 ;
    wire new_AGEMA_signal_20377 ;
    wire new_AGEMA_signal_20378 ;
    wire new_AGEMA_signal_20379 ;
    wire new_AGEMA_signal_20380 ;
    wire new_AGEMA_signal_20381 ;
    wire new_AGEMA_signal_20382 ;
    wire new_AGEMA_signal_20383 ;
    wire new_AGEMA_signal_20384 ;
    wire new_AGEMA_signal_20385 ;
    wire new_AGEMA_signal_20386 ;
    wire new_AGEMA_signal_20387 ;
    wire new_AGEMA_signal_20388 ;
    wire new_AGEMA_signal_20389 ;
    wire new_AGEMA_signal_20390 ;
    wire new_AGEMA_signal_20391 ;
    wire new_AGEMA_signal_20392 ;
    wire new_AGEMA_signal_20393 ;
    wire new_AGEMA_signal_20394 ;
    wire new_AGEMA_signal_20395 ;
    wire new_AGEMA_signal_20396 ;
    wire new_AGEMA_signal_20397 ;
    wire new_AGEMA_signal_20398 ;
    wire new_AGEMA_signal_20399 ;
    wire new_AGEMA_signal_20400 ;
    wire new_AGEMA_signal_20401 ;
    wire new_AGEMA_signal_20402 ;
    wire new_AGEMA_signal_20403 ;
    wire new_AGEMA_signal_20404 ;
    wire new_AGEMA_signal_20405 ;
    wire new_AGEMA_signal_20406 ;
    wire new_AGEMA_signal_20407 ;
    wire new_AGEMA_signal_20408 ;
    wire new_AGEMA_signal_20409 ;
    wire new_AGEMA_signal_20410 ;
    wire new_AGEMA_signal_20411 ;
    wire new_AGEMA_signal_20412 ;
    wire new_AGEMA_signal_20413 ;
    wire new_AGEMA_signal_20414 ;
    wire new_AGEMA_signal_20415 ;
    wire new_AGEMA_signal_20416 ;
    wire new_AGEMA_signal_20417 ;
    wire new_AGEMA_signal_20418 ;
    wire new_AGEMA_signal_20419 ;
    wire new_AGEMA_signal_20420 ;
    wire new_AGEMA_signal_20421 ;
    wire new_AGEMA_signal_20422 ;
    wire new_AGEMA_signal_20423 ;
    wire new_AGEMA_signal_20424 ;
    wire new_AGEMA_signal_20425 ;
    wire new_AGEMA_signal_20426 ;
    wire new_AGEMA_signal_20427 ;
    wire new_AGEMA_signal_20428 ;
    wire new_AGEMA_signal_20429 ;
    wire new_AGEMA_signal_20430 ;
    wire new_AGEMA_signal_20431 ;
    wire new_AGEMA_signal_20432 ;
    wire new_AGEMA_signal_20433 ;
    wire new_AGEMA_signal_20434 ;
    wire new_AGEMA_signal_20435 ;
    wire new_AGEMA_signal_20436 ;
    wire new_AGEMA_signal_20437 ;
    wire new_AGEMA_signal_20438 ;
    wire new_AGEMA_signal_20439 ;
    wire new_AGEMA_signal_20440 ;
    wire new_AGEMA_signal_20441 ;
    wire new_AGEMA_signal_20442 ;
    wire new_AGEMA_signal_20443 ;
    wire new_AGEMA_signal_20444 ;
    wire new_AGEMA_signal_20445 ;
    wire new_AGEMA_signal_20446 ;
    wire new_AGEMA_signal_20447 ;
    wire new_AGEMA_signal_20448 ;
    wire new_AGEMA_signal_20449 ;
    wire new_AGEMA_signal_20450 ;
    wire new_AGEMA_signal_20451 ;
    wire new_AGEMA_signal_20452 ;
    wire new_AGEMA_signal_20453 ;
    wire new_AGEMA_signal_20454 ;
    wire new_AGEMA_signal_20455 ;
    wire new_AGEMA_signal_20456 ;
    wire new_AGEMA_signal_20457 ;
    wire new_AGEMA_signal_20458 ;
    wire new_AGEMA_signal_20459 ;
    wire new_AGEMA_signal_20460 ;
    wire new_AGEMA_signal_20461 ;
    wire new_AGEMA_signal_20462 ;
    wire new_AGEMA_signal_20463 ;
    wire new_AGEMA_signal_20464 ;
    wire new_AGEMA_signal_20465 ;
    wire new_AGEMA_signal_20466 ;
    wire new_AGEMA_signal_20467 ;
    wire new_AGEMA_signal_20468 ;
    wire new_AGEMA_signal_20469 ;
    wire new_AGEMA_signal_20470 ;
    wire new_AGEMA_signal_20471 ;
    wire new_AGEMA_signal_20472 ;
    wire new_AGEMA_signal_20473 ;
    wire new_AGEMA_signal_20474 ;
    wire new_AGEMA_signal_20475 ;
    wire new_AGEMA_signal_20476 ;
    wire new_AGEMA_signal_20477 ;
    wire new_AGEMA_signal_20478 ;
    wire new_AGEMA_signal_20479 ;
    wire new_AGEMA_signal_20480 ;
    wire new_AGEMA_signal_20481 ;
    wire new_AGEMA_signal_20482 ;
    wire new_AGEMA_signal_20483 ;
    wire new_AGEMA_signal_20484 ;
    wire new_AGEMA_signal_20485 ;
    wire new_AGEMA_signal_20486 ;
    wire new_AGEMA_signal_20487 ;
    wire new_AGEMA_signal_20488 ;
    wire new_AGEMA_signal_20489 ;
    wire new_AGEMA_signal_20490 ;
    wire new_AGEMA_signal_20491 ;
    wire new_AGEMA_signal_20492 ;
    wire new_AGEMA_signal_20493 ;
    wire new_AGEMA_signal_20494 ;
    wire new_AGEMA_signal_20495 ;
    wire new_AGEMA_signal_20496 ;
    wire new_AGEMA_signal_20497 ;
    wire new_AGEMA_signal_20498 ;
    wire new_AGEMA_signal_20499 ;
    wire new_AGEMA_signal_20500 ;
    wire new_AGEMA_signal_20501 ;
    wire new_AGEMA_signal_20502 ;
    wire new_AGEMA_signal_20503 ;
    wire new_AGEMA_signal_20504 ;
    wire new_AGEMA_signal_20505 ;
    wire new_AGEMA_signal_20506 ;
    wire new_AGEMA_signal_20507 ;
    wire new_AGEMA_signal_20508 ;
    wire new_AGEMA_signal_20509 ;
    wire new_AGEMA_signal_20510 ;
    wire new_AGEMA_signal_20511 ;
    wire new_AGEMA_signal_20512 ;
    wire new_AGEMA_signal_20513 ;
    wire new_AGEMA_signal_20514 ;
    wire new_AGEMA_signal_20515 ;
    wire new_AGEMA_signal_20516 ;
    wire new_AGEMA_signal_20517 ;
    wire new_AGEMA_signal_20518 ;
    wire new_AGEMA_signal_20519 ;
    wire new_AGEMA_signal_20520 ;
    wire new_AGEMA_signal_20521 ;
    wire new_AGEMA_signal_20522 ;
    wire new_AGEMA_signal_20523 ;
    wire new_AGEMA_signal_20524 ;
    wire new_AGEMA_signal_20525 ;
    wire new_AGEMA_signal_20526 ;
    wire new_AGEMA_signal_20527 ;
    wire new_AGEMA_signal_20528 ;
    wire new_AGEMA_signal_20529 ;
    wire new_AGEMA_signal_20530 ;
    wire new_AGEMA_signal_20531 ;
    wire new_AGEMA_signal_20532 ;
    wire new_AGEMA_signal_20533 ;
    wire new_AGEMA_signal_20534 ;
    wire new_AGEMA_signal_20535 ;
    wire new_AGEMA_signal_20536 ;
    wire new_AGEMA_signal_20537 ;
    wire new_AGEMA_signal_20538 ;
    wire new_AGEMA_signal_20539 ;
    wire new_AGEMA_signal_20540 ;
    wire new_AGEMA_signal_20541 ;
    wire new_AGEMA_signal_20542 ;
    wire new_AGEMA_signal_20543 ;
    wire new_AGEMA_signal_20544 ;
    wire new_AGEMA_signal_20545 ;
    wire new_AGEMA_signal_20546 ;
    wire new_AGEMA_signal_20547 ;
    wire new_AGEMA_signal_20548 ;
    wire new_AGEMA_signal_20549 ;
    wire new_AGEMA_signal_20550 ;
    wire new_AGEMA_signal_20551 ;
    wire new_AGEMA_signal_20552 ;
    wire new_AGEMA_signal_20553 ;
    wire new_AGEMA_signal_20554 ;
    wire new_AGEMA_signal_20555 ;
    wire new_AGEMA_signal_20556 ;
    wire new_AGEMA_signal_20557 ;
    wire new_AGEMA_signal_20558 ;
    wire new_AGEMA_signal_20559 ;
    wire new_AGEMA_signal_20560 ;
    wire new_AGEMA_signal_20561 ;
    wire new_AGEMA_signal_20562 ;
    wire new_AGEMA_signal_20563 ;
    wire new_AGEMA_signal_20564 ;
    wire new_AGEMA_signal_20565 ;
    wire new_AGEMA_signal_20566 ;
    wire new_AGEMA_signal_20567 ;
    wire new_AGEMA_signal_20568 ;
    wire new_AGEMA_signal_20569 ;
    wire new_AGEMA_signal_20570 ;
    wire new_AGEMA_signal_20571 ;
    wire new_AGEMA_signal_20572 ;
    wire new_AGEMA_signal_20573 ;
    wire new_AGEMA_signal_20574 ;
    wire new_AGEMA_signal_20575 ;
    wire new_AGEMA_signal_20576 ;
    wire new_AGEMA_signal_20577 ;
    wire new_AGEMA_signal_20578 ;
    wire new_AGEMA_signal_20579 ;
    wire new_AGEMA_signal_20580 ;
    wire new_AGEMA_signal_20581 ;
    wire new_AGEMA_signal_20582 ;
    wire new_AGEMA_signal_20583 ;
    wire new_AGEMA_signal_20584 ;
    wire new_AGEMA_signal_20585 ;
    wire new_AGEMA_signal_20586 ;
    wire new_AGEMA_signal_20587 ;
    wire new_AGEMA_signal_20588 ;
    wire new_AGEMA_signal_20589 ;
    wire new_AGEMA_signal_20590 ;
    wire new_AGEMA_signal_20591 ;
    wire new_AGEMA_signal_20592 ;
    wire new_AGEMA_signal_20593 ;
    wire new_AGEMA_signal_20594 ;
    wire new_AGEMA_signal_20595 ;
    wire new_AGEMA_signal_20596 ;
    wire new_AGEMA_signal_20597 ;
    wire new_AGEMA_signal_20598 ;
    wire new_AGEMA_signal_20599 ;
    wire new_AGEMA_signal_20600 ;
    wire new_AGEMA_signal_20601 ;
    wire new_AGEMA_signal_20602 ;
    wire new_AGEMA_signal_20603 ;
    wire new_AGEMA_signal_20604 ;
    wire new_AGEMA_signal_20605 ;
    wire new_AGEMA_signal_20606 ;
    wire new_AGEMA_signal_20607 ;
    wire new_AGEMA_signal_20608 ;
    wire new_AGEMA_signal_20609 ;
    wire new_AGEMA_signal_20610 ;
    wire new_AGEMA_signal_20611 ;
    wire new_AGEMA_signal_20612 ;
    wire new_AGEMA_signal_20613 ;
    wire new_AGEMA_signal_20614 ;
    wire new_AGEMA_signal_20615 ;
    wire new_AGEMA_signal_20616 ;
    wire new_AGEMA_signal_20617 ;
    wire new_AGEMA_signal_20618 ;
    wire new_AGEMA_signal_20619 ;
    wire new_AGEMA_signal_20620 ;
    wire new_AGEMA_signal_20621 ;
    wire new_AGEMA_signal_20622 ;
    wire new_AGEMA_signal_20623 ;
    wire new_AGEMA_signal_20624 ;
    wire new_AGEMA_signal_20625 ;
    wire new_AGEMA_signal_20626 ;
    wire new_AGEMA_signal_20627 ;
    wire new_AGEMA_signal_20628 ;
    wire new_AGEMA_signal_20629 ;
    wire new_AGEMA_signal_20630 ;
    wire new_AGEMA_signal_20631 ;
    wire new_AGEMA_signal_20632 ;
    wire new_AGEMA_signal_20633 ;
    wire new_AGEMA_signal_20634 ;
    wire new_AGEMA_signal_20635 ;
    wire new_AGEMA_signal_20636 ;
    wire new_AGEMA_signal_20637 ;
    wire new_AGEMA_signal_20638 ;
    wire new_AGEMA_signal_20639 ;
    wire new_AGEMA_signal_20640 ;
    wire new_AGEMA_signal_20641 ;
    wire new_AGEMA_signal_20642 ;
    wire new_AGEMA_signal_20643 ;
    wire new_AGEMA_signal_20644 ;
    wire new_AGEMA_signal_20645 ;
    wire new_AGEMA_signal_20646 ;
    wire new_AGEMA_signal_20647 ;
    wire new_AGEMA_signal_20648 ;
    wire new_AGEMA_signal_20649 ;
    wire new_AGEMA_signal_20650 ;
    wire new_AGEMA_signal_20651 ;
    wire new_AGEMA_signal_20652 ;
    wire new_AGEMA_signal_20653 ;
    wire new_AGEMA_signal_20654 ;
    wire new_AGEMA_signal_20655 ;
    wire new_AGEMA_signal_20656 ;
    wire new_AGEMA_signal_20657 ;
    wire new_AGEMA_signal_20658 ;
    wire new_AGEMA_signal_20659 ;
    wire new_AGEMA_signal_20660 ;
    wire new_AGEMA_signal_20661 ;
    wire new_AGEMA_signal_20662 ;
    wire new_AGEMA_signal_20663 ;
    wire new_AGEMA_signal_20664 ;
    wire new_AGEMA_signal_20665 ;
    wire new_AGEMA_signal_20666 ;
    wire new_AGEMA_signal_20667 ;
    wire new_AGEMA_signal_20668 ;
    wire new_AGEMA_signal_20669 ;
    wire new_AGEMA_signal_20670 ;
    wire new_AGEMA_signal_20671 ;
    wire new_AGEMA_signal_20672 ;
    wire new_AGEMA_signal_20673 ;
    wire new_AGEMA_signal_20674 ;
    wire new_AGEMA_signal_20675 ;
    wire new_AGEMA_signal_20676 ;
    wire new_AGEMA_signal_20677 ;
    wire new_AGEMA_signal_20678 ;
    wire new_AGEMA_signal_20679 ;
    wire new_AGEMA_signal_20680 ;
    wire new_AGEMA_signal_20681 ;
    wire new_AGEMA_signal_20682 ;
    wire new_AGEMA_signal_20683 ;
    wire new_AGEMA_signal_20684 ;
    wire new_AGEMA_signal_20685 ;
    wire new_AGEMA_signal_20686 ;
    wire new_AGEMA_signal_20687 ;
    wire new_AGEMA_signal_20688 ;
    wire new_AGEMA_signal_20689 ;
    wire new_AGEMA_signal_20690 ;
    wire new_AGEMA_signal_20691 ;
    wire new_AGEMA_signal_20692 ;
    wire new_AGEMA_signal_20693 ;
    wire new_AGEMA_signal_20694 ;
    wire new_AGEMA_signal_20695 ;
    wire new_AGEMA_signal_20696 ;
    wire new_AGEMA_signal_20697 ;
    wire new_AGEMA_signal_20698 ;
    wire new_AGEMA_signal_20699 ;
    wire new_AGEMA_signal_20700 ;
    wire new_AGEMA_signal_20701 ;
    wire new_AGEMA_signal_20702 ;
    wire new_AGEMA_signal_20703 ;
    wire new_AGEMA_signal_20704 ;
    wire new_AGEMA_signal_20705 ;
    wire new_AGEMA_signal_20706 ;
    wire new_AGEMA_signal_20707 ;
    wire new_AGEMA_signal_20708 ;
    wire new_AGEMA_signal_20709 ;
    wire new_AGEMA_signal_20710 ;
    wire new_AGEMA_signal_20711 ;
    wire new_AGEMA_signal_20712 ;
    wire new_AGEMA_signal_20713 ;
    wire new_AGEMA_signal_20714 ;
    wire new_AGEMA_signal_20715 ;
    wire new_AGEMA_signal_20716 ;
    wire new_AGEMA_signal_20717 ;
    wire new_AGEMA_signal_20718 ;
    wire new_AGEMA_signal_20719 ;
    wire new_AGEMA_signal_20720 ;
    wire new_AGEMA_signal_20721 ;
    wire new_AGEMA_signal_20722 ;
    wire new_AGEMA_signal_20723 ;
    wire new_AGEMA_signal_20724 ;
    wire new_AGEMA_signal_20725 ;
    wire new_AGEMA_signal_20726 ;
    wire new_AGEMA_signal_20727 ;
    wire new_AGEMA_signal_20728 ;
    wire new_AGEMA_signal_20729 ;
    wire new_AGEMA_signal_20730 ;
    wire new_AGEMA_signal_20731 ;
    wire new_AGEMA_signal_20732 ;
    wire new_AGEMA_signal_20733 ;
    wire new_AGEMA_signal_20734 ;
    wire new_AGEMA_signal_20735 ;
    wire new_AGEMA_signal_20736 ;
    wire new_AGEMA_signal_20737 ;
    wire new_AGEMA_signal_20738 ;
    wire new_AGEMA_signal_20739 ;
    wire new_AGEMA_signal_20740 ;
    wire new_AGEMA_signal_20741 ;
    wire new_AGEMA_signal_20742 ;
    wire new_AGEMA_signal_20743 ;
    wire new_AGEMA_signal_20744 ;
    wire new_AGEMA_signal_20745 ;
    wire new_AGEMA_signal_20746 ;
    wire new_AGEMA_signal_20747 ;
    wire new_AGEMA_signal_20748 ;
    wire new_AGEMA_signal_20749 ;
    wire new_AGEMA_signal_20750 ;
    wire new_AGEMA_signal_20751 ;
    wire new_AGEMA_signal_20752 ;
    wire new_AGEMA_signal_20753 ;
    wire new_AGEMA_signal_20754 ;
    wire new_AGEMA_signal_20755 ;
    wire new_AGEMA_signal_20756 ;
    wire new_AGEMA_signal_20757 ;
    wire new_AGEMA_signal_20758 ;
    wire new_AGEMA_signal_20759 ;
    wire new_AGEMA_signal_20760 ;
    wire new_AGEMA_signal_20761 ;
    wire new_AGEMA_signal_20762 ;
    wire new_AGEMA_signal_20763 ;
    wire new_AGEMA_signal_20764 ;
    wire new_AGEMA_signal_20765 ;
    wire new_AGEMA_signal_20766 ;
    wire new_AGEMA_signal_20767 ;
    wire new_AGEMA_signal_20768 ;
    wire new_AGEMA_signal_20769 ;
    wire new_AGEMA_signal_20770 ;
    wire new_AGEMA_signal_20771 ;
    wire new_AGEMA_signal_20772 ;
    wire new_AGEMA_signal_20773 ;
    wire new_AGEMA_signal_20774 ;
    wire new_AGEMA_signal_20775 ;
    wire new_AGEMA_signal_20776 ;
    wire new_AGEMA_signal_20777 ;
    wire new_AGEMA_signal_20778 ;
    wire new_AGEMA_signal_20779 ;
    wire new_AGEMA_signal_20780 ;
    wire new_AGEMA_signal_20781 ;
    wire new_AGEMA_signal_20782 ;
    wire new_AGEMA_signal_20783 ;
    wire new_AGEMA_signal_20784 ;
    wire new_AGEMA_signal_20785 ;
    wire new_AGEMA_signal_20786 ;
    wire new_AGEMA_signal_20787 ;
    wire new_AGEMA_signal_20788 ;
    wire new_AGEMA_signal_20789 ;
    wire new_AGEMA_signal_20790 ;
    wire new_AGEMA_signal_20791 ;
    wire new_AGEMA_signal_20792 ;
    wire new_AGEMA_signal_20793 ;
    wire new_AGEMA_signal_20794 ;
    wire new_AGEMA_signal_20795 ;
    wire new_AGEMA_signal_20796 ;
    wire new_AGEMA_signal_20797 ;
    wire new_AGEMA_signal_20798 ;
    wire new_AGEMA_signal_20799 ;
    wire new_AGEMA_signal_20800 ;
    wire new_AGEMA_signal_20801 ;
    wire new_AGEMA_signal_20802 ;
    wire new_AGEMA_signal_20803 ;
    wire new_AGEMA_signal_20804 ;
    wire new_AGEMA_signal_20805 ;
    wire new_AGEMA_signal_20806 ;
    wire new_AGEMA_signal_20807 ;
    wire new_AGEMA_signal_20808 ;
    wire new_AGEMA_signal_20809 ;
    wire new_AGEMA_signal_20810 ;
    wire new_AGEMA_signal_20811 ;
    wire new_AGEMA_signal_20812 ;
    wire new_AGEMA_signal_20813 ;
    wire new_AGEMA_signal_20814 ;
    wire new_AGEMA_signal_20815 ;
    wire new_AGEMA_signal_20816 ;
    wire new_AGEMA_signal_20817 ;
    wire new_AGEMA_signal_20818 ;
    wire new_AGEMA_signal_20819 ;
    wire new_AGEMA_signal_20820 ;
    wire new_AGEMA_signal_20821 ;
    wire new_AGEMA_signal_20822 ;
    wire new_AGEMA_signal_20823 ;
    wire new_AGEMA_signal_20824 ;
    wire new_AGEMA_signal_20825 ;
    wire new_AGEMA_signal_20826 ;
    wire new_AGEMA_signal_20827 ;
    wire new_AGEMA_signal_20828 ;
    wire new_AGEMA_signal_20829 ;
    wire new_AGEMA_signal_20830 ;
    wire new_AGEMA_signal_20831 ;
    wire new_AGEMA_signal_20832 ;
    wire new_AGEMA_signal_20833 ;
    wire new_AGEMA_signal_20834 ;
    wire new_AGEMA_signal_20835 ;
    wire new_AGEMA_signal_20836 ;
    wire new_AGEMA_signal_20837 ;
    wire new_AGEMA_signal_20838 ;
    wire new_AGEMA_signal_20839 ;
    wire new_AGEMA_signal_20840 ;
    wire new_AGEMA_signal_20841 ;
    wire new_AGEMA_signal_20842 ;
    wire new_AGEMA_signal_20843 ;
    wire new_AGEMA_signal_20844 ;
    wire new_AGEMA_signal_20845 ;
    wire new_AGEMA_signal_20846 ;
    wire new_AGEMA_signal_20847 ;
    wire new_AGEMA_signal_20848 ;
    wire new_AGEMA_signal_20849 ;
    wire new_AGEMA_signal_20850 ;
    wire new_AGEMA_signal_20851 ;
    wire new_AGEMA_signal_20852 ;
    wire new_AGEMA_signal_20853 ;
    wire new_AGEMA_signal_20854 ;
    wire new_AGEMA_signal_20855 ;
    wire new_AGEMA_signal_20856 ;
    wire new_AGEMA_signal_20857 ;
    wire new_AGEMA_signal_20858 ;
    wire new_AGEMA_signal_20859 ;
    wire new_AGEMA_signal_20860 ;
    wire new_AGEMA_signal_20861 ;
    wire new_AGEMA_signal_20862 ;
    wire new_AGEMA_signal_20863 ;
    wire new_AGEMA_signal_20864 ;
    wire new_AGEMA_signal_20865 ;
    wire new_AGEMA_signal_20866 ;
    wire new_AGEMA_signal_20867 ;
    wire new_AGEMA_signal_20868 ;
    wire new_AGEMA_signal_20869 ;
    wire new_AGEMA_signal_20870 ;
    wire new_AGEMA_signal_20871 ;
    wire new_AGEMA_signal_20872 ;
    wire new_AGEMA_signal_20873 ;
    wire new_AGEMA_signal_20874 ;
    wire new_AGEMA_signal_20875 ;
    wire new_AGEMA_signal_20876 ;
    wire new_AGEMA_signal_20877 ;
    wire new_AGEMA_signal_20878 ;
    wire new_AGEMA_signal_20879 ;
    wire new_AGEMA_signal_20880 ;
    wire new_AGEMA_signal_20881 ;
    wire new_AGEMA_signal_20882 ;
    wire new_AGEMA_signal_20883 ;
    wire new_AGEMA_signal_20884 ;
    wire new_AGEMA_signal_20885 ;
    wire new_AGEMA_signal_20886 ;
    wire new_AGEMA_signal_20887 ;
    wire new_AGEMA_signal_20888 ;
    wire new_AGEMA_signal_20889 ;
    wire new_AGEMA_signal_20890 ;
    wire new_AGEMA_signal_20891 ;
    wire new_AGEMA_signal_20892 ;
    wire new_AGEMA_signal_20893 ;
    wire new_AGEMA_signal_20894 ;
    wire new_AGEMA_signal_20895 ;
    wire new_AGEMA_signal_20896 ;
    wire new_AGEMA_signal_20897 ;
    wire new_AGEMA_signal_20898 ;
    wire new_AGEMA_signal_20899 ;
    wire new_AGEMA_signal_20900 ;
    wire new_AGEMA_signal_20901 ;
    wire new_AGEMA_signal_20902 ;
    wire new_AGEMA_signal_20903 ;
    wire new_AGEMA_signal_20904 ;
    wire new_AGEMA_signal_20905 ;
    wire new_AGEMA_signal_20906 ;
    wire new_AGEMA_signal_20907 ;
    wire new_AGEMA_signal_20908 ;
    wire new_AGEMA_signal_20909 ;
    wire new_AGEMA_signal_20910 ;
    wire new_AGEMA_signal_20911 ;
    wire new_AGEMA_signal_20912 ;
    wire new_AGEMA_signal_20913 ;
    wire new_AGEMA_signal_20914 ;
    wire new_AGEMA_signal_20915 ;
    wire new_AGEMA_signal_20916 ;
    wire new_AGEMA_signal_20917 ;
    wire new_AGEMA_signal_20918 ;
    wire new_AGEMA_signal_20919 ;
    wire new_AGEMA_signal_20920 ;
    wire new_AGEMA_signal_20921 ;
    wire new_AGEMA_signal_20922 ;
    wire new_AGEMA_signal_20923 ;
    wire new_AGEMA_signal_20924 ;
    wire new_AGEMA_signal_20925 ;
    wire new_AGEMA_signal_20926 ;
    wire new_AGEMA_signal_20927 ;
    wire new_AGEMA_signal_20928 ;
    wire new_AGEMA_signal_20929 ;
    wire new_AGEMA_signal_20930 ;
    wire new_AGEMA_signal_20931 ;
    wire new_AGEMA_signal_20932 ;
    wire new_AGEMA_signal_20933 ;
    wire new_AGEMA_signal_20934 ;
    wire new_AGEMA_signal_20935 ;
    wire new_AGEMA_signal_20936 ;
    wire new_AGEMA_signal_20937 ;
    wire new_AGEMA_signal_20938 ;
    wire new_AGEMA_signal_20939 ;
    wire new_AGEMA_signal_20940 ;
    wire new_AGEMA_signal_20941 ;
    wire new_AGEMA_signal_20942 ;
    wire new_AGEMA_signal_20943 ;
    wire new_AGEMA_signal_20944 ;
    wire new_AGEMA_signal_20945 ;
    wire new_AGEMA_signal_20946 ;
    wire new_AGEMA_signal_20947 ;
    wire new_AGEMA_signal_20948 ;
    wire new_AGEMA_signal_20949 ;
    wire new_AGEMA_signal_20950 ;
    wire new_AGEMA_signal_20951 ;
    wire new_AGEMA_signal_20952 ;
    wire new_AGEMA_signal_20953 ;
    wire new_AGEMA_signal_20954 ;
    wire new_AGEMA_signal_20955 ;
    wire new_AGEMA_signal_20956 ;
    wire new_AGEMA_signal_20957 ;
    wire new_AGEMA_signal_20958 ;
    wire new_AGEMA_signal_20959 ;
    wire new_AGEMA_signal_20960 ;
    wire new_AGEMA_signal_20961 ;
    wire new_AGEMA_signal_20962 ;
    wire new_AGEMA_signal_20963 ;
    wire new_AGEMA_signal_20964 ;
    wire new_AGEMA_signal_20965 ;
    wire new_AGEMA_signal_20966 ;
    wire new_AGEMA_signal_20967 ;
    wire new_AGEMA_signal_20968 ;
    wire new_AGEMA_signal_20969 ;
    wire new_AGEMA_signal_20970 ;
    wire new_AGEMA_signal_20971 ;
    wire new_AGEMA_signal_20972 ;
    wire new_AGEMA_signal_20973 ;
    wire new_AGEMA_signal_20974 ;
    wire new_AGEMA_signal_20975 ;
    wire new_AGEMA_signal_20976 ;
    wire new_AGEMA_signal_20977 ;
    wire new_AGEMA_signal_20978 ;
    wire new_AGEMA_signal_20979 ;
    wire new_AGEMA_signal_20980 ;
    wire new_AGEMA_signal_20981 ;
    wire new_AGEMA_signal_20982 ;
    wire new_AGEMA_signal_20983 ;
    wire new_AGEMA_signal_20984 ;
    wire new_AGEMA_signal_20985 ;
    wire new_AGEMA_signal_20986 ;
    wire new_AGEMA_signal_20987 ;
    wire new_AGEMA_signal_20988 ;
    wire new_AGEMA_signal_20989 ;
    wire new_AGEMA_signal_20990 ;
    wire new_AGEMA_signal_20991 ;
    wire new_AGEMA_signal_20992 ;
    wire new_AGEMA_signal_20993 ;
    wire new_AGEMA_signal_20994 ;
    wire new_AGEMA_signal_20995 ;
    wire new_AGEMA_signal_20996 ;
    wire new_AGEMA_signal_20997 ;
    wire new_AGEMA_signal_20998 ;
    wire new_AGEMA_signal_20999 ;
    wire new_AGEMA_signal_21000 ;
    wire new_AGEMA_signal_21001 ;
    wire new_AGEMA_signal_21002 ;
    wire new_AGEMA_signal_21003 ;
    wire new_AGEMA_signal_21004 ;
    wire new_AGEMA_signal_21005 ;
    wire new_AGEMA_signal_21006 ;
    wire new_AGEMA_signal_21007 ;
    wire new_AGEMA_signal_21008 ;
    wire new_AGEMA_signal_21009 ;
    wire new_AGEMA_signal_21010 ;
    wire new_AGEMA_signal_21011 ;
    wire new_AGEMA_signal_21012 ;
    wire new_AGEMA_signal_21013 ;
    wire new_AGEMA_signal_21014 ;
    wire new_AGEMA_signal_21015 ;
    wire new_AGEMA_signal_21016 ;
    wire new_AGEMA_signal_21017 ;
    wire new_AGEMA_signal_21018 ;
    wire new_AGEMA_signal_21019 ;
    wire new_AGEMA_signal_21020 ;
    wire new_AGEMA_signal_21021 ;
    wire new_AGEMA_signal_21022 ;
    wire new_AGEMA_signal_21023 ;
    wire new_AGEMA_signal_21024 ;
    wire new_AGEMA_signal_21025 ;
    wire new_AGEMA_signal_21026 ;
    wire new_AGEMA_signal_21027 ;
    wire new_AGEMA_signal_21028 ;
    wire new_AGEMA_signal_21029 ;
    wire new_AGEMA_signal_21030 ;
    wire new_AGEMA_signal_21031 ;
    wire new_AGEMA_signal_21032 ;
    wire new_AGEMA_signal_21033 ;
    wire new_AGEMA_signal_21034 ;
    wire new_AGEMA_signal_21035 ;
    wire new_AGEMA_signal_21036 ;
    wire new_AGEMA_signal_21037 ;
    wire new_AGEMA_signal_21038 ;
    wire new_AGEMA_signal_21039 ;
    wire new_AGEMA_signal_21040 ;
    wire new_AGEMA_signal_21041 ;
    wire new_AGEMA_signal_21042 ;
    wire new_AGEMA_signal_21043 ;
    wire new_AGEMA_signal_21044 ;
    wire new_AGEMA_signal_21045 ;
    wire new_AGEMA_signal_21046 ;
    wire new_AGEMA_signal_21047 ;
    wire new_AGEMA_signal_21048 ;
    wire new_AGEMA_signal_21049 ;
    wire new_AGEMA_signal_21050 ;
    wire new_AGEMA_signal_21051 ;
    wire new_AGEMA_signal_21052 ;
    wire new_AGEMA_signal_21053 ;
    wire new_AGEMA_signal_21054 ;
    wire new_AGEMA_signal_21055 ;
    wire new_AGEMA_signal_21056 ;
    wire new_AGEMA_signal_21057 ;
    wire new_AGEMA_signal_21058 ;
    wire new_AGEMA_signal_21059 ;
    wire new_AGEMA_signal_21060 ;
    wire new_AGEMA_signal_21061 ;
    wire new_AGEMA_signal_21062 ;
    wire new_AGEMA_signal_21063 ;
    wire new_AGEMA_signal_21064 ;
    wire new_AGEMA_signal_21065 ;
    wire new_AGEMA_signal_21066 ;
    wire new_AGEMA_signal_21067 ;
    wire new_AGEMA_signal_21068 ;
    wire new_AGEMA_signal_21069 ;
    wire new_AGEMA_signal_21070 ;
    wire new_AGEMA_signal_21071 ;
    wire new_AGEMA_signal_21072 ;
    wire new_AGEMA_signal_21073 ;
    wire new_AGEMA_signal_21074 ;
    wire new_AGEMA_signal_21075 ;
    wire new_AGEMA_signal_21076 ;
    wire new_AGEMA_signal_21077 ;
    wire new_AGEMA_signal_21078 ;
    wire new_AGEMA_signal_21079 ;
    wire new_AGEMA_signal_21080 ;
    wire new_AGEMA_signal_21081 ;
    wire new_AGEMA_signal_21082 ;
    wire new_AGEMA_signal_21083 ;
    wire new_AGEMA_signal_21084 ;
    wire new_AGEMA_signal_21085 ;
    wire new_AGEMA_signal_21086 ;
    wire new_AGEMA_signal_21087 ;
    wire new_AGEMA_signal_21088 ;
    wire new_AGEMA_signal_21089 ;
    wire new_AGEMA_signal_21090 ;
    wire new_AGEMA_signal_21091 ;
    wire new_AGEMA_signal_21092 ;
    wire new_AGEMA_signal_21093 ;
    wire new_AGEMA_signal_21094 ;
    wire new_AGEMA_signal_21095 ;
    wire new_AGEMA_signal_21096 ;
    wire new_AGEMA_signal_21097 ;
    wire new_AGEMA_signal_21098 ;
    wire new_AGEMA_signal_21099 ;
    wire new_AGEMA_signal_21100 ;
    wire new_AGEMA_signal_21101 ;
    wire new_AGEMA_signal_21102 ;
    wire new_AGEMA_signal_21103 ;
    wire new_AGEMA_signal_21104 ;
    wire new_AGEMA_signal_21105 ;
    wire new_AGEMA_signal_21106 ;
    wire new_AGEMA_signal_21107 ;
    wire new_AGEMA_signal_21108 ;
    wire new_AGEMA_signal_21109 ;
    wire new_AGEMA_signal_21110 ;
    wire new_AGEMA_signal_21111 ;
    wire new_AGEMA_signal_21112 ;
    wire new_AGEMA_signal_21113 ;
    wire new_AGEMA_signal_21114 ;
    wire new_AGEMA_signal_21115 ;
    wire new_AGEMA_signal_21116 ;
    wire new_AGEMA_signal_21117 ;
    wire new_AGEMA_signal_21118 ;
    wire new_AGEMA_signal_21119 ;
    wire new_AGEMA_signal_21120 ;
    wire new_AGEMA_signal_21121 ;
    wire new_AGEMA_signal_21122 ;
    wire new_AGEMA_signal_21123 ;
    wire new_AGEMA_signal_21124 ;
    wire new_AGEMA_signal_21125 ;
    wire new_AGEMA_signal_21126 ;
    wire new_AGEMA_signal_21127 ;
    wire new_AGEMA_signal_21128 ;
    wire new_AGEMA_signal_21129 ;
    wire new_AGEMA_signal_21130 ;
    wire new_AGEMA_signal_21131 ;
    wire new_AGEMA_signal_21132 ;
    wire new_AGEMA_signal_21133 ;
    wire new_AGEMA_signal_21134 ;
    wire new_AGEMA_signal_21135 ;
    wire new_AGEMA_signal_21136 ;
    wire new_AGEMA_signal_21137 ;
    wire new_AGEMA_signal_21138 ;
    wire new_AGEMA_signal_21139 ;
    wire new_AGEMA_signal_21140 ;
    wire new_AGEMA_signal_21141 ;
    wire new_AGEMA_signal_21142 ;
    wire new_AGEMA_signal_21143 ;
    wire new_AGEMA_signal_21144 ;
    wire new_AGEMA_signal_21145 ;
    wire new_AGEMA_signal_21146 ;
    wire new_AGEMA_signal_21147 ;
    wire new_AGEMA_signal_21148 ;
    wire new_AGEMA_signal_21149 ;
    wire new_AGEMA_signal_21150 ;
    wire new_AGEMA_signal_21151 ;
    wire new_AGEMA_signal_21152 ;
    wire new_AGEMA_signal_21153 ;
    wire new_AGEMA_signal_21154 ;
    wire new_AGEMA_signal_21155 ;
    wire new_AGEMA_signal_21156 ;
    wire new_AGEMA_signal_21157 ;
    wire new_AGEMA_signal_21158 ;
    wire new_AGEMA_signal_21159 ;
    wire new_AGEMA_signal_21160 ;
    wire new_AGEMA_signal_21161 ;
    wire new_AGEMA_signal_21162 ;
    wire new_AGEMA_signal_21163 ;
    wire new_AGEMA_signal_21164 ;
    wire new_AGEMA_signal_21165 ;
    wire new_AGEMA_signal_21166 ;
    wire new_AGEMA_signal_21167 ;
    wire new_AGEMA_signal_21168 ;
    wire new_AGEMA_signal_21169 ;
    wire new_AGEMA_signal_21170 ;
    wire new_AGEMA_signal_21171 ;
    wire new_AGEMA_signal_21172 ;
    wire new_AGEMA_signal_21173 ;
    wire new_AGEMA_signal_21174 ;
    wire new_AGEMA_signal_21175 ;
    wire new_AGEMA_signal_21176 ;
    wire new_AGEMA_signal_21177 ;
    wire new_AGEMA_signal_21178 ;
    wire new_AGEMA_signal_21179 ;
    wire new_AGEMA_signal_21180 ;
    wire new_AGEMA_signal_21181 ;
    wire new_AGEMA_signal_21182 ;
    wire new_AGEMA_signal_21183 ;
    wire new_AGEMA_signal_21184 ;
    wire new_AGEMA_signal_21185 ;
    wire new_AGEMA_signal_21186 ;
    wire new_AGEMA_signal_21187 ;
    wire new_AGEMA_signal_21188 ;
    wire new_AGEMA_signal_21189 ;
    wire new_AGEMA_signal_21190 ;
    wire new_AGEMA_signal_21191 ;
    wire new_AGEMA_signal_21192 ;
    wire new_AGEMA_signal_21193 ;
    wire new_AGEMA_signal_21194 ;
    wire new_AGEMA_signal_21195 ;
    wire new_AGEMA_signal_21196 ;
    wire new_AGEMA_signal_21197 ;
    wire new_AGEMA_signal_21198 ;
    wire new_AGEMA_signal_21199 ;
    wire new_AGEMA_signal_21200 ;
    wire new_AGEMA_signal_21201 ;
    wire new_AGEMA_signal_21202 ;
    wire new_AGEMA_signal_21203 ;
    wire new_AGEMA_signal_21204 ;
    wire new_AGEMA_signal_21205 ;
    wire new_AGEMA_signal_21206 ;
    wire new_AGEMA_signal_21207 ;
    wire new_AGEMA_signal_21208 ;
    wire new_AGEMA_signal_21209 ;
    wire new_AGEMA_signal_21210 ;
    wire new_AGEMA_signal_21211 ;
    wire new_AGEMA_signal_21212 ;
    wire new_AGEMA_signal_21213 ;
    wire new_AGEMA_signal_21214 ;
    wire new_AGEMA_signal_21215 ;
    wire new_AGEMA_signal_21216 ;
    wire new_AGEMA_signal_21217 ;
    wire new_AGEMA_signal_21218 ;
    wire new_AGEMA_signal_21219 ;
    wire new_AGEMA_signal_21220 ;
    wire new_AGEMA_signal_21221 ;
    wire new_AGEMA_signal_21222 ;
    wire new_AGEMA_signal_21223 ;
    wire new_AGEMA_signal_21224 ;
    wire new_AGEMA_signal_21225 ;
    wire new_AGEMA_signal_21226 ;
    wire new_AGEMA_signal_21227 ;
    wire new_AGEMA_signal_21228 ;
    wire new_AGEMA_signal_21229 ;
    wire new_AGEMA_signal_21230 ;
    wire new_AGEMA_signal_21231 ;
    wire new_AGEMA_signal_21232 ;
    wire new_AGEMA_signal_21233 ;
    wire new_AGEMA_signal_21234 ;
    wire new_AGEMA_signal_21235 ;
    wire new_AGEMA_signal_21236 ;
    wire new_AGEMA_signal_21237 ;
    wire new_AGEMA_signal_21238 ;
    wire new_AGEMA_signal_21239 ;
    wire new_AGEMA_signal_21240 ;
    wire new_AGEMA_signal_21241 ;
    wire new_AGEMA_signal_21242 ;
    wire new_AGEMA_signal_21243 ;
    wire new_AGEMA_signal_21244 ;
    wire new_AGEMA_signal_21245 ;
    wire new_AGEMA_signal_21246 ;
    wire new_AGEMA_signal_21247 ;
    wire new_AGEMA_signal_21248 ;
    wire new_AGEMA_signal_21249 ;
    wire new_AGEMA_signal_21250 ;
    wire new_AGEMA_signal_21251 ;
    wire new_AGEMA_signal_21252 ;
    wire new_AGEMA_signal_21253 ;
    wire new_AGEMA_signal_21254 ;
    wire new_AGEMA_signal_21255 ;
    wire new_AGEMA_signal_21256 ;
    wire new_AGEMA_signal_21257 ;
    wire new_AGEMA_signal_21258 ;
    wire new_AGEMA_signal_21259 ;
    wire new_AGEMA_signal_21260 ;
    wire new_AGEMA_signal_21261 ;
    wire new_AGEMA_signal_21262 ;
    wire new_AGEMA_signal_21263 ;
    wire new_AGEMA_signal_21264 ;
    wire new_AGEMA_signal_21265 ;
    wire new_AGEMA_signal_21266 ;
    wire new_AGEMA_signal_21267 ;
    wire new_AGEMA_signal_21268 ;
    wire new_AGEMA_signal_21269 ;
    wire new_AGEMA_signal_21270 ;
    wire new_AGEMA_signal_21271 ;
    wire new_AGEMA_signal_21272 ;
    wire new_AGEMA_signal_21273 ;
    wire new_AGEMA_signal_21274 ;
    wire new_AGEMA_signal_21275 ;
    wire new_AGEMA_signal_21276 ;
    wire new_AGEMA_signal_21277 ;
    wire new_AGEMA_signal_21278 ;
    wire new_AGEMA_signal_21279 ;
    wire new_AGEMA_signal_21280 ;
    wire new_AGEMA_signal_21281 ;
    wire new_AGEMA_signal_21282 ;
    wire new_AGEMA_signal_21283 ;
    wire new_AGEMA_signal_21284 ;
    wire new_AGEMA_signal_21285 ;
    wire new_AGEMA_signal_21286 ;
    wire new_AGEMA_signal_21287 ;
    wire new_AGEMA_signal_21288 ;
    wire new_AGEMA_signal_21289 ;
    wire new_AGEMA_signal_21290 ;
    wire new_AGEMA_signal_21291 ;
    wire new_AGEMA_signal_21292 ;
    wire new_AGEMA_signal_21293 ;
    wire new_AGEMA_signal_21294 ;
    wire new_AGEMA_signal_21295 ;
    wire new_AGEMA_signal_21296 ;
    wire new_AGEMA_signal_21297 ;
    wire new_AGEMA_signal_21298 ;
    wire new_AGEMA_signal_21299 ;
    wire new_AGEMA_signal_21300 ;
    wire new_AGEMA_signal_21301 ;
    wire new_AGEMA_signal_21302 ;
    wire new_AGEMA_signal_21303 ;
    wire new_AGEMA_signal_21304 ;
    wire new_AGEMA_signal_21305 ;
    wire new_AGEMA_signal_21306 ;
    wire new_AGEMA_signal_21307 ;
    wire new_AGEMA_signal_21308 ;
    wire new_AGEMA_signal_21309 ;
    wire new_AGEMA_signal_21310 ;
    wire new_AGEMA_signal_21311 ;
    wire new_AGEMA_signal_21312 ;
    wire new_AGEMA_signal_21313 ;
    wire new_AGEMA_signal_21314 ;
    wire new_AGEMA_signal_21315 ;
    wire new_AGEMA_signal_21316 ;
    wire new_AGEMA_signal_21317 ;
    wire new_AGEMA_signal_21318 ;
    wire new_AGEMA_signal_21319 ;
    wire new_AGEMA_signal_21320 ;
    wire new_AGEMA_signal_21321 ;
    wire new_AGEMA_signal_21322 ;
    wire new_AGEMA_signal_21323 ;
    wire new_AGEMA_signal_21324 ;
    wire new_AGEMA_signal_21325 ;
    wire new_AGEMA_signal_21326 ;
    wire new_AGEMA_signal_21327 ;
    wire new_AGEMA_signal_21328 ;
    wire new_AGEMA_signal_21329 ;
    wire new_AGEMA_signal_21330 ;
    wire new_AGEMA_signal_21331 ;
    wire new_AGEMA_signal_21332 ;
    wire new_AGEMA_signal_21333 ;
    wire new_AGEMA_signal_21334 ;
    wire new_AGEMA_signal_21335 ;
    wire new_AGEMA_signal_21336 ;
    wire new_AGEMA_signal_21337 ;
    wire new_AGEMA_signal_21338 ;
    wire new_AGEMA_signal_21339 ;
    wire new_AGEMA_signal_21340 ;
    wire new_AGEMA_signal_21341 ;
    wire new_AGEMA_signal_21342 ;
    wire new_AGEMA_signal_21343 ;
    wire new_AGEMA_signal_21344 ;
    wire new_AGEMA_signal_21345 ;
    wire new_AGEMA_signal_21346 ;
    wire new_AGEMA_signal_21347 ;
    wire new_AGEMA_signal_21348 ;
    wire new_AGEMA_signal_21349 ;
    wire new_AGEMA_signal_21350 ;
    wire new_AGEMA_signal_21351 ;
    wire new_AGEMA_signal_21352 ;
    wire new_AGEMA_signal_21353 ;
    wire new_AGEMA_signal_21354 ;
    wire new_AGEMA_signal_21355 ;
    wire new_AGEMA_signal_21356 ;
    wire new_AGEMA_signal_21357 ;
    wire new_AGEMA_signal_21358 ;
    wire new_AGEMA_signal_21359 ;
    wire new_AGEMA_signal_21360 ;
    wire new_AGEMA_signal_21361 ;
    wire new_AGEMA_signal_21362 ;
    wire new_AGEMA_signal_21363 ;
    wire new_AGEMA_signal_21364 ;
    wire new_AGEMA_signal_21365 ;
    wire new_AGEMA_signal_21366 ;
    wire new_AGEMA_signal_21367 ;
    wire new_AGEMA_signal_21368 ;
    wire new_AGEMA_signal_21369 ;
    wire new_AGEMA_signal_21370 ;
    wire new_AGEMA_signal_21371 ;
    wire new_AGEMA_signal_21372 ;
    wire new_AGEMA_signal_21373 ;
    wire new_AGEMA_signal_21374 ;
    wire new_AGEMA_signal_21375 ;
    wire new_AGEMA_signal_21376 ;
    wire new_AGEMA_signal_21377 ;
    wire new_AGEMA_signal_21378 ;
    wire new_AGEMA_signal_21379 ;
    wire new_AGEMA_signal_21380 ;
    wire new_AGEMA_signal_21381 ;
    wire new_AGEMA_signal_21382 ;
    wire new_AGEMA_signal_21383 ;
    wire new_AGEMA_signal_21384 ;
    wire new_AGEMA_signal_21385 ;
    wire new_AGEMA_signal_21386 ;
    wire new_AGEMA_signal_21387 ;
    wire new_AGEMA_signal_21388 ;
    wire new_AGEMA_signal_21389 ;
    wire new_AGEMA_signal_21390 ;
    wire new_AGEMA_signal_21391 ;
    wire new_AGEMA_signal_21392 ;
    wire new_AGEMA_signal_21393 ;
    wire new_AGEMA_signal_21394 ;
    wire new_AGEMA_signal_21395 ;
    wire new_AGEMA_signal_21396 ;
    wire new_AGEMA_signal_21397 ;
    wire new_AGEMA_signal_21398 ;
    wire new_AGEMA_signal_21399 ;
    wire new_AGEMA_signal_21400 ;
    wire new_AGEMA_signal_21401 ;
    wire new_AGEMA_signal_21402 ;
    wire new_AGEMA_signal_21403 ;
    wire new_AGEMA_signal_21404 ;
    wire new_AGEMA_signal_21405 ;
    wire new_AGEMA_signal_21406 ;
    wire new_AGEMA_signal_21407 ;
    wire new_AGEMA_signal_21408 ;
    wire new_AGEMA_signal_21409 ;
    wire new_AGEMA_signal_21410 ;
    wire new_AGEMA_signal_21411 ;
    wire new_AGEMA_signal_21412 ;
    wire new_AGEMA_signal_21413 ;
    wire new_AGEMA_signal_21414 ;
    wire new_AGEMA_signal_21415 ;
    wire new_AGEMA_signal_21416 ;
    wire new_AGEMA_signal_21417 ;
    wire new_AGEMA_signal_21418 ;
    wire new_AGEMA_signal_21419 ;
    wire new_AGEMA_signal_21420 ;
    wire new_AGEMA_signal_21421 ;
    wire new_AGEMA_signal_21422 ;
    wire new_AGEMA_signal_21423 ;
    wire new_AGEMA_signal_21424 ;
    wire new_AGEMA_signal_21425 ;
    wire new_AGEMA_signal_21426 ;
    wire new_AGEMA_signal_21427 ;
    wire new_AGEMA_signal_21428 ;
    wire new_AGEMA_signal_21429 ;
    wire new_AGEMA_signal_21430 ;
    wire new_AGEMA_signal_21431 ;
    wire new_AGEMA_signal_21432 ;
    wire new_AGEMA_signal_21433 ;
    wire new_AGEMA_signal_21434 ;
    wire new_AGEMA_signal_21435 ;
    wire new_AGEMA_signal_21436 ;
    wire new_AGEMA_signal_21437 ;
    wire new_AGEMA_signal_21438 ;
    wire new_AGEMA_signal_21439 ;
    wire new_AGEMA_signal_21440 ;
    wire new_AGEMA_signal_21441 ;
    wire new_AGEMA_signal_21442 ;
    wire new_AGEMA_signal_21443 ;
    wire new_AGEMA_signal_21444 ;
    wire new_AGEMA_signal_21445 ;
    wire new_AGEMA_signal_21446 ;
    wire new_AGEMA_signal_21447 ;
    wire new_AGEMA_signal_21448 ;
    wire new_AGEMA_signal_21449 ;
    wire new_AGEMA_signal_21450 ;
    wire new_AGEMA_signal_21451 ;
    wire new_AGEMA_signal_21452 ;
    wire new_AGEMA_signal_21453 ;
    wire new_AGEMA_signal_21454 ;
    wire new_AGEMA_signal_21455 ;
    wire new_AGEMA_signal_21456 ;
    wire new_AGEMA_signal_21457 ;
    wire new_AGEMA_signal_21458 ;
    wire new_AGEMA_signal_21459 ;
    wire new_AGEMA_signal_21460 ;
    wire new_AGEMA_signal_21461 ;
    wire new_AGEMA_signal_21462 ;
    wire new_AGEMA_signal_21463 ;
    wire new_AGEMA_signal_21464 ;
    wire new_AGEMA_signal_21465 ;
    wire new_AGEMA_signal_21466 ;
    wire new_AGEMA_signal_21467 ;
    wire new_AGEMA_signal_21468 ;
    wire new_AGEMA_signal_21469 ;
    wire new_AGEMA_signal_21470 ;
    wire new_AGEMA_signal_21471 ;
    wire new_AGEMA_signal_21472 ;
    wire new_AGEMA_signal_21473 ;
    wire new_AGEMA_signal_21474 ;
    wire new_AGEMA_signal_21475 ;
    wire new_AGEMA_signal_21476 ;
    wire new_AGEMA_signal_21477 ;
    wire new_AGEMA_signal_21478 ;
    wire new_AGEMA_signal_21479 ;
    wire new_AGEMA_signal_21480 ;
    wire new_AGEMA_signal_21481 ;
    wire new_AGEMA_signal_21482 ;
    wire new_AGEMA_signal_21483 ;
    wire new_AGEMA_signal_21484 ;
    wire new_AGEMA_signal_21485 ;
    wire new_AGEMA_signal_21486 ;
    wire new_AGEMA_signal_21487 ;
    wire new_AGEMA_signal_21488 ;
    wire new_AGEMA_signal_21489 ;
    wire new_AGEMA_signal_21490 ;
    wire new_AGEMA_signal_21491 ;
    wire new_AGEMA_signal_21492 ;
    wire new_AGEMA_signal_21493 ;
    wire new_AGEMA_signal_21494 ;
    wire new_AGEMA_signal_21495 ;
    wire new_AGEMA_signal_21496 ;
    wire new_AGEMA_signal_21497 ;
    wire new_AGEMA_signal_21498 ;
    wire new_AGEMA_signal_21499 ;
    wire new_AGEMA_signal_21500 ;
    wire new_AGEMA_signal_21501 ;
    wire new_AGEMA_signal_21502 ;
    wire new_AGEMA_signal_21503 ;
    wire new_AGEMA_signal_21504 ;
    wire new_AGEMA_signal_21505 ;
    wire new_AGEMA_signal_21506 ;
    wire new_AGEMA_signal_21507 ;
    wire new_AGEMA_signal_21508 ;
    wire new_AGEMA_signal_21509 ;
    wire new_AGEMA_signal_21510 ;
    wire new_AGEMA_signal_21511 ;
    wire new_AGEMA_signal_21512 ;
    wire new_AGEMA_signal_21513 ;
    wire new_AGEMA_signal_21514 ;
    wire new_AGEMA_signal_21515 ;
    wire new_AGEMA_signal_21516 ;
    wire new_AGEMA_signal_21517 ;
    wire new_AGEMA_signal_21518 ;
    wire new_AGEMA_signal_21519 ;
    wire new_AGEMA_signal_21520 ;
    wire new_AGEMA_signal_21521 ;
    wire new_AGEMA_signal_21522 ;
    wire new_AGEMA_signal_21523 ;
    wire new_AGEMA_signal_21524 ;
    wire new_AGEMA_signal_21525 ;
    wire new_AGEMA_signal_21526 ;
    wire new_AGEMA_signal_21527 ;
    wire new_AGEMA_signal_21528 ;
    wire new_AGEMA_signal_21529 ;
    wire new_AGEMA_signal_21530 ;
    wire new_AGEMA_signal_21531 ;
    wire new_AGEMA_signal_21532 ;
    wire new_AGEMA_signal_21533 ;
    wire new_AGEMA_signal_21534 ;
    wire new_AGEMA_signal_21535 ;
    wire new_AGEMA_signal_21536 ;
    wire new_AGEMA_signal_21537 ;
    wire new_AGEMA_signal_21538 ;
    wire new_AGEMA_signal_21539 ;
    wire new_AGEMA_signal_21540 ;
    wire new_AGEMA_signal_21541 ;
    wire new_AGEMA_signal_21542 ;
    wire new_AGEMA_signal_21543 ;
    wire new_AGEMA_signal_21544 ;
    wire new_AGEMA_signal_21545 ;
    wire new_AGEMA_signal_21546 ;
    wire new_AGEMA_signal_21547 ;
    wire new_AGEMA_signal_21548 ;
    wire new_AGEMA_signal_21549 ;
    wire new_AGEMA_signal_21550 ;
    wire new_AGEMA_signal_21551 ;
    wire new_AGEMA_signal_21552 ;
    wire new_AGEMA_signal_21553 ;
    wire new_AGEMA_signal_21554 ;
    wire new_AGEMA_signal_21555 ;
    wire new_AGEMA_signal_21556 ;
    wire new_AGEMA_signal_21557 ;
    wire new_AGEMA_signal_21558 ;
    wire new_AGEMA_signal_21559 ;
    wire new_AGEMA_signal_21560 ;
    wire new_AGEMA_signal_21561 ;
    wire new_AGEMA_signal_21562 ;
    wire new_AGEMA_signal_21563 ;
    wire new_AGEMA_signal_21564 ;
    wire new_AGEMA_signal_21565 ;
    wire new_AGEMA_signal_21566 ;
    wire new_AGEMA_signal_21567 ;
    wire new_AGEMA_signal_21568 ;
    wire new_AGEMA_signal_21569 ;
    wire new_AGEMA_signal_21570 ;
    wire new_AGEMA_signal_21571 ;
    wire new_AGEMA_signal_21572 ;
    wire new_AGEMA_signal_21573 ;
    wire new_AGEMA_signal_21574 ;
    wire new_AGEMA_signal_21575 ;
    wire new_AGEMA_signal_21576 ;
    wire new_AGEMA_signal_21577 ;
    wire new_AGEMA_signal_21578 ;
    wire new_AGEMA_signal_21579 ;
    wire new_AGEMA_signal_21580 ;
    wire new_AGEMA_signal_21581 ;
    wire new_AGEMA_signal_21582 ;
    wire new_AGEMA_signal_21583 ;
    wire new_AGEMA_signal_21584 ;
    wire new_AGEMA_signal_21585 ;
    wire new_AGEMA_signal_21586 ;
    wire new_AGEMA_signal_21587 ;
    wire new_AGEMA_signal_21588 ;
    wire new_AGEMA_signal_21589 ;
    wire new_AGEMA_signal_21590 ;
    wire new_AGEMA_signal_21591 ;
    wire new_AGEMA_signal_21592 ;
    wire new_AGEMA_signal_21593 ;
    wire new_AGEMA_signal_21594 ;
    wire new_AGEMA_signal_21595 ;
    wire new_AGEMA_signal_21596 ;
    wire new_AGEMA_signal_21597 ;
    wire new_AGEMA_signal_21598 ;
    wire new_AGEMA_signal_21599 ;
    wire new_AGEMA_signal_21600 ;
    wire new_AGEMA_signal_21601 ;
    wire new_AGEMA_signal_21602 ;
    wire new_AGEMA_signal_21603 ;
    wire new_AGEMA_signal_21604 ;
    wire new_AGEMA_signal_21605 ;
    wire new_AGEMA_signal_21606 ;
    wire new_AGEMA_signal_21607 ;
    wire new_AGEMA_signal_21608 ;
    wire new_AGEMA_signal_21609 ;
    wire new_AGEMA_signal_21610 ;
    wire new_AGEMA_signal_21611 ;
    wire new_AGEMA_signal_21612 ;
    wire new_AGEMA_signal_21613 ;
    wire new_AGEMA_signal_21614 ;
    wire new_AGEMA_signal_21615 ;
    wire new_AGEMA_signal_21616 ;
    wire new_AGEMA_signal_21617 ;
    wire new_AGEMA_signal_21618 ;
    wire new_AGEMA_signal_21619 ;
    wire new_AGEMA_signal_21620 ;
    wire new_AGEMA_signal_21621 ;
    wire new_AGEMA_signal_21622 ;
    wire new_AGEMA_signal_21623 ;
    wire new_AGEMA_signal_21624 ;
    wire new_AGEMA_signal_21625 ;
    wire new_AGEMA_signal_21626 ;
    wire new_AGEMA_signal_21627 ;
    wire new_AGEMA_signal_21628 ;
    wire new_AGEMA_signal_21629 ;
    wire new_AGEMA_signal_21630 ;
    wire new_AGEMA_signal_21631 ;
    wire new_AGEMA_signal_21632 ;
    wire new_AGEMA_signal_21633 ;
    wire new_AGEMA_signal_21634 ;
    wire new_AGEMA_signal_21635 ;
    wire new_AGEMA_signal_21636 ;
    wire new_AGEMA_signal_21637 ;
    wire new_AGEMA_signal_21638 ;
    wire new_AGEMA_signal_21639 ;
    wire new_AGEMA_signal_21640 ;
    wire new_AGEMA_signal_21641 ;
    wire new_AGEMA_signal_21642 ;
    wire new_AGEMA_signal_21643 ;
    wire new_AGEMA_signal_21644 ;
    wire new_AGEMA_signal_21645 ;
    wire new_AGEMA_signal_21646 ;
    wire new_AGEMA_signal_21647 ;
    wire new_AGEMA_signal_21648 ;
    wire new_AGEMA_signal_21649 ;
    wire new_AGEMA_signal_21650 ;
    wire new_AGEMA_signal_21651 ;
    wire new_AGEMA_signal_21652 ;
    wire new_AGEMA_signal_21653 ;
    wire new_AGEMA_signal_21654 ;
    wire new_AGEMA_signal_21655 ;
    wire new_AGEMA_signal_21656 ;
    wire new_AGEMA_signal_21657 ;
    wire new_AGEMA_signal_21658 ;
    wire new_AGEMA_signal_21659 ;
    wire new_AGEMA_signal_21660 ;
    wire new_AGEMA_signal_21661 ;
    wire new_AGEMA_signal_21662 ;
    wire new_AGEMA_signal_21663 ;
    wire new_AGEMA_signal_21664 ;
    wire new_AGEMA_signal_21665 ;
    wire new_AGEMA_signal_21666 ;
    wire new_AGEMA_signal_21667 ;
    wire new_AGEMA_signal_21668 ;
    wire new_AGEMA_signal_21669 ;
    wire new_AGEMA_signal_21670 ;
    wire new_AGEMA_signal_21671 ;
    wire new_AGEMA_signal_21672 ;
    wire new_AGEMA_signal_21673 ;
    wire new_AGEMA_signal_21674 ;
    wire new_AGEMA_signal_21675 ;
    wire new_AGEMA_signal_21676 ;
    wire new_AGEMA_signal_21677 ;
    wire new_AGEMA_signal_21678 ;
    wire new_AGEMA_signal_21679 ;
    wire new_AGEMA_signal_21680 ;
    wire new_AGEMA_signal_21681 ;
    wire new_AGEMA_signal_21682 ;
    wire new_AGEMA_signal_21683 ;
    wire new_AGEMA_signal_21684 ;
    wire new_AGEMA_signal_21685 ;
    wire new_AGEMA_signal_21686 ;
    wire new_AGEMA_signal_21687 ;
    wire new_AGEMA_signal_21688 ;
    wire new_AGEMA_signal_21689 ;
    wire new_AGEMA_signal_21690 ;
    wire new_AGEMA_signal_21691 ;
    wire new_AGEMA_signal_21692 ;
    wire new_AGEMA_signal_21693 ;
    wire new_AGEMA_signal_21694 ;
    wire new_AGEMA_signal_21695 ;
    wire new_AGEMA_signal_21696 ;
    wire new_AGEMA_signal_21697 ;
    wire new_AGEMA_signal_21698 ;
    wire new_AGEMA_signal_21699 ;
    wire new_AGEMA_signal_21700 ;
    wire new_AGEMA_signal_21701 ;
    wire new_AGEMA_signal_21702 ;
    wire new_AGEMA_signal_21703 ;
    wire new_AGEMA_signal_21704 ;
    wire new_AGEMA_signal_21705 ;
    wire new_AGEMA_signal_21706 ;
    wire new_AGEMA_signal_21707 ;
    wire new_AGEMA_signal_21708 ;
    wire new_AGEMA_signal_21709 ;
    wire new_AGEMA_signal_21710 ;
    wire new_AGEMA_signal_21711 ;
    wire new_AGEMA_signal_21712 ;
    wire new_AGEMA_signal_21713 ;
    wire new_AGEMA_signal_21714 ;
    wire new_AGEMA_signal_21715 ;
    wire new_AGEMA_signal_21716 ;
    wire new_AGEMA_signal_21717 ;
    wire new_AGEMA_signal_21718 ;
    wire new_AGEMA_signal_21719 ;
    wire new_AGEMA_signal_21720 ;
    wire new_AGEMA_signal_21721 ;
    wire new_AGEMA_signal_21722 ;
    wire new_AGEMA_signal_21723 ;
    wire new_AGEMA_signal_21724 ;
    wire new_AGEMA_signal_21725 ;
    wire new_AGEMA_signal_21726 ;
    wire new_AGEMA_signal_21727 ;
    wire new_AGEMA_signal_21728 ;
    wire new_AGEMA_signal_21729 ;
    wire new_AGEMA_signal_21730 ;
    wire new_AGEMA_signal_21731 ;
    wire new_AGEMA_signal_21732 ;
    wire new_AGEMA_signal_21733 ;
    wire new_AGEMA_signal_21734 ;
    wire new_AGEMA_signal_21735 ;
    wire new_AGEMA_signal_21736 ;
    wire new_AGEMA_signal_21737 ;
    wire new_AGEMA_signal_21738 ;
    wire new_AGEMA_signal_21739 ;
    wire new_AGEMA_signal_21740 ;
    wire new_AGEMA_signal_21741 ;
    wire new_AGEMA_signal_21742 ;
    wire new_AGEMA_signal_21743 ;
    wire new_AGEMA_signal_21744 ;
    wire new_AGEMA_signal_21745 ;
    wire new_AGEMA_signal_21746 ;
    wire new_AGEMA_signal_21747 ;
    wire new_AGEMA_signal_21748 ;
    wire new_AGEMA_signal_21749 ;
    wire new_AGEMA_signal_21750 ;
    wire new_AGEMA_signal_21751 ;
    wire new_AGEMA_signal_21752 ;
    wire new_AGEMA_signal_21753 ;
    wire new_AGEMA_signal_21754 ;
    wire new_AGEMA_signal_21755 ;
    wire new_AGEMA_signal_21756 ;
    wire new_AGEMA_signal_21757 ;
    wire new_AGEMA_signal_21758 ;
    wire new_AGEMA_signal_21759 ;
    wire new_AGEMA_signal_21760 ;
    wire new_AGEMA_signal_21761 ;
    wire new_AGEMA_signal_21762 ;
    wire new_AGEMA_signal_21763 ;
    wire new_AGEMA_signal_21764 ;
    wire new_AGEMA_signal_21765 ;
    wire new_AGEMA_signal_21766 ;
    wire new_AGEMA_signal_21767 ;
    wire new_AGEMA_signal_21768 ;
    wire new_AGEMA_signal_21769 ;
    wire new_AGEMA_signal_21770 ;
    wire new_AGEMA_signal_21771 ;
    wire new_AGEMA_signal_21772 ;
    wire new_AGEMA_signal_21773 ;
    wire new_AGEMA_signal_21774 ;
    wire new_AGEMA_signal_21775 ;
    wire new_AGEMA_signal_21776 ;
    wire new_AGEMA_signal_21777 ;
    wire new_AGEMA_signal_21778 ;
    wire new_AGEMA_signal_21779 ;
    wire new_AGEMA_signal_21780 ;
    wire new_AGEMA_signal_21781 ;
    wire new_AGEMA_signal_21782 ;
    wire new_AGEMA_signal_21783 ;
    wire new_AGEMA_signal_21784 ;
    wire new_AGEMA_signal_21785 ;
    wire new_AGEMA_signal_21786 ;
    wire new_AGEMA_signal_21787 ;
    wire new_AGEMA_signal_21788 ;
    wire new_AGEMA_signal_21789 ;
    wire new_AGEMA_signal_21790 ;
    wire new_AGEMA_signal_21791 ;
    wire new_AGEMA_signal_21792 ;
    wire new_AGEMA_signal_21793 ;
    wire new_AGEMA_signal_21794 ;
    wire new_AGEMA_signal_21795 ;
    wire new_AGEMA_signal_21796 ;
    wire new_AGEMA_signal_21797 ;
    wire new_AGEMA_signal_21798 ;
    wire new_AGEMA_signal_21799 ;
    wire new_AGEMA_signal_21800 ;
    wire new_AGEMA_signal_21801 ;
    wire new_AGEMA_signal_21802 ;
    wire new_AGEMA_signal_21803 ;
    wire new_AGEMA_signal_21804 ;
    wire new_AGEMA_signal_21805 ;
    wire new_AGEMA_signal_21806 ;
    wire new_AGEMA_signal_21807 ;
    wire new_AGEMA_signal_21808 ;
    wire new_AGEMA_signal_21809 ;
    wire new_AGEMA_signal_21810 ;
    wire new_AGEMA_signal_21811 ;
    wire new_AGEMA_signal_21812 ;
    wire new_AGEMA_signal_21813 ;
    wire new_AGEMA_signal_21814 ;
    wire new_AGEMA_signal_21815 ;
    wire new_AGEMA_signal_21816 ;
    wire new_AGEMA_signal_21817 ;
    wire new_AGEMA_signal_21818 ;
    wire new_AGEMA_signal_21819 ;
    wire new_AGEMA_signal_21820 ;
    wire new_AGEMA_signal_21821 ;
    wire new_AGEMA_signal_21822 ;
    wire new_AGEMA_signal_21823 ;
    wire new_AGEMA_signal_21824 ;
    wire new_AGEMA_signal_21825 ;
    wire new_AGEMA_signal_21826 ;
    wire new_AGEMA_signal_21827 ;
    wire new_AGEMA_signal_21828 ;
    wire new_AGEMA_signal_21829 ;
    wire new_AGEMA_signal_21830 ;
    wire new_AGEMA_signal_21831 ;
    wire new_AGEMA_signal_21832 ;
    wire new_AGEMA_signal_21833 ;
    wire new_AGEMA_signal_21834 ;
    wire new_AGEMA_signal_21835 ;
    wire new_AGEMA_signal_21836 ;
    wire new_AGEMA_signal_21837 ;
    wire new_AGEMA_signal_21838 ;
    wire new_AGEMA_signal_21839 ;
    wire new_AGEMA_signal_21840 ;
    wire new_AGEMA_signal_21841 ;
    wire new_AGEMA_signal_21842 ;
    wire new_AGEMA_signal_21843 ;
    wire new_AGEMA_signal_21844 ;
    wire new_AGEMA_signal_21845 ;
    wire new_AGEMA_signal_21846 ;
    wire new_AGEMA_signal_21847 ;
    wire new_AGEMA_signal_21848 ;
    wire new_AGEMA_signal_21849 ;
    wire new_AGEMA_signal_21850 ;
    wire new_AGEMA_signal_21851 ;
    wire new_AGEMA_signal_21852 ;
    wire new_AGEMA_signal_21853 ;
    wire new_AGEMA_signal_21854 ;
    wire new_AGEMA_signal_21855 ;
    wire new_AGEMA_signal_21856 ;
    wire new_AGEMA_signal_21857 ;
    wire new_AGEMA_signal_21858 ;
    wire new_AGEMA_signal_21859 ;
    wire new_AGEMA_signal_21860 ;
    wire new_AGEMA_signal_21861 ;
    wire new_AGEMA_signal_21862 ;
    wire new_AGEMA_signal_21863 ;
    wire new_AGEMA_signal_21864 ;
    wire new_AGEMA_signal_21865 ;
    wire new_AGEMA_signal_21866 ;
    wire new_AGEMA_signal_21867 ;
    wire new_AGEMA_signal_21868 ;
    wire new_AGEMA_signal_21869 ;
    wire new_AGEMA_signal_21870 ;
    wire new_AGEMA_signal_21871 ;
    wire new_AGEMA_signal_21872 ;
    wire new_AGEMA_signal_21873 ;
    wire new_AGEMA_signal_21874 ;
    wire new_AGEMA_signal_21875 ;
    wire new_AGEMA_signal_21876 ;
    wire new_AGEMA_signal_21877 ;
    wire new_AGEMA_signal_21878 ;
    wire new_AGEMA_signal_21879 ;
    wire new_AGEMA_signal_21880 ;
    wire new_AGEMA_signal_21881 ;
    wire new_AGEMA_signal_21882 ;
    wire new_AGEMA_signal_21883 ;
    wire new_AGEMA_signal_21884 ;
    wire new_AGEMA_signal_21885 ;
    wire new_AGEMA_signal_21886 ;
    wire new_AGEMA_signal_21887 ;
    wire new_AGEMA_signal_21888 ;
    wire new_AGEMA_signal_21889 ;
    wire new_AGEMA_signal_21890 ;
    wire new_AGEMA_signal_21891 ;
    wire new_AGEMA_signal_21892 ;
    wire new_AGEMA_signal_21893 ;
    wire new_AGEMA_signal_21894 ;
    wire new_AGEMA_signal_21895 ;
    wire new_AGEMA_signal_21896 ;
    wire new_AGEMA_signal_21897 ;
    wire new_AGEMA_signal_21898 ;
    wire new_AGEMA_signal_21899 ;
    wire new_AGEMA_signal_21900 ;
    wire new_AGEMA_signal_21901 ;
    wire new_AGEMA_signal_21902 ;
    wire new_AGEMA_signal_21903 ;
    wire new_AGEMA_signal_21904 ;
    wire new_AGEMA_signal_21905 ;
    wire new_AGEMA_signal_21906 ;
    wire new_AGEMA_signal_21907 ;
    wire new_AGEMA_signal_21908 ;
    wire new_AGEMA_signal_21909 ;
    wire new_AGEMA_signal_21910 ;
    wire new_AGEMA_signal_21911 ;
    wire new_AGEMA_signal_21912 ;
    wire new_AGEMA_signal_21913 ;
    wire new_AGEMA_signal_21914 ;
    wire new_AGEMA_signal_21915 ;
    wire new_AGEMA_signal_21916 ;
    wire new_AGEMA_signal_21917 ;
    wire new_AGEMA_signal_21918 ;
    wire new_AGEMA_signal_21919 ;
    wire new_AGEMA_signal_21920 ;
    wire new_AGEMA_signal_21921 ;
    wire new_AGEMA_signal_21922 ;
    wire new_AGEMA_signal_21923 ;
    wire new_AGEMA_signal_21924 ;
    wire new_AGEMA_signal_21925 ;
    wire new_AGEMA_signal_21926 ;
    wire new_AGEMA_signal_21927 ;
    wire new_AGEMA_signal_21928 ;
    wire new_AGEMA_signal_21929 ;
    wire new_AGEMA_signal_21930 ;
    wire new_AGEMA_signal_21931 ;
    wire new_AGEMA_signal_21932 ;
    wire new_AGEMA_signal_21933 ;
    wire new_AGEMA_signal_21934 ;
    wire new_AGEMA_signal_21935 ;
    wire new_AGEMA_signal_21936 ;
    wire new_AGEMA_signal_21937 ;
    wire new_AGEMA_signal_21938 ;
    wire new_AGEMA_signal_21939 ;
    wire new_AGEMA_signal_21940 ;
    wire new_AGEMA_signal_21941 ;
    wire new_AGEMA_signal_21942 ;
    wire new_AGEMA_signal_21943 ;
    wire new_AGEMA_signal_21944 ;
    wire new_AGEMA_signal_21945 ;
    wire new_AGEMA_signal_21946 ;
    wire new_AGEMA_signal_21947 ;
    wire new_AGEMA_signal_21948 ;
    wire new_AGEMA_signal_21949 ;
    wire new_AGEMA_signal_21950 ;
    wire new_AGEMA_signal_21951 ;
    wire new_AGEMA_signal_21952 ;
    wire new_AGEMA_signal_21953 ;
    wire new_AGEMA_signal_21954 ;
    wire new_AGEMA_signal_21955 ;
    wire new_AGEMA_signal_21956 ;
    wire new_AGEMA_signal_21957 ;
    wire new_AGEMA_signal_21958 ;
    wire new_AGEMA_signal_21959 ;
    wire new_AGEMA_signal_21960 ;
    wire new_AGEMA_signal_21961 ;
    wire new_AGEMA_signal_21962 ;
    wire new_AGEMA_signal_21963 ;
    wire new_AGEMA_signal_21964 ;
    wire new_AGEMA_signal_21965 ;
    wire new_AGEMA_signal_21966 ;
    wire new_AGEMA_signal_21967 ;
    wire new_AGEMA_signal_21968 ;
    wire new_AGEMA_signal_21969 ;
    wire new_AGEMA_signal_21970 ;
    wire new_AGEMA_signal_21971 ;
    wire new_AGEMA_signal_21972 ;
    wire new_AGEMA_signal_21973 ;
    wire new_AGEMA_signal_21974 ;
    wire new_AGEMA_signal_21975 ;
    wire new_AGEMA_signal_21976 ;
    wire new_AGEMA_signal_21977 ;
    wire new_AGEMA_signal_21978 ;
    wire new_AGEMA_signal_21979 ;
    wire new_AGEMA_signal_21980 ;
    wire new_AGEMA_signal_21981 ;
    wire new_AGEMA_signal_21982 ;
    wire new_AGEMA_signal_21983 ;
    wire new_AGEMA_signal_21984 ;
    wire new_AGEMA_signal_21985 ;
    wire new_AGEMA_signal_21986 ;
    wire new_AGEMA_signal_21987 ;
    wire new_AGEMA_signal_21988 ;
    wire new_AGEMA_signal_21989 ;
    wire new_AGEMA_signal_21990 ;
    wire new_AGEMA_signal_21991 ;
    wire new_AGEMA_signal_21992 ;
    wire new_AGEMA_signal_21993 ;
    wire new_AGEMA_signal_21994 ;
    wire new_AGEMA_signal_21995 ;
    wire new_AGEMA_signal_21996 ;
    wire new_AGEMA_signal_21997 ;
    wire new_AGEMA_signal_21998 ;
    wire new_AGEMA_signal_21999 ;
    wire new_AGEMA_signal_22000 ;
    wire new_AGEMA_signal_22001 ;
    wire new_AGEMA_signal_22002 ;
    wire new_AGEMA_signal_22003 ;
    wire new_AGEMA_signal_22004 ;
    wire new_AGEMA_signal_22005 ;
    wire new_AGEMA_signal_22006 ;
    wire new_AGEMA_signal_22007 ;
    wire new_AGEMA_signal_22008 ;
    wire new_AGEMA_signal_22009 ;
    wire new_AGEMA_signal_22010 ;
    wire new_AGEMA_signal_22011 ;
    wire new_AGEMA_signal_22012 ;
    wire new_AGEMA_signal_22013 ;
    wire new_AGEMA_signal_22014 ;
    wire new_AGEMA_signal_22015 ;
    wire new_AGEMA_signal_22016 ;
    wire new_AGEMA_signal_22017 ;
    wire new_AGEMA_signal_22018 ;
    wire new_AGEMA_signal_22019 ;
    wire new_AGEMA_signal_22020 ;
    wire new_AGEMA_signal_22021 ;
    wire new_AGEMA_signal_22022 ;
    wire new_AGEMA_signal_22023 ;
    wire new_AGEMA_signal_22024 ;
    wire new_AGEMA_signal_22025 ;
    wire new_AGEMA_signal_22026 ;
    wire new_AGEMA_signal_22027 ;
    wire new_AGEMA_signal_22028 ;
    wire new_AGEMA_signal_22029 ;
    wire new_AGEMA_signal_22030 ;
    wire new_AGEMA_signal_22031 ;
    wire new_AGEMA_signal_22032 ;
    wire new_AGEMA_signal_22033 ;
    wire new_AGEMA_signal_22034 ;
    wire new_AGEMA_signal_22035 ;
    wire new_AGEMA_signal_22036 ;
    wire new_AGEMA_signal_22037 ;
    wire new_AGEMA_signal_22038 ;
    wire new_AGEMA_signal_22039 ;
    wire new_AGEMA_signal_22040 ;
    wire new_AGEMA_signal_22041 ;
    wire new_AGEMA_signal_22042 ;
    wire new_AGEMA_signal_22043 ;
    wire new_AGEMA_signal_22044 ;
    wire new_AGEMA_signal_22045 ;
    wire new_AGEMA_signal_22046 ;
    wire new_AGEMA_signal_22047 ;
    wire new_AGEMA_signal_22048 ;
    wire new_AGEMA_signal_22049 ;
    wire new_AGEMA_signal_22050 ;
    wire new_AGEMA_signal_22051 ;
    wire new_AGEMA_signal_22052 ;
    wire new_AGEMA_signal_22053 ;
    wire new_AGEMA_signal_22054 ;
    wire new_AGEMA_signal_22055 ;
    wire new_AGEMA_signal_22056 ;
    wire new_AGEMA_signal_22057 ;
    wire new_AGEMA_signal_22058 ;
    wire new_AGEMA_signal_22059 ;
    wire new_AGEMA_signal_22060 ;
    wire new_AGEMA_signal_22061 ;
    wire new_AGEMA_signal_22062 ;
    wire new_AGEMA_signal_22063 ;
    wire new_AGEMA_signal_22064 ;
    wire new_AGEMA_signal_22065 ;
    wire new_AGEMA_signal_22066 ;
    wire new_AGEMA_signal_22067 ;
    wire new_AGEMA_signal_22068 ;
    wire new_AGEMA_signal_22069 ;
    wire new_AGEMA_signal_22070 ;
    wire new_AGEMA_signal_22071 ;
    wire new_AGEMA_signal_22072 ;
    wire new_AGEMA_signal_22073 ;
    wire new_AGEMA_signal_22074 ;
    wire new_AGEMA_signal_22075 ;
    wire new_AGEMA_signal_22076 ;
    wire new_AGEMA_signal_22077 ;
    wire new_AGEMA_signal_22078 ;
    wire new_AGEMA_signal_22079 ;
    wire new_AGEMA_signal_22080 ;
    wire new_AGEMA_signal_22081 ;
    wire new_AGEMA_signal_22082 ;
    wire new_AGEMA_signal_22083 ;
    wire new_AGEMA_signal_22084 ;
    wire new_AGEMA_signal_22085 ;
    wire new_AGEMA_signal_22086 ;
    wire new_AGEMA_signal_22087 ;
    wire new_AGEMA_signal_22088 ;
    wire new_AGEMA_signal_22089 ;
    wire new_AGEMA_signal_22090 ;
    wire new_AGEMA_signal_22091 ;
    wire new_AGEMA_signal_22092 ;
    wire new_AGEMA_signal_22093 ;
    wire new_AGEMA_signal_22094 ;
    wire new_AGEMA_signal_22095 ;
    wire new_AGEMA_signal_22096 ;
    wire new_AGEMA_signal_22097 ;
    wire new_AGEMA_signal_22098 ;
    wire new_AGEMA_signal_22099 ;
    wire new_AGEMA_signal_22100 ;
    wire new_AGEMA_signal_22101 ;
    wire new_AGEMA_signal_22102 ;
    wire new_AGEMA_signal_22103 ;
    wire new_AGEMA_signal_22104 ;
    wire new_AGEMA_signal_22105 ;
    wire new_AGEMA_signal_22106 ;
    wire new_AGEMA_signal_22107 ;
    wire new_AGEMA_signal_22108 ;
    wire new_AGEMA_signal_22109 ;
    wire new_AGEMA_signal_22110 ;
    wire new_AGEMA_signal_22111 ;
    wire new_AGEMA_signal_22112 ;
    wire new_AGEMA_signal_22113 ;
    wire new_AGEMA_signal_22114 ;
    wire new_AGEMA_signal_22115 ;
    wire new_AGEMA_signal_22116 ;
    wire new_AGEMA_signal_22117 ;
    wire new_AGEMA_signal_22118 ;
    wire new_AGEMA_signal_22119 ;
    wire new_AGEMA_signal_22120 ;
    wire new_AGEMA_signal_22121 ;
    wire new_AGEMA_signal_22122 ;
    wire new_AGEMA_signal_22123 ;
    wire new_AGEMA_signal_22124 ;
    wire new_AGEMA_signal_22125 ;
    wire new_AGEMA_signal_22126 ;
    wire new_AGEMA_signal_22127 ;
    wire new_AGEMA_signal_22128 ;
    wire new_AGEMA_signal_22129 ;
    wire new_AGEMA_signal_22130 ;
    wire new_AGEMA_signal_22131 ;
    wire new_AGEMA_signal_22132 ;
    wire new_AGEMA_signal_22133 ;
    wire new_AGEMA_signal_22134 ;
    wire new_AGEMA_signal_22135 ;
    wire new_AGEMA_signal_22136 ;
    wire new_AGEMA_signal_22137 ;
    wire new_AGEMA_signal_22138 ;
    wire new_AGEMA_signal_22139 ;
    wire new_AGEMA_signal_22140 ;
    wire new_AGEMA_signal_22141 ;
    wire new_AGEMA_signal_22142 ;
    wire new_AGEMA_signal_22143 ;
    wire new_AGEMA_signal_22144 ;
    wire new_AGEMA_signal_22145 ;
    wire new_AGEMA_signal_22146 ;
    wire new_AGEMA_signal_22147 ;
    wire new_AGEMA_signal_22148 ;
    wire new_AGEMA_signal_22149 ;
    wire new_AGEMA_signal_22150 ;
    wire new_AGEMA_signal_22151 ;
    wire new_AGEMA_signal_22152 ;
    wire new_AGEMA_signal_22153 ;
    wire new_AGEMA_signal_22154 ;
    wire new_AGEMA_signal_22155 ;
    wire new_AGEMA_signal_22156 ;
    wire new_AGEMA_signal_22157 ;
    wire new_AGEMA_signal_22158 ;
    wire new_AGEMA_signal_22159 ;
    wire new_AGEMA_signal_22160 ;
    wire new_AGEMA_signal_22161 ;
    wire new_AGEMA_signal_22162 ;
    wire new_AGEMA_signal_22163 ;
    wire new_AGEMA_signal_22164 ;
    wire new_AGEMA_signal_22165 ;
    wire new_AGEMA_signal_22166 ;
    wire new_AGEMA_signal_22167 ;
    wire new_AGEMA_signal_22168 ;
    wire new_AGEMA_signal_22169 ;
    wire new_AGEMA_signal_22170 ;
    wire new_AGEMA_signal_22171 ;
    wire new_AGEMA_signal_22172 ;
    wire new_AGEMA_signal_22173 ;
    wire new_AGEMA_signal_22174 ;
    wire new_AGEMA_signal_22175 ;
    wire new_AGEMA_signal_22176 ;
    wire new_AGEMA_signal_22177 ;
    wire new_AGEMA_signal_22178 ;
    wire new_AGEMA_signal_22179 ;
    wire new_AGEMA_signal_22180 ;
    wire new_AGEMA_signal_22181 ;
    wire new_AGEMA_signal_22182 ;
    wire new_AGEMA_signal_22183 ;
    wire new_AGEMA_signal_22184 ;
    wire new_AGEMA_signal_22185 ;
    wire new_AGEMA_signal_22186 ;
    wire new_AGEMA_signal_22187 ;
    wire new_AGEMA_signal_22188 ;
    wire new_AGEMA_signal_22189 ;
    wire new_AGEMA_signal_22190 ;
    wire new_AGEMA_signal_22191 ;
    wire new_AGEMA_signal_22192 ;
    wire new_AGEMA_signal_22193 ;
    wire new_AGEMA_signal_22194 ;
    wire new_AGEMA_signal_22195 ;
    wire new_AGEMA_signal_22196 ;
    wire new_AGEMA_signal_22197 ;
    wire new_AGEMA_signal_22198 ;
    wire new_AGEMA_signal_22199 ;
    wire new_AGEMA_signal_22200 ;
    wire new_AGEMA_signal_22201 ;
    wire new_AGEMA_signal_22202 ;
    wire new_AGEMA_signal_22203 ;
    wire new_AGEMA_signal_22204 ;
    wire new_AGEMA_signal_22205 ;
    wire new_AGEMA_signal_22206 ;
    wire new_AGEMA_signal_22207 ;
    wire new_AGEMA_signal_22208 ;
    wire new_AGEMA_signal_22209 ;
    wire new_AGEMA_signal_22210 ;
    wire new_AGEMA_signal_22211 ;
    wire new_AGEMA_signal_22212 ;
    wire new_AGEMA_signal_22213 ;
    wire new_AGEMA_signal_22214 ;
    wire new_AGEMA_signal_22215 ;
    wire new_AGEMA_signal_22216 ;
    wire new_AGEMA_signal_22217 ;
    wire new_AGEMA_signal_22218 ;
    wire new_AGEMA_signal_22219 ;
    wire new_AGEMA_signal_22220 ;
    wire new_AGEMA_signal_22221 ;
    wire new_AGEMA_signal_22222 ;
    wire new_AGEMA_signal_22223 ;
    wire new_AGEMA_signal_22224 ;
    wire new_AGEMA_signal_22225 ;
    wire new_AGEMA_signal_22226 ;
    wire new_AGEMA_signal_22227 ;
    wire new_AGEMA_signal_22228 ;
    wire new_AGEMA_signal_22229 ;
    wire new_AGEMA_signal_22230 ;
    wire new_AGEMA_signal_22231 ;
    wire new_AGEMA_signal_22232 ;
    wire new_AGEMA_signal_22233 ;
    wire new_AGEMA_signal_22234 ;
    wire new_AGEMA_signal_22235 ;
    wire new_AGEMA_signal_22236 ;
    wire new_AGEMA_signal_22237 ;
    wire new_AGEMA_signal_22238 ;
    wire new_AGEMA_signal_22239 ;
    wire new_AGEMA_signal_22240 ;
    wire new_AGEMA_signal_22241 ;
    wire new_AGEMA_signal_22242 ;
    wire new_AGEMA_signal_22243 ;
    wire new_AGEMA_signal_22244 ;
    wire new_AGEMA_signal_22245 ;
    wire new_AGEMA_signal_22246 ;
    wire new_AGEMA_signal_22247 ;
    wire new_AGEMA_signal_22248 ;
    wire new_AGEMA_signal_22249 ;
    wire new_AGEMA_signal_22250 ;
    wire new_AGEMA_signal_22251 ;
    wire new_AGEMA_signal_22252 ;
    wire new_AGEMA_signal_22253 ;
    wire new_AGEMA_signal_22254 ;
    wire new_AGEMA_signal_22255 ;
    wire new_AGEMA_signal_22256 ;
    wire new_AGEMA_signal_22257 ;
    wire new_AGEMA_signal_22258 ;
    wire new_AGEMA_signal_22259 ;
    wire new_AGEMA_signal_22260 ;
    wire new_AGEMA_signal_22261 ;
    wire new_AGEMA_signal_22262 ;
    wire new_AGEMA_signal_22263 ;
    wire new_AGEMA_signal_22264 ;
    wire new_AGEMA_signal_22265 ;
    wire new_AGEMA_signal_22266 ;
    wire new_AGEMA_signal_22267 ;
    wire new_AGEMA_signal_22268 ;
    wire new_AGEMA_signal_22269 ;
    wire new_AGEMA_signal_22270 ;
    wire new_AGEMA_signal_22271 ;
    wire new_AGEMA_signal_22272 ;
    wire new_AGEMA_signal_22273 ;
    wire new_AGEMA_signal_22274 ;
    wire new_AGEMA_signal_22275 ;
    wire new_AGEMA_signal_22276 ;
    wire new_AGEMA_signal_22277 ;
    wire new_AGEMA_signal_22278 ;
    wire new_AGEMA_signal_22279 ;
    wire new_AGEMA_signal_22280 ;
    wire new_AGEMA_signal_22281 ;
    wire new_AGEMA_signal_22282 ;
    wire new_AGEMA_signal_22283 ;
    wire new_AGEMA_signal_22284 ;
    wire new_AGEMA_signal_22285 ;
    wire new_AGEMA_signal_22286 ;
    wire new_AGEMA_signal_22287 ;
    wire new_AGEMA_signal_22288 ;
    wire new_AGEMA_signal_22289 ;
    wire new_AGEMA_signal_22290 ;
    wire new_AGEMA_signal_22291 ;
    wire new_AGEMA_signal_22292 ;
    wire new_AGEMA_signal_22293 ;
    wire new_AGEMA_signal_22294 ;
    wire new_AGEMA_signal_22295 ;
    wire new_AGEMA_signal_22296 ;
    wire new_AGEMA_signal_22297 ;
    wire new_AGEMA_signal_22298 ;
    wire new_AGEMA_signal_22299 ;
    wire new_AGEMA_signal_22300 ;
    wire new_AGEMA_signal_22301 ;
    wire new_AGEMA_signal_22302 ;
    wire new_AGEMA_signal_22303 ;
    wire new_AGEMA_signal_22304 ;
    wire new_AGEMA_signal_22305 ;
    wire new_AGEMA_signal_22306 ;
    wire new_AGEMA_signal_22307 ;
    wire new_AGEMA_signal_22308 ;
    wire new_AGEMA_signal_22309 ;
    wire new_AGEMA_signal_22310 ;
    wire new_AGEMA_signal_22311 ;
    wire new_AGEMA_signal_22312 ;
    wire new_AGEMA_signal_22313 ;
    wire new_AGEMA_signal_22314 ;
    wire new_AGEMA_signal_22315 ;
    wire new_AGEMA_signal_22316 ;
    wire new_AGEMA_signal_22317 ;
    wire new_AGEMA_signal_22318 ;
    wire new_AGEMA_signal_22319 ;
    wire new_AGEMA_signal_22320 ;
    wire new_AGEMA_signal_22321 ;
    wire new_AGEMA_signal_22322 ;
    wire new_AGEMA_signal_22323 ;
    wire new_AGEMA_signal_22324 ;
    wire new_AGEMA_signal_22325 ;
    wire new_AGEMA_signal_22326 ;
    wire new_AGEMA_signal_22327 ;
    wire new_AGEMA_signal_22328 ;
    wire new_AGEMA_signal_22329 ;
    wire new_AGEMA_signal_22330 ;
    wire new_AGEMA_signal_22331 ;
    wire new_AGEMA_signal_22332 ;
    wire new_AGEMA_signal_22333 ;
    wire new_AGEMA_signal_22334 ;
    wire new_AGEMA_signal_22335 ;
    wire new_AGEMA_signal_22336 ;
    wire new_AGEMA_signal_22337 ;
    wire new_AGEMA_signal_22338 ;
    wire new_AGEMA_signal_22339 ;
    wire new_AGEMA_signal_22340 ;
    wire new_AGEMA_signal_22341 ;
    wire new_AGEMA_signal_22342 ;
    wire new_AGEMA_signal_22343 ;
    wire new_AGEMA_signal_22344 ;
    wire new_AGEMA_signal_22345 ;
    wire new_AGEMA_signal_22346 ;
    wire new_AGEMA_signal_22347 ;
    wire new_AGEMA_signal_22348 ;
    wire new_AGEMA_signal_22349 ;
    wire new_AGEMA_signal_22350 ;
    wire new_AGEMA_signal_22351 ;
    wire new_AGEMA_signal_22352 ;
    wire new_AGEMA_signal_22353 ;
    wire new_AGEMA_signal_22354 ;
    wire new_AGEMA_signal_22355 ;
    wire new_AGEMA_signal_22356 ;
    wire new_AGEMA_signal_22357 ;
    wire new_AGEMA_signal_22358 ;
    wire new_AGEMA_signal_22359 ;
    wire new_AGEMA_signal_22360 ;
    wire new_AGEMA_signal_22361 ;
    wire new_AGEMA_signal_22362 ;
    wire new_AGEMA_signal_22363 ;
    wire new_AGEMA_signal_22364 ;
    wire new_AGEMA_signal_22365 ;
    wire new_AGEMA_signal_22366 ;
    wire new_AGEMA_signal_22367 ;
    wire new_AGEMA_signal_22368 ;
    wire new_AGEMA_signal_22369 ;
    wire new_AGEMA_signal_22370 ;
    wire new_AGEMA_signal_22371 ;
    wire new_AGEMA_signal_22372 ;
    wire new_AGEMA_signal_22373 ;
    wire new_AGEMA_signal_22374 ;
    wire new_AGEMA_signal_22375 ;
    wire new_AGEMA_signal_22376 ;
    wire new_AGEMA_signal_22377 ;
    wire new_AGEMA_signal_22378 ;
    wire new_AGEMA_signal_22379 ;
    wire new_AGEMA_signal_22380 ;
    wire new_AGEMA_signal_22381 ;
    wire new_AGEMA_signal_22382 ;
    wire new_AGEMA_signal_22383 ;
    wire new_AGEMA_signal_22384 ;
    wire new_AGEMA_signal_22385 ;
    wire new_AGEMA_signal_22386 ;
    wire new_AGEMA_signal_22387 ;
    wire new_AGEMA_signal_22388 ;
    wire new_AGEMA_signal_22389 ;
    wire new_AGEMA_signal_22390 ;
    wire new_AGEMA_signal_22391 ;
    wire new_AGEMA_signal_22392 ;
    wire new_AGEMA_signal_22393 ;
    wire new_AGEMA_signal_22394 ;
    wire new_AGEMA_signal_22395 ;
    wire new_AGEMA_signal_22396 ;
    wire new_AGEMA_signal_22397 ;
    wire new_AGEMA_signal_22398 ;
    wire new_AGEMA_signal_22399 ;
    wire new_AGEMA_signal_22400 ;
    wire new_AGEMA_signal_22401 ;
    wire new_AGEMA_signal_22402 ;
    wire new_AGEMA_signal_22403 ;
    wire new_AGEMA_signal_22404 ;
    wire new_AGEMA_signal_22405 ;
    wire new_AGEMA_signal_22406 ;
    wire new_AGEMA_signal_22407 ;
    wire new_AGEMA_signal_22408 ;
    wire new_AGEMA_signal_22409 ;
    wire new_AGEMA_signal_22410 ;
    wire new_AGEMA_signal_22411 ;
    wire new_AGEMA_signal_22412 ;
    wire new_AGEMA_signal_22413 ;
    wire new_AGEMA_signal_22414 ;
    wire new_AGEMA_signal_22415 ;
    wire new_AGEMA_signal_22416 ;
    wire new_AGEMA_signal_22417 ;
    wire new_AGEMA_signal_22418 ;
    wire new_AGEMA_signal_22419 ;
    wire new_AGEMA_signal_22420 ;
    wire new_AGEMA_signal_22421 ;
    wire new_AGEMA_signal_22422 ;
    wire new_AGEMA_signal_22423 ;
    wire new_AGEMA_signal_22424 ;
    wire new_AGEMA_signal_22425 ;
    wire new_AGEMA_signal_22426 ;
    wire new_AGEMA_signal_22427 ;
    wire new_AGEMA_signal_22428 ;
    wire new_AGEMA_signal_22429 ;
    wire new_AGEMA_signal_22430 ;
    wire new_AGEMA_signal_22431 ;
    wire new_AGEMA_signal_22432 ;
    wire new_AGEMA_signal_22433 ;
    wire new_AGEMA_signal_22434 ;
    wire new_AGEMA_signal_22435 ;
    wire new_AGEMA_signal_22436 ;
    wire new_AGEMA_signal_22437 ;
    wire new_AGEMA_signal_22438 ;
    wire new_AGEMA_signal_22439 ;
    wire new_AGEMA_signal_22440 ;
    wire new_AGEMA_signal_22441 ;
    wire new_AGEMA_signal_22442 ;
    wire new_AGEMA_signal_22443 ;
    wire new_AGEMA_signal_22444 ;
    wire new_AGEMA_signal_22445 ;
    wire new_AGEMA_signal_22446 ;
    wire new_AGEMA_signal_22447 ;
    wire new_AGEMA_signal_22448 ;
    wire new_AGEMA_signal_22449 ;
    wire new_AGEMA_signal_22450 ;
    wire new_AGEMA_signal_22451 ;
    wire new_AGEMA_signal_22452 ;
    wire new_AGEMA_signal_22453 ;
    wire new_AGEMA_signal_22454 ;
    wire new_AGEMA_signal_22455 ;
    wire new_AGEMA_signal_22456 ;
    wire new_AGEMA_signal_22457 ;
    wire new_AGEMA_signal_22458 ;
    wire new_AGEMA_signal_22459 ;
    wire new_AGEMA_signal_22460 ;
    wire new_AGEMA_signal_22461 ;
    wire new_AGEMA_signal_22462 ;
    wire new_AGEMA_signal_22463 ;
    wire new_AGEMA_signal_22464 ;
    wire new_AGEMA_signal_22465 ;
    wire new_AGEMA_signal_22466 ;
    wire new_AGEMA_signal_22467 ;
    wire new_AGEMA_signal_22468 ;
    wire new_AGEMA_signal_22469 ;
    wire new_AGEMA_signal_22470 ;
    wire new_AGEMA_signal_22471 ;
    wire new_AGEMA_signal_22472 ;
    wire new_AGEMA_signal_22473 ;
    wire new_AGEMA_signal_22474 ;
    wire new_AGEMA_signal_22475 ;
    wire new_AGEMA_signal_22476 ;
    wire new_AGEMA_signal_22477 ;
    wire new_AGEMA_signal_22478 ;
    wire new_AGEMA_signal_22479 ;
    wire new_AGEMA_signal_22480 ;
    wire new_AGEMA_signal_22481 ;
    wire new_AGEMA_signal_22482 ;
    wire new_AGEMA_signal_22483 ;
    wire new_AGEMA_signal_22484 ;
    wire new_AGEMA_signal_22485 ;
    wire new_AGEMA_signal_22486 ;
    wire new_AGEMA_signal_22487 ;
    wire new_AGEMA_signal_22488 ;
    wire new_AGEMA_signal_22489 ;
    wire new_AGEMA_signal_22490 ;
    wire new_AGEMA_signal_22491 ;
    wire new_AGEMA_signal_22492 ;
    wire new_AGEMA_signal_22493 ;
    wire new_AGEMA_signal_22494 ;
    wire new_AGEMA_signal_22495 ;
    wire new_AGEMA_signal_22496 ;
    wire new_AGEMA_signal_22497 ;
    wire new_AGEMA_signal_22498 ;
    wire new_AGEMA_signal_22499 ;
    wire new_AGEMA_signal_22500 ;
    wire new_AGEMA_signal_22501 ;
    wire new_AGEMA_signal_22502 ;
    wire new_AGEMA_signal_22503 ;
    wire new_AGEMA_signal_22504 ;
    wire new_AGEMA_signal_22505 ;
    wire new_AGEMA_signal_22506 ;
    wire new_AGEMA_signal_22507 ;
    wire new_AGEMA_signal_22508 ;
    wire new_AGEMA_signal_22509 ;
    wire new_AGEMA_signal_22510 ;
    wire new_AGEMA_signal_22511 ;
    wire new_AGEMA_signal_22512 ;
    wire new_AGEMA_signal_22513 ;
    wire new_AGEMA_signal_22514 ;
    wire new_AGEMA_signal_22515 ;
    wire new_AGEMA_signal_22516 ;
    wire new_AGEMA_signal_22517 ;
    wire new_AGEMA_signal_22518 ;
    wire new_AGEMA_signal_22519 ;
    wire new_AGEMA_signal_22520 ;
    wire new_AGEMA_signal_22521 ;
    wire new_AGEMA_signal_22522 ;
    wire new_AGEMA_signal_22523 ;
    wire new_AGEMA_signal_22524 ;
    wire new_AGEMA_signal_22525 ;
    wire new_AGEMA_signal_22526 ;
    wire new_AGEMA_signal_22527 ;
    wire new_AGEMA_signal_22528 ;
    wire new_AGEMA_signal_22529 ;
    wire new_AGEMA_signal_22530 ;
    wire new_AGEMA_signal_22531 ;
    wire new_AGEMA_signal_22532 ;
    wire new_AGEMA_signal_22533 ;
    wire new_AGEMA_signal_22534 ;
    wire new_AGEMA_signal_22535 ;
    wire new_AGEMA_signal_22536 ;
    wire new_AGEMA_signal_22537 ;
    wire new_AGEMA_signal_22538 ;
    wire new_AGEMA_signal_22539 ;
    wire new_AGEMA_signal_22540 ;
    wire new_AGEMA_signal_22541 ;
    wire new_AGEMA_signal_22542 ;
    wire new_AGEMA_signal_22543 ;
    wire new_AGEMA_signal_22544 ;
    wire new_AGEMA_signal_22545 ;
    wire new_AGEMA_signal_22546 ;
    wire new_AGEMA_signal_22547 ;
    wire new_AGEMA_signal_22548 ;
    wire new_AGEMA_signal_22549 ;
    wire new_AGEMA_signal_22550 ;
    wire new_AGEMA_signal_22551 ;
    wire new_AGEMA_signal_22552 ;
    wire new_AGEMA_signal_22553 ;
    wire new_AGEMA_signal_22554 ;
    wire new_AGEMA_signal_22555 ;
    wire new_AGEMA_signal_22556 ;
    wire new_AGEMA_signal_22557 ;
    wire new_AGEMA_signal_22558 ;
    wire new_AGEMA_signal_22559 ;
    wire new_AGEMA_signal_22560 ;
    wire new_AGEMA_signal_22561 ;
    wire new_AGEMA_signal_22562 ;
    wire new_AGEMA_signal_22563 ;
    wire new_AGEMA_signal_22564 ;
    wire new_AGEMA_signal_22565 ;
    wire new_AGEMA_signal_22566 ;
    wire new_AGEMA_signal_22567 ;
    wire new_AGEMA_signal_22568 ;
    wire new_AGEMA_signal_22569 ;
    wire new_AGEMA_signal_22570 ;
    wire new_AGEMA_signal_22571 ;
    wire new_AGEMA_signal_22572 ;
    wire new_AGEMA_signal_22573 ;
    wire new_AGEMA_signal_22574 ;
    wire new_AGEMA_signal_22575 ;
    wire new_AGEMA_signal_22576 ;
    wire new_AGEMA_signal_22577 ;
    wire new_AGEMA_signal_22578 ;
    wire new_AGEMA_signal_22579 ;
    wire new_AGEMA_signal_22580 ;
    wire new_AGEMA_signal_22581 ;
    wire new_AGEMA_signal_22582 ;
    wire new_AGEMA_signal_22583 ;
    wire new_AGEMA_signal_22584 ;
    wire new_AGEMA_signal_22585 ;
    wire new_AGEMA_signal_22586 ;
    wire new_AGEMA_signal_22587 ;
    wire new_AGEMA_signal_22588 ;
    wire new_AGEMA_signal_22589 ;
    wire new_AGEMA_signal_22590 ;
    wire new_AGEMA_signal_22591 ;
    wire new_AGEMA_signal_22592 ;
    wire new_AGEMA_signal_22593 ;
    wire new_AGEMA_signal_22594 ;
    wire new_AGEMA_signal_22595 ;
    wire new_AGEMA_signal_22596 ;
    wire new_AGEMA_signal_22597 ;
    wire new_AGEMA_signal_22598 ;
    wire new_AGEMA_signal_22599 ;
    wire new_AGEMA_signal_22600 ;
    wire new_AGEMA_signal_22601 ;
    wire new_AGEMA_signal_22602 ;
    wire new_AGEMA_signal_22603 ;
    wire new_AGEMA_signal_22604 ;
    wire new_AGEMA_signal_22605 ;
    wire new_AGEMA_signal_22606 ;
    wire new_AGEMA_signal_22607 ;
    wire new_AGEMA_signal_22608 ;
    wire new_AGEMA_signal_22609 ;
    wire new_AGEMA_signal_22610 ;
    wire new_AGEMA_signal_22611 ;
    wire new_AGEMA_signal_22612 ;
    wire new_AGEMA_signal_22613 ;
    wire new_AGEMA_signal_22614 ;
    wire new_AGEMA_signal_22615 ;
    wire new_AGEMA_signal_22616 ;
    wire new_AGEMA_signal_22617 ;
    wire new_AGEMA_signal_22618 ;
    wire new_AGEMA_signal_22619 ;
    wire new_AGEMA_signal_22620 ;
    wire new_AGEMA_signal_22621 ;
    wire new_AGEMA_signal_22622 ;
    wire new_AGEMA_signal_22623 ;
    wire new_AGEMA_signal_22624 ;
    wire new_AGEMA_signal_22625 ;
    wire new_AGEMA_signal_22626 ;
    wire new_AGEMA_signal_22627 ;
    wire new_AGEMA_signal_22628 ;
    wire new_AGEMA_signal_22629 ;
    wire new_AGEMA_signal_22630 ;
    wire new_AGEMA_signal_22631 ;
    wire new_AGEMA_signal_22632 ;
    wire new_AGEMA_signal_22633 ;
    wire new_AGEMA_signal_22634 ;
    wire new_AGEMA_signal_22635 ;
    wire new_AGEMA_signal_22636 ;
    wire new_AGEMA_signal_22637 ;
    wire new_AGEMA_signal_22638 ;
    wire new_AGEMA_signal_22639 ;
    wire new_AGEMA_signal_22640 ;
    wire new_AGEMA_signal_22641 ;
    wire new_AGEMA_signal_22642 ;
    wire new_AGEMA_signal_22643 ;
    wire new_AGEMA_signal_22644 ;
    wire new_AGEMA_signal_22645 ;
    wire new_AGEMA_signal_22646 ;
    wire new_AGEMA_signal_22647 ;
    wire new_AGEMA_signal_22648 ;
    wire new_AGEMA_signal_22649 ;
    wire new_AGEMA_signal_22650 ;
    wire new_AGEMA_signal_22651 ;
    wire new_AGEMA_signal_22652 ;
    wire new_AGEMA_signal_22653 ;
    wire new_AGEMA_signal_22654 ;
    wire new_AGEMA_signal_22655 ;
    wire new_AGEMA_signal_22656 ;
    wire new_AGEMA_signal_22657 ;
    wire new_AGEMA_signal_22658 ;
    wire new_AGEMA_signal_22659 ;
    wire new_AGEMA_signal_22660 ;
    wire new_AGEMA_signal_22661 ;
    wire new_AGEMA_signal_22662 ;
    wire new_AGEMA_signal_22663 ;
    wire new_AGEMA_signal_22664 ;
    wire new_AGEMA_signal_22665 ;
    wire new_AGEMA_signal_22666 ;
    wire new_AGEMA_signal_22667 ;
    wire new_AGEMA_signal_22668 ;
    wire new_AGEMA_signal_22669 ;
    wire new_AGEMA_signal_22670 ;
    wire new_AGEMA_signal_22671 ;
    wire new_AGEMA_signal_22672 ;
    wire new_AGEMA_signal_22673 ;
    wire new_AGEMA_signal_22674 ;
    wire new_AGEMA_signal_22675 ;
    wire new_AGEMA_signal_22676 ;
    wire new_AGEMA_signal_22677 ;
    wire new_AGEMA_signal_22678 ;
    wire new_AGEMA_signal_22679 ;
    wire new_AGEMA_signal_22680 ;
    wire new_AGEMA_signal_22681 ;
    wire new_AGEMA_signal_22682 ;
    wire new_AGEMA_signal_22683 ;
    wire new_AGEMA_signal_22684 ;
    wire new_AGEMA_signal_22685 ;
    wire new_AGEMA_signal_22686 ;
    wire new_AGEMA_signal_22687 ;
    wire new_AGEMA_signal_22688 ;
    wire new_AGEMA_signal_22689 ;
    wire new_AGEMA_signal_22690 ;
    wire new_AGEMA_signal_22691 ;
    wire new_AGEMA_signal_22692 ;
    wire new_AGEMA_signal_22693 ;
    wire new_AGEMA_signal_22694 ;
    wire new_AGEMA_signal_22695 ;
    wire new_AGEMA_signal_22696 ;
    wire new_AGEMA_signal_22697 ;
    wire new_AGEMA_signal_22698 ;
    wire new_AGEMA_signal_22699 ;
    wire new_AGEMA_signal_22700 ;
    wire new_AGEMA_signal_22701 ;
    wire new_AGEMA_signal_22702 ;
    wire new_AGEMA_signal_22703 ;
    wire new_AGEMA_signal_22704 ;
    wire new_AGEMA_signal_22705 ;
    wire new_AGEMA_signal_22706 ;
    wire new_AGEMA_signal_22707 ;
    wire new_AGEMA_signal_22708 ;
    wire new_AGEMA_signal_22709 ;
    wire new_AGEMA_signal_22710 ;
    wire new_AGEMA_signal_22711 ;
    wire new_AGEMA_signal_22712 ;
    wire new_AGEMA_signal_22713 ;
    wire new_AGEMA_signal_22714 ;
    wire new_AGEMA_signal_22715 ;
    wire new_AGEMA_signal_22716 ;
    wire new_AGEMA_signal_22717 ;
    wire new_AGEMA_signal_22718 ;
    wire new_AGEMA_signal_22719 ;
    wire new_AGEMA_signal_22720 ;
    wire new_AGEMA_signal_22721 ;
    wire new_AGEMA_signal_22722 ;
    wire new_AGEMA_signal_22723 ;
    wire new_AGEMA_signal_22724 ;
    wire new_AGEMA_signal_22725 ;
    wire new_AGEMA_signal_22726 ;
    wire new_AGEMA_signal_22727 ;
    wire new_AGEMA_signal_22728 ;
    wire new_AGEMA_signal_22729 ;
    wire new_AGEMA_signal_22730 ;
    wire new_AGEMA_signal_22731 ;
    wire new_AGEMA_signal_22732 ;
    wire new_AGEMA_signal_22733 ;
    wire new_AGEMA_signal_22734 ;
    wire new_AGEMA_signal_22735 ;
    wire new_AGEMA_signal_22736 ;
    wire new_AGEMA_signal_22737 ;
    wire new_AGEMA_signal_22738 ;
    wire new_AGEMA_signal_22739 ;
    wire new_AGEMA_signal_22740 ;
    wire new_AGEMA_signal_22741 ;
    wire new_AGEMA_signal_22742 ;
    wire new_AGEMA_signal_22743 ;
    wire new_AGEMA_signal_22744 ;
    wire new_AGEMA_signal_22745 ;
    wire new_AGEMA_signal_22746 ;
    wire new_AGEMA_signal_22747 ;
    wire new_AGEMA_signal_22748 ;
    wire new_AGEMA_signal_22749 ;
    wire new_AGEMA_signal_22750 ;
    wire new_AGEMA_signal_22751 ;
    wire new_AGEMA_signal_22752 ;
    wire new_AGEMA_signal_22753 ;
    wire new_AGEMA_signal_22754 ;
    wire new_AGEMA_signal_22755 ;
    wire new_AGEMA_signal_22756 ;
    wire new_AGEMA_signal_22757 ;
    wire new_AGEMA_signal_22758 ;
    wire new_AGEMA_signal_22759 ;
    wire new_AGEMA_signal_22760 ;
    wire new_AGEMA_signal_22761 ;
    wire new_AGEMA_signal_22762 ;
    wire new_AGEMA_signal_22763 ;
    wire new_AGEMA_signal_22764 ;
    wire new_AGEMA_signal_22765 ;
    wire new_AGEMA_signal_22766 ;
    wire new_AGEMA_signal_22767 ;
    wire new_AGEMA_signal_22768 ;
    wire new_AGEMA_signal_22769 ;
    wire new_AGEMA_signal_22770 ;
    wire new_AGEMA_signal_22771 ;
    wire new_AGEMA_signal_22772 ;
    wire new_AGEMA_signal_22773 ;
    wire new_AGEMA_signal_22774 ;
    wire new_AGEMA_signal_22775 ;
    wire new_AGEMA_signal_22776 ;
    wire new_AGEMA_signal_22777 ;
    wire new_AGEMA_signal_22778 ;
    wire new_AGEMA_signal_22779 ;
    wire new_AGEMA_signal_22780 ;
    wire new_AGEMA_signal_22781 ;
    wire new_AGEMA_signal_22782 ;
    wire new_AGEMA_signal_22783 ;
    wire new_AGEMA_signal_22784 ;
    wire new_AGEMA_signal_22785 ;
    wire new_AGEMA_signal_22786 ;
    wire new_AGEMA_signal_22787 ;
    wire new_AGEMA_signal_22788 ;
    wire new_AGEMA_signal_22789 ;
    wire new_AGEMA_signal_22790 ;
    wire new_AGEMA_signal_22791 ;
    wire new_AGEMA_signal_22792 ;
    wire new_AGEMA_signal_22793 ;
    wire new_AGEMA_signal_22794 ;
    wire new_AGEMA_signal_22795 ;
    wire new_AGEMA_signal_22796 ;
    wire new_AGEMA_signal_22797 ;
    wire new_AGEMA_signal_22798 ;
    wire new_AGEMA_signal_22799 ;
    wire new_AGEMA_signal_22800 ;
    wire new_AGEMA_signal_22801 ;
    wire new_AGEMA_signal_22802 ;
    wire new_AGEMA_signal_22803 ;
    wire new_AGEMA_signal_22804 ;
    wire new_AGEMA_signal_22805 ;
    wire new_AGEMA_signal_22806 ;
    wire new_AGEMA_signal_22807 ;
    wire new_AGEMA_signal_22808 ;
    wire new_AGEMA_signal_22809 ;
    wire new_AGEMA_signal_22810 ;
    wire new_AGEMA_signal_22811 ;
    wire new_AGEMA_signal_22812 ;
    wire new_AGEMA_signal_22813 ;
    wire new_AGEMA_signal_22814 ;
    wire new_AGEMA_signal_22815 ;
    wire new_AGEMA_signal_22816 ;
    wire new_AGEMA_signal_22817 ;
    wire new_AGEMA_signal_22818 ;
    wire new_AGEMA_signal_22819 ;
    wire new_AGEMA_signal_22820 ;
    wire new_AGEMA_signal_22821 ;
    wire new_AGEMA_signal_22822 ;
    wire new_AGEMA_signal_22823 ;
    wire new_AGEMA_signal_22824 ;
    wire new_AGEMA_signal_22825 ;
    wire new_AGEMA_signal_22826 ;
    wire new_AGEMA_signal_22827 ;
    wire new_AGEMA_signal_22828 ;
    wire new_AGEMA_signal_22829 ;
    wire new_AGEMA_signal_22830 ;
    wire new_AGEMA_signal_22831 ;
    wire new_AGEMA_signal_22832 ;
    wire new_AGEMA_signal_22833 ;
    wire new_AGEMA_signal_22834 ;
    wire new_AGEMA_signal_22835 ;
    wire new_AGEMA_signal_22836 ;
    wire new_AGEMA_signal_22837 ;
    wire new_AGEMA_signal_22838 ;
    wire new_AGEMA_signal_22839 ;
    wire new_AGEMA_signal_22840 ;
    wire new_AGEMA_signal_22841 ;
    wire new_AGEMA_signal_22842 ;
    wire new_AGEMA_signal_22843 ;
    wire new_AGEMA_signal_22844 ;
    wire new_AGEMA_signal_22845 ;
    wire new_AGEMA_signal_22846 ;
    wire new_AGEMA_signal_22847 ;
    wire new_AGEMA_signal_22848 ;
    wire new_AGEMA_signal_22849 ;
    wire new_AGEMA_signal_22850 ;
    wire new_AGEMA_signal_22851 ;
    wire new_AGEMA_signal_22852 ;
    wire new_AGEMA_signal_22853 ;
    wire new_AGEMA_signal_22854 ;
    wire new_AGEMA_signal_22855 ;
    wire new_AGEMA_signal_22856 ;
    wire new_AGEMA_signal_22857 ;
    wire new_AGEMA_signal_22858 ;
    wire new_AGEMA_signal_22859 ;
    wire new_AGEMA_signal_22860 ;
    wire new_AGEMA_signal_22861 ;
    wire new_AGEMA_signal_22862 ;
    wire new_AGEMA_signal_22863 ;
    wire new_AGEMA_signal_22864 ;
    wire new_AGEMA_signal_22865 ;
    wire new_AGEMA_signal_22866 ;
    wire new_AGEMA_signal_22867 ;
    wire new_AGEMA_signal_22868 ;
    wire new_AGEMA_signal_22869 ;
    wire new_AGEMA_signal_22870 ;
    wire new_AGEMA_signal_22871 ;
    wire new_AGEMA_signal_22872 ;
    wire new_AGEMA_signal_22873 ;
    wire new_AGEMA_signal_22874 ;
    wire new_AGEMA_signal_22875 ;
    wire new_AGEMA_signal_22876 ;
    wire new_AGEMA_signal_22877 ;
    wire new_AGEMA_signal_22878 ;
    wire new_AGEMA_signal_22879 ;
    wire new_AGEMA_signal_22880 ;
    wire new_AGEMA_signal_22881 ;
    wire new_AGEMA_signal_22882 ;
    wire new_AGEMA_signal_22883 ;
    wire new_AGEMA_signal_22884 ;
    wire new_AGEMA_signal_22885 ;
    wire new_AGEMA_signal_22886 ;
    wire new_AGEMA_signal_22887 ;
    wire new_AGEMA_signal_22888 ;
    wire new_AGEMA_signal_22889 ;
    wire new_AGEMA_signal_22890 ;
    wire new_AGEMA_signal_22891 ;
    wire new_AGEMA_signal_22892 ;
    wire new_AGEMA_signal_22893 ;
    wire new_AGEMA_signal_22894 ;
    wire new_AGEMA_signal_22895 ;
    wire new_AGEMA_signal_22896 ;
    wire new_AGEMA_signal_22897 ;
    wire new_AGEMA_signal_22898 ;
    wire new_AGEMA_signal_22899 ;
    wire new_AGEMA_signal_22900 ;
    wire new_AGEMA_signal_22901 ;
    wire new_AGEMA_signal_22902 ;
    wire new_AGEMA_signal_22903 ;
    wire new_AGEMA_signal_22904 ;
    wire new_AGEMA_signal_22905 ;
    wire new_AGEMA_signal_22906 ;
    wire new_AGEMA_signal_22907 ;
    wire new_AGEMA_signal_22908 ;
    wire new_AGEMA_signal_22909 ;
    wire new_AGEMA_signal_22910 ;
    wire new_AGEMA_signal_22911 ;
    wire new_AGEMA_signal_22912 ;
    wire new_AGEMA_signal_22913 ;
    wire new_AGEMA_signal_22914 ;
    wire new_AGEMA_signal_22915 ;
    wire new_AGEMA_signal_22916 ;
    wire new_AGEMA_signal_22917 ;
    wire new_AGEMA_signal_22918 ;
    wire new_AGEMA_signal_22919 ;
    wire new_AGEMA_signal_22920 ;
    wire new_AGEMA_signal_22921 ;
    wire new_AGEMA_signal_22922 ;
    wire new_AGEMA_signal_22923 ;
    wire new_AGEMA_signal_22924 ;
    wire new_AGEMA_signal_22925 ;
    wire new_AGEMA_signal_22926 ;
    wire new_AGEMA_signal_22927 ;
    wire new_AGEMA_signal_22928 ;
    wire new_AGEMA_signal_22929 ;
    wire new_AGEMA_signal_22930 ;
    wire new_AGEMA_signal_22931 ;
    wire new_AGEMA_signal_22932 ;
    wire new_AGEMA_signal_22933 ;
    wire new_AGEMA_signal_22934 ;
    wire new_AGEMA_signal_22935 ;
    wire new_AGEMA_signal_22936 ;
    wire new_AGEMA_signal_22937 ;
    wire new_AGEMA_signal_22938 ;
    wire new_AGEMA_signal_22939 ;
    wire new_AGEMA_signal_22940 ;
    wire new_AGEMA_signal_22941 ;
    wire new_AGEMA_signal_22942 ;
    wire new_AGEMA_signal_22943 ;
    wire new_AGEMA_signal_22944 ;
    wire new_AGEMA_signal_22945 ;
    wire new_AGEMA_signal_22946 ;
    wire new_AGEMA_signal_22947 ;
    wire new_AGEMA_signal_22948 ;
    wire new_AGEMA_signal_22949 ;
    wire new_AGEMA_signal_22950 ;
    wire new_AGEMA_signal_22951 ;
    wire new_AGEMA_signal_22952 ;
    wire new_AGEMA_signal_22953 ;
    wire new_AGEMA_signal_22954 ;
    wire new_AGEMA_signal_22955 ;
    wire new_AGEMA_signal_22956 ;
    wire new_AGEMA_signal_22957 ;
    wire new_AGEMA_signal_22958 ;
    wire new_AGEMA_signal_22959 ;
    wire new_AGEMA_signal_22960 ;
    wire new_AGEMA_signal_22961 ;
    wire new_AGEMA_signal_22962 ;
    wire new_AGEMA_signal_22963 ;
    wire new_AGEMA_signal_22964 ;
    wire new_AGEMA_signal_22965 ;
    wire new_AGEMA_signal_22966 ;
    wire new_AGEMA_signal_22967 ;
    wire new_AGEMA_signal_22968 ;
    wire new_AGEMA_signal_22969 ;
    wire new_AGEMA_signal_22970 ;
    wire new_AGEMA_signal_22971 ;
    wire new_AGEMA_signal_22972 ;
    wire new_AGEMA_signal_22973 ;
    wire new_AGEMA_signal_22974 ;
    wire new_AGEMA_signal_22975 ;
    wire new_AGEMA_signal_22976 ;
    wire new_AGEMA_signal_22977 ;
    wire new_AGEMA_signal_22978 ;
    wire new_AGEMA_signal_22979 ;
    wire new_AGEMA_signal_22980 ;
    wire new_AGEMA_signal_22981 ;
    wire new_AGEMA_signal_22982 ;
    wire new_AGEMA_signal_22983 ;
    wire new_AGEMA_signal_22984 ;
    wire new_AGEMA_signal_22985 ;
    wire new_AGEMA_signal_22986 ;
    wire new_AGEMA_signal_22987 ;
    wire new_AGEMA_signal_22988 ;
    wire new_AGEMA_signal_22989 ;
    wire new_AGEMA_signal_22990 ;
    wire new_AGEMA_signal_22991 ;
    wire new_AGEMA_signal_22992 ;
    wire new_AGEMA_signal_22993 ;
    wire new_AGEMA_signal_22994 ;
    wire new_AGEMA_signal_22995 ;
    wire new_AGEMA_signal_22996 ;
    wire new_AGEMA_signal_22997 ;
    wire new_AGEMA_signal_22998 ;
    wire new_AGEMA_signal_22999 ;
    wire new_AGEMA_signal_23000 ;
    wire new_AGEMA_signal_23001 ;
    wire new_AGEMA_signal_23002 ;
    wire new_AGEMA_signal_23003 ;
    wire new_AGEMA_signal_23004 ;
    wire new_AGEMA_signal_23005 ;
    wire new_AGEMA_signal_23006 ;
    wire new_AGEMA_signal_23007 ;
    wire new_AGEMA_signal_23008 ;
    wire new_AGEMA_signal_23009 ;
    wire new_AGEMA_signal_23010 ;
    wire new_AGEMA_signal_23011 ;
    wire new_AGEMA_signal_23012 ;
    wire new_AGEMA_signal_23013 ;
    wire new_AGEMA_signal_23014 ;
    wire new_AGEMA_signal_23015 ;
    wire new_AGEMA_signal_23016 ;
    wire new_AGEMA_signal_23017 ;
    wire new_AGEMA_signal_23018 ;
    wire new_AGEMA_signal_23019 ;
    wire new_AGEMA_signal_23020 ;
    wire new_AGEMA_signal_23021 ;
    wire new_AGEMA_signal_23022 ;
    wire new_AGEMA_signal_23023 ;
    wire new_AGEMA_signal_23024 ;
    wire new_AGEMA_signal_23025 ;
    wire new_AGEMA_signal_23026 ;
    wire new_AGEMA_signal_23027 ;
    wire new_AGEMA_signal_23028 ;
    wire new_AGEMA_signal_23029 ;
    wire new_AGEMA_signal_23030 ;
    wire new_AGEMA_signal_23031 ;
    wire new_AGEMA_signal_23032 ;
    wire new_AGEMA_signal_23033 ;
    wire new_AGEMA_signal_23034 ;
    wire new_AGEMA_signal_23035 ;
    wire new_AGEMA_signal_23036 ;
    wire new_AGEMA_signal_23037 ;
    wire new_AGEMA_signal_23038 ;
    wire new_AGEMA_signal_23039 ;
    wire new_AGEMA_signal_23040 ;
    wire new_AGEMA_signal_23041 ;
    wire new_AGEMA_signal_23042 ;
    wire new_AGEMA_signal_23043 ;
    wire new_AGEMA_signal_23044 ;
    wire new_AGEMA_signal_23045 ;
    wire new_AGEMA_signal_23046 ;
    wire new_AGEMA_signal_23047 ;
    wire new_AGEMA_signal_23048 ;
    wire new_AGEMA_signal_23049 ;
    wire new_AGEMA_signal_23050 ;
    wire new_AGEMA_signal_23051 ;
    wire new_AGEMA_signal_23052 ;
    wire new_AGEMA_signal_23053 ;
    wire new_AGEMA_signal_23054 ;
    wire new_AGEMA_signal_23055 ;
    wire new_AGEMA_signal_23056 ;
    wire new_AGEMA_signal_23057 ;
    wire new_AGEMA_signal_23058 ;
    wire new_AGEMA_signal_23059 ;
    wire new_AGEMA_signal_23060 ;
    wire new_AGEMA_signal_23061 ;
    wire new_AGEMA_signal_23062 ;
    wire new_AGEMA_signal_23063 ;
    wire new_AGEMA_signal_23064 ;
    wire new_AGEMA_signal_23065 ;
    wire new_AGEMA_signal_23066 ;
    wire new_AGEMA_signal_23067 ;
    wire new_AGEMA_signal_23068 ;
    wire new_AGEMA_signal_23069 ;
    wire new_AGEMA_signal_23070 ;
    wire new_AGEMA_signal_23071 ;
    wire new_AGEMA_signal_23072 ;
    wire new_AGEMA_signal_23073 ;
    wire new_AGEMA_signal_23074 ;
    wire new_AGEMA_signal_23075 ;
    wire new_AGEMA_signal_23076 ;
    wire new_AGEMA_signal_23077 ;
    wire new_AGEMA_signal_23078 ;
    wire new_AGEMA_signal_23079 ;
    wire new_AGEMA_signal_23080 ;
    wire new_AGEMA_signal_23081 ;
    wire new_AGEMA_signal_23082 ;
    wire new_AGEMA_signal_23083 ;
    wire new_AGEMA_signal_23084 ;
    wire new_AGEMA_signal_23085 ;
    wire new_AGEMA_signal_23086 ;
    wire new_AGEMA_signal_23087 ;
    wire new_AGEMA_signal_23088 ;
    wire new_AGEMA_signal_23089 ;
    wire new_AGEMA_signal_23090 ;
    wire new_AGEMA_signal_23091 ;
    wire new_AGEMA_signal_23092 ;
    wire new_AGEMA_signal_23093 ;
    wire new_AGEMA_signal_23094 ;
    wire new_AGEMA_signal_23095 ;
    wire new_AGEMA_signal_23096 ;
    wire new_AGEMA_signal_23097 ;
    wire new_AGEMA_signal_23098 ;
    wire new_AGEMA_signal_23099 ;
    wire new_AGEMA_signal_23100 ;
    wire new_AGEMA_signal_23101 ;
    wire new_AGEMA_signal_23102 ;
    wire new_AGEMA_signal_23103 ;
    wire new_AGEMA_signal_23104 ;
    wire new_AGEMA_signal_23105 ;
    wire new_AGEMA_signal_23106 ;
    wire new_AGEMA_signal_23107 ;
    wire new_AGEMA_signal_23108 ;
    wire new_AGEMA_signal_23109 ;
    wire new_AGEMA_signal_23110 ;
    wire new_AGEMA_signal_23111 ;
    wire new_AGEMA_signal_23112 ;
    wire new_AGEMA_signal_23113 ;
    wire new_AGEMA_signal_23114 ;
    wire new_AGEMA_signal_23115 ;
    wire new_AGEMA_signal_23116 ;
    wire new_AGEMA_signal_23117 ;
    wire new_AGEMA_signal_23118 ;
    wire new_AGEMA_signal_23119 ;
    wire new_AGEMA_signal_23120 ;
    wire new_AGEMA_signal_23121 ;
    wire new_AGEMA_signal_23122 ;
    wire new_AGEMA_signal_23123 ;
    wire new_AGEMA_signal_23124 ;
    wire new_AGEMA_signal_23125 ;
    wire new_AGEMA_signal_23126 ;
    wire new_AGEMA_signal_23127 ;
    wire new_AGEMA_signal_23128 ;
    wire new_AGEMA_signal_23129 ;
    wire new_AGEMA_signal_23130 ;
    wire new_AGEMA_signal_23131 ;
    wire new_AGEMA_signal_23132 ;
    wire new_AGEMA_signal_23133 ;
    wire new_AGEMA_signal_23134 ;
    wire new_AGEMA_signal_23135 ;
    wire new_AGEMA_signal_23136 ;
    wire new_AGEMA_signal_23137 ;
    wire new_AGEMA_signal_23138 ;
    wire new_AGEMA_signal_23139 ;
    wire new_AGEMA_signal_23140 ;
    wire new_AGEMA_signal_23141 ;
    wire new_AGEMA_signal_23142 ;
    wire new_AGEMA_signal_23143 ;
    wire new_AGEMA_signal_23144 ;
    wire new_AGEMA_signal_23145 ;
    wire new_AGEMA_signal_23146 ;
    wire new_AGEMA_signal_23147 ;
    wire new_AGEMA_signal_23148 ;
    wire new_AGEMA_signal_23149 ;
    wire new_AGEMA_signal_23150 ;
    wire new_AGEMA_signal_23151 ;
    wire new_AGEMA_signal_23152 ;
    wire new_AGEMA_signal_23153 ;
    wire new_AGEMA_signal_23154 ;
    wire new_AGEMA_signal_23155 ;
    wire new_AGEMA_signal_23156 ;
    wire new_AGEMA_signal_23157 ;
    wire new_AGEMA_signal_23158 ;
    wire new_AGEMA_signal_23159 ;
    wire new_AGEMA_signal_23160 ;
    wire new_AGEMA_signal_23161 ;
    wire new_AGEMA_signal_23162 ;
    wire new_AGEMA_signal_23163 ;
    wire new_AGEMA_signal_23164 ;
    wire new_AGEMA_signal_23165 ;
    wire new_AGEMA_signal_23166 ;
    wire new_AGEMA_signal_23167 ;
    wire new_AGEMA_signal_23168 ;
    wire new_AGEMA_signal_23169 ;
    wire new_AGEMA_signal_23170 ;
    wire new_AGEMA_signal_23171 ;
    wire new_AGEMA_signal_23172 ;
    wire new_AGEMA_signal_23173 ;
    wire new_AGEMA_signal_23174 ;
    wire new_AGEMA_signal_23175 ;
    wire new_AGEMA_signal_23176 ;
    wire new_AGEMA_signal_23177 ;
    wire new_AGEMA_signal_23178 ;
    wire new_AGEMA_signal_23179 ;
    wire new_AGEMA_signal_23180 ;
    wire new_AGEMA_signal_23181 ;
    wire new_AGEMA_signal_23182 ;
    wire new_AGEMA_signal_23183 ;
    wire new_AGEMA_signal_23184 ;
    wire new_AGEMA_signal_23185 ;
    wire new_AGEMA_signal_23186 ;
    wire new_AGEMA_signal_23187 ;
    wire new_AGEMA_signal_23188 ;
    wire new_AGEMA_signal_23189 ;
    wire new_AGEMA_signal_23190 ;
    wire new_AGEMA_signal_23191 ;
    wire new_AGEMA_signal_23192 ;
    wire new_AGEMA_signal_23193 ;
    wire new_AGEMA_signal_23194 ;
    wire new_AGEMA_signal_23195 ;
    wire new_AGEMA_signal_23196 ;
    wire new_AGEMA_signal_23197 ;
    wire new_AGEMA_signal_23198 ;
    wire new_AGEMA_signal_23199 ;
    wire new_AGEMA_signal_23200 ;
    wire new_AGEMA_signal_23201 ;
    wire new_AGEMA_signal_23202 ;
    wire new_AGEMA_signal_23203 ;
    wire new_AGEMA_signal_23204 ;
    wire new_AGEMA_signal_23205 ;
    wire new_AGEMA_signal_23206 ;
    wire new_AGEMA_signal_23207 ;
    wire new_AGEMA_signal_23208 ;
    wire new_AGEMA_signal_23209 ;
    wire new_AGEMA_signal_23210 ;
    wire new_AGEMA_signal_23211 ;
    wire new_AGEMA_signal_23212 ;
    wire new_AGEMA_signal_23213 ;
    wire new_AGEMA_signal_23214 ;
    wire new_AGEMA_signal_23215 ;
    wire new_AGEMA_signal_23216 ;
    wire new_AGEMA_signal_23217 ;
    wire new_AGEMA_signal_23218 ;
    wire new_AGEMA_signal_23219 ;
    wire new_AGEMA_signal_23220 ;
    wire new_AGEMA_signal_23221 ;
    wire new_AGEMA_signal_23222 ;
    wire new_AGEMA_signal_23223 ;
    wire new_AGEMA_signal_23224 ;
    wire new_AGEMA_signal_23225 ;
    wire new_AGEMA_signal_23226 ;
    wire new_AGEMA_signal_23227 ;
    wire new_AGEMA_signal_23228 ;
    wire new_AGEMA_signal_23229 ;
    wire new_AGEMA_signal_23230 ;
    wire new_AGEMA_signal_23231 ;
    wire new_AGEMA_signal_23232 ;
    wire new_AGEMA_signal_23233 ;
    wire new_AGEMA_signal_23234 ;
    wire new_AGEMA_signal_23235 ;
    wire new_AGEMA_signal_23236 ;
    wire new_AGEMA_signal_23237 ;
    wire new_AGEMA_signal_23238 ;
    wire new_AGEMA_signal_23239 ;
    wire new_AGEMA_signal_23240 ;
    wire new_AGEMA_signal_23241 ;
    wire new_AGEMA_signal_23242 ;
    wire new_AGEMA_signal_23243 ;
    wire new_AGEMA_signal_23244 ;
    wire new_AGEMA_signal_23245 ;
    wire new_AGEMA_signal_23246 ;
    wire new_AGEMA_signal_23247 ;
    wire new_AGEMA_signal_23248 ;
    wire new_AGEMA_signal_23249 ;
    wire new_AGEMA_signal_23250 ;
    wire new_AGEMA_signal_23251 ;
    wire new_AGEMA_signal_23252 ;
    wire new_AGEMA_signal_23253 ;
    wire new_AGEMA_signal_23254 ;
    wire new_AGEMA_signal_23255 ;
    wire new_AGEMA_signal_23256 ;
    wire new_AGEMA_signal_23257 ;
    wire new_AGEMA_signal_23258 ;
    wire new_AGEMA_signal_23259 ;
    wire new_AGEMA_signal_23260 ;
    wire new_AGEMA_signal_23261 ;
    wire new_AGEMA_signal_23262 ;
    wire new_AGEMA_signal_23263 ;
    wire new_AGEMA_signal_23264 ;
    wire new_AGEMA_signal_23265 ;
    wire new_AGEMA_signal_23266 ;
    wire new_AGEMA_signal_23267 ;
    wire new_AGEMA_signal_23268 ;
    wire new_AGEMA_signal_23269 ;
    wire new_AGEMA_signal_23270 ;
    wire new_AGEMA_signal_23271 ;
    wire new_AGEMA_signal_23272 ;
    wire new_AGEMA_signal_23273 ;
    wire new_AGEMA_signal_23274 ;
    wire new_AGEMA_signal_23275 ;
    wire new_AGEMA_signal_23276 ;
    wire new_AGEMA_signal_23277 ;
    wire new_AGEMA_signal_23278 ;
    wire new_AGEMA_signal_23279 ;
    wire new_AGEMA_signal_23280 ;
    wire new_AGEMA_signal_23281 ;
    wire new_AGEMA_signal_23282 ;
    wire new_AGEMA_signal_23283 ;
    wire new_AGEMA_signal_23284 ;
    wire new_AGEMA_signal_23285 ;
    wire new_AGEMA_signal_23286 ;
    wire new_AGEMA_signal_23287 ;
    wire new_AGEMA_signal_23288 ;
    wire new_AGEMA_signal_23289 ;
    wire new_AGEMA_signal_23290 ;
    wire new_AGEMA_signal_23291 ;
    wire new_AGEMA_signal_23292 ;
    wire new_AGEMA_signal_23293 ;
    wire new_AGEMA_signal_23294 ;
    wire new_AGEMA_signal_23295 ;
    wire new_AGEMA_signal_23296 ;
    wire new_AGEMA_signal_23297 ;
    wire new_AGEMA_signal_23298 ;
    wire new_AGEMA_signal_23299 ;
    wire new_AGEMA_signal_23300 ;
    wire new_AGEMA_signal_23301 ;
    wire new_AGEMA_signal_23302 ;
    wire new_AGEMA_signal_23303 ;
    wire new_AGEMA_signal_23304 ;
    wire new_AGEMA_signal_23305 ;
    wire new_AGEMA_signal_23306 ;
    wire new_AGEMA_signal_23307 ;
    wire new_AGEMA_signal_23308 ;
    wire new_AGEMA_signal_23309 ;
    wire new_AGEMA_signal_23310 ;
    wire new_AGEMA_signal_23311 ;
    wire new_AGEMA_signal_23312 ;
    wire new_AGEMA_signal_23313 ;
    wire new_AGEMA_signal_23314 ;
    wire new_AGEMA_signal_23315 ;
    wire new_AGEMA_signal_23316 ;
    wire new_AGEMA_signal_23317 ;
    wire new_AGEMA_signal_23318 ;
    wire new_AGEMA_signal_23319 ;
    wire new_AGEMA_signal_23320 ;
    wire new_AGEMA_signal_23321 ;
    wire new_AGEMA_signal_23322 ;
    wire new_AGEMA_signal_23323 ;
    wire new_AGEMA_signal_23324 ;
    wire new_AGEMA_signal_23325 ;
    wire new_AGEMA_signal_23326 ;
    wire new_AGEMA_signal_23327 ;
    wire new_AGEMA_signal_23328 ;
    wire new_AGEMA_signal_23329 ;
    wire new_AGEMA_signal_23330 ;
    wire new_AGEMA_signal_23331 ;
    wire new_AGEMA_signal_23332 ;
    wire new_AGEMA_signal_23333 ;
    wire new_AGEMA_signal_23334 ;
    wire new_AGEMA_signal_23335 ;
    wire new_AGEMA_signal_23336 ;
    wire new_AGEMA_signal_23337 ;
    wire new_AGEMA_signal_23338 ;
    wire new_AGEMA_signal_23339 ;
    wire new_AGEMA_signal_23340 ;
    wire new_AGEMA_signal_23341 ;
    wire new_AGEMA_signal_23342 ;
    wire new_AGEMA_signal_23343 ;
    wire new_AGEMA_signal_23344 ;
    wire new_AGEMA_signal_23345 ;
    wire new_AGEMA_signal_23346 ;
    wire new_AGEMA_signal_23347 ;
    wire new_AGEMA_signal_23348 ;
    wire new_AGEMA_signal_23349 ;
    wire new_AGEMA_signal_23350 ;
    wire new_AGEMA_signal_23351 ;
    wire new_AGEMA_signal_23352 ;
    wire new_AGEMA_signal_23353 ;
    wire new_AGEMA_signal_23354 ;
    wire new_AGEMA_signal_23355 ;
    wire new_AGEMA_signal_23356 ;
    wire new_AGEMA_signal_23357 ;
    wire new_AGEMA_signal_23358 ;
    wire new_AGEMA_signal_23359 ;
    wire new_AGEMA_signal_23360 ;
    wire new_AGEMA_signal_23361 ;
    wire new_AGEMA_signal_23362 ;
    wire new_AGEMA_signal_23363 ;
    wire new_AGEMA_signal_23364 ;
    wire new_AGEMA_signal_23365 ;
    wire new_AGEMA_signal_23366 ;
    wire new_AGEMA_signal_23367 ;
    wire new_AGEMA_signal_23368 ;
    wire new_AGEMA_signal_23369 ;
    wire new_AGEMA_signal_23370 ;
    wire new_AGEMA_signal_23371 ;
    wire new_AGEMA_signal_23372 ;
    wire new_AGEMA_signal_23373 ;
    wire new_AGEMA_signal_23374 ;
    wire new_AGEMA_signal_23375 ;
    wire new_AGEMA_signal_23376 ;
    wire new_AGEMA_signal_23377 ;
    wire new_AGEMA_signal_23378 ;
    wire new_AGEMA_signal_23379 ;
    wire new_AGEMA_signal_23380 ;
    wire new_AGEMA_signal_23381 ;
    wire new_AGEMA_signal_23382 ;
    wire new_AGEMA_signal_23383 ;
    wire new_AGEMA_signal_23384 ;
    wire new_AGEMA_signal_23385 ;
    wire new_AGEMA_signal_23386 ;
    wire new_AGEMA_signal_23387 ;
    wire new_AGEMA_signal_23388 ;
    wire new_AGEMA_signal_23389 ;
    wire new_AGEMA_signal_23390 ;
    wire new_AGEMA_signal_23391 ;
    wire new_AGEMA_signal_23392 ;
    wire new_AGEMA_signal_23393 ;
    wire new_AGEMA_signal_23394 ;
    wire new_AGEMA_signal_23395 ;
    wire new_AGEMA_signal_23396 ;
    wire new_AGEMA_signal_23397 ;
    wire new_AGEMA_signal_23398 ;
    wire new_AGEMA_signal_23399 ;
    wire new_AGEMA_signal_23400 ;
    wire new_AGEMA_signal_23401 ;
    wire new_AGEMA_signal_23402 ;
    wire new_AGEMA_signal_23403 ;
    wire new_AGEMA_signal_23404 ;
    wire new_AGEMA_signal_23405 ;
    wire new_AGEMA_signal_23406 ;
    wire new_AGEMA_signal_23407 ;
    wire new_AGEMA_signal_23408 ;
    wire new_AGEMA_signal_23409 ;
    wire new_AGEMA_signal_23410 ;
    wire new_AGEMA_signal_23411 ;
    wire new_AGEMA_signal_23412 ;
    wire new_AGEMA_signal_23413 ;
    wire new_AGEMA_signal_23414 ;
    wire new_AGEMA_signal_23415 ;
    wire new_AGEMA_signal_23416 ;
    wire new_AGEMA_signal_23417 ;
    wire new_AGEMA_signal_23418 ;
    wire new_AGEMA_signal_23419 ;
    wire new_AGEMA_signal_23420 ;
    wire new_AGEMA_signal_23421 ;
    wire new_AGEMA_signal_23422 ;
    wire new_AGEMA_signal_23423 ;
    wire new_AGEMA_signal_23424 ;
    wire new_AGEMA_signal_23425 ;
    wire new_AGEMA_signal_23426 ;
    wire new_AGEMA_signal_23427 ;
    wire new_AGEMA_signal_23428 ;
    wire new_AGEMA_signal_23429 ;
    wire new_AGEMA_signal_23430 ;
    wire new_AGEMA_signal_23431 ;
    wire new_AGEMA_signal_23432 ;
    wire new_AGEMA_signal_23433 ;
    wire new_AGEMA_signal_23434 ;
    wire new_AGEMA_signal_23435 ;
    wire new_AGEMA_signal_23436 ;
    wire new_AGEMA_signal_23437 ;
    wire new_AGEMA_signal_23438 ;
    wire new_AGEMA_signal_23439 ;
    wire new_AGEMA_signal_23440 ;
    wire new_AGEMA_signal_23441 ;
    wire new_AGEMA_signal_23442 ;
    wire new_AGEMA_signal_23443 ;
    wire new_AGEMA_signal_23444 ;
    wire new_AGEMA_signal_23445 ;
    wire new_AGEMA_signal_23446 ;
    wire new_AGEMA_signal_23447 ;
    wire new_AGEMA_signal_23448 ;
    wire new_AGEMA_signal_23449 ;
    wire new_AGEMA_signal_23450 ;
    wire new_AGEMA_signal_23451 ;
    wire new_AGEMA_signal_23452 ;
    wire new_AGEMA_signal_23453 ;
    wire new_AGEMA_signal_23454 ;
    wire new_AGEMA_signal_23455 ;
    wire new_AGEMA_signal_23456 ;
    wire new_AGEMA_signal_23457 ;
    wire new_AGEMA_signal_23458 ;
    wire new_AGEMA_signal_23459 ;
    wire new_AGEMA_signal_23460 ;
    wire new_AGEMA_signal_23461 ;
    wire new_AGEMA_signal_23462 ;
    wire new_AGEMA_signal_23463 ;
    wire new_AGEMA_signal_23464 ;
    wire new_AGEMA_signal_23465 ;
    wire new_AGEMA_signal_23466 ;
    wire new_AGEMA_signal_23467 ;
    wire new_AGEMA_signal_23468 ;
    wire new_AGEMA_signal_23469 ;
    wire new_AGEMA_signal_23470 ;
    wire new_AGEMA_signal_23471 ;
    wire new_AGEMA_signal_23472 ;
    wire new_AGEMA_signal_23473 ;
    wire new_AGEMA_signal_23474 ;
    wire new_AGEMA_signal_23475 ;
    wire new_AGEMA_signal_23476 ;
    wire new_AGEMA_signal_23477 ;
    wire new_AGEMA_signal_23478 ;
    wire new_AGEMA_signal_23479 ;
    wire new_AGEMA_signal_23480 ;
    wire new_AGEMA_signal_23481 ;
    wire new_AGEMA_signal_23482 ;
    wire new_AGEMA_signal_23483 ;
    wire new_AGEMA_signal_23484 ;
    wire new_AGEMA_signal_23485 ;
    wire new_AGEMA_signal_23486 ;
    wire new_AGEMA_signal_23487 ;
    wire new_AGEMA_signal_23488 ;
    wire new_AGEMA_signal_23489 ;
    wire new_AGEMA_signal_23490 ;
    wire new_AGEMA_signal_23491 ;
    wire new_AGEMA_signal_23492 ;
    wire new_AGEMA_signal_23493 ;
    wire new_AGEMA_signal_23494 ;
    wire new_AGEMA_signal_23495 ;
    wire new_AGEMA_signal_23496 ;
    wire new_AGEMA_signal_23497 ;
    wire new_AGEMA_signal_23498 ;
    wire new_AGEMA_signal_23499 ;
    wire new_AGEMA_signal_23500 ;
    wire new_AGEMA_signal_23501 ;
    wire new_AGEMA_signal_23502 ;
    wire new_AGEMA_signal_23503 ;
    wire new_AGEMA_signal_23504 ;
    wire new_AGEMA_signal_23505 ;
    wire new_AGEMA_signal_23506 ;
    wire new_AGEMA_signal_23507 ;
    wire new_AGEMA_signal_23508 ;
    wire new_AGEMA_signal_23509 ;
    wire new_AGEMA_signal_23510 ;
    wire new_AGEMA_signal_23511 ;
    wire new_AGEMA_signal_23512 ;
    wire new_AGEMA_signal_23513 ;
    wire new_AGEMA_signal_23514 ;
    wire new_AGEMA_signal_23515 ;
    wire new_AGEMA_signal_23516 ;
    wire new_AGEMA_signal_23517 ;
    wire new_AGEMA_signal_23518 ;
    wire new_AGEMA_signal_23519 ;
    wire new_AGEMA_signal_23520 ;
    wire new_AGEMA_signal_23521 ;
    wire new_AGEMA_signal_23522 ;
    wire new_AGEMA_signal_23523 ;
    wire new_AGEMA_signal_23524 ;
    wire new_AGEMA_signal_23525 ;
    wire new_AGEMA_signal_23526 ;
    wire new_AGEMA_signal_23527 ;
    wire new_AGEMA_signal_23528 ;
    wire new_AGEMA_signal_23529 ;
    wire new_AGEMA_signal_23530 ;
    wire new_AGEMA_signal_23531 ;
    wire new_AGEMA_signal_23532 ;
    wire new_AGEMA_signal_23533 ;
    wire new_AGEMA_signal_23534 ;
    wire new_AGEMA_signal_23535 ;
    wire new_AGEMA_signal_23536 ;
    wire new_AGEMA_signal_23537 ;
    wire new_AGEMA_signal_23538 ;
    wire new_AGEMA_signal_23539 ;
    wire new_AGEMA_signal_23540 ;
    wire new_AGEMA_signal_23541 ;
    wire new_AGEMA_signal_23542 ;
    wire new_AGEMA_signal_23543 ;
    wire new_AGEMA_signal_23544 ;
    wire new_AGEMA_signal_23545 ;
    wire new_AGEMA_signal_23546 ;
    wire new_AGEMA_signal_23547 ;
    wire new_AGEMA_signal_23548 ;
    wire new_AGEMA_signal_23549 ;
    wire new_AGEMA_signal_23550 ;
    wire new_AGEMA_signal_23551 ;
    wire new_AGEMA_signal_23552 ;
    wire new_AGEMA_signal_23553 ;
    wire new_AGEMA_signal_23554 ;
    wire new_AGEMA_signal_23555 ;
    wire new_AGEMA_signal_23556 ;
    wire new_AGEMA_signal_23557 ;
    wire new_AGEMA_signal_23558 ;
    wire new_AGEMA_signal_23559 ;
    wire new_AGEMA_signal_23560 ;
    wire new_AGEMA_signal_23561 ;
    wire new_AGEMA_signal_23562 ;
    wire new_AGEMA_signal_23563 ;
    wire new_AGEMA_signal_23564 ;
    wire new_AGEMA_signal_23565 ;
    wire new_AGEMA_signal_23566 ;
    wire new_AGEMA_signal_23567 ;
    wire new_AGEMA_signal_23568 ;
    wire new_AGEMA_signal_23569 ;
    wire new_AGEMA_signal_23570 ;
    wire new_AGEMA_signal_23571 ;
    wire new_AGEMA_signal_23572 ;
    wire new_AGEMA_signal_23573 ;
    wire new_AGEMA_signal_23574 ;
    wire new_AGEMA_signal_23575 ;
    wire new_AGEMA_signal_23576 ;
    wire new_AGEMA_signal_23577 ;
    wire new_AGEMA_signal_23578 ;
    wire new_AGEMA_signal_23579 ;
    wire new_AGEMA_signal_23580 ;
    wire new_AGEMA_signal_23581 ;
    wire new_AGEMA_signal_23582 ;
    wire new_AGEMA_signal_23583 ;
    wire new_AGEMA_signal_23584 ;
    wire new_AGEMA_signal_23585 ;
    wire new_AGEMA_signal_23586 ;
    wire new_AGEMA_signal_23587 ;
    wire new_AGEMA_signal_23588 ;
    wire new_AGEMA_signal_23589 ;
    wire new_AGEMA_signal_23590 ;
    wire new_AGEMA_signal_23591 ;
    wire new_AGEMA_signal_23592 ;
    wire new_AGEMA_signal_23593 ;
    wire new_AGEMA_signal_23594 ;
    wire new_AGEMA_signal_23595 ;
    wire new_AGEMA_signal_23596 ;
    wire new_AGEMA_signal_23597 ;
    wire new_AGEMA_signal_23598 ;
    wire new_AGEMA_signal_23599 ;
    wire new_AGEMA_signal_23600 ;
    wire new_AGEMA_signal_23601 ;
    wire new_AGEMA_signal_23602 ;
    wire new_AGEMA_signal_23603 ;
    wire new_AGEMA_signal_23604 ;
    wire new_AGEMA_signal_23605 ;
    wire new_AGEMA_signal_23606 ;
    wire new_AGEMA_signal_23607 ;
    wire new_AGEMA_signal_23608 ;
    wire new_AGEMA_signal_23609 ;
    wire new_AGEMA_signal_23610 ;
    wire new_AGEMA_signal_23611 ;
    wire new_AGEMA_signal_23612 ;
    wire new_AGEMA_signal_23613 ;
    wire new_AGEMA_signal_23614 ;
    wire new_AGEMA_signal_23615 ;
    wire new_AGEMA_signal_23616 ;
    wire new_AGEMA_signal_23617 ;
    wire new_AGEMA_signal_23618 ;
    wire new_AGEMA_signal_23619 ;
    wire new_AGEMA_signal_23620 ;
    wire new_AGEMA_signal_23621 ;
    wire new_AGEMA_signal_23622 ;
    wire new_AGEMA_signal_23623 ;
    wire new_AGEMA_signal_23624 ;
    wire new_AGEMA_signal_23625 ;
    wire new_AGEMA_signal_23626 ;
    wire new_AGEMA_signal_23627 ;
    wire new_AGEMA_signal_23628 ;
    wire new_AGEMA_signal_23629 ;
    wire new_AGEMA_signal_23630 ;
    wire new_AGEMA_signal_23631 ;
    wire new_AGEMA_signal_23632 ;
    wire new_AGEMA_signal_23633 ;
    wire new_AGEMA_signal_23634 ;
    wire new_AGEMA_signal_23635 ;
    wire new_AGEMA_signal_23636 ;
    wire new_AGEMA_signal_23637 ;
    wire new_AGEMA_signal_23638 ;
    wire new_AGEMA_signal_23639 ;
    wire new_AGEMA_signal_23640 ;
    wire new_AGEMA_signal_23641 ;
    wire new_AGEMA_signal_23642 ;
    wire new_AGEMA_signal_23643 ;
    wire new_AGEMA_signal_23644 ;
    wire new_AGEMA_signal_23645 ;
    wire new_AGEMA_signal_23646 ;
    wire new_AGEMA_signal_23647 ;
    wire new_AGEMA_signal_23648 ;
    wire new_AGEMA_signal_23649 ;
    wire new_AGEMA_signal_23650 ;
    wire new_AGEMA_signal_23651 ;
    wire new_AGEMA_signal_23652 ;
    wire new_AGEMA_signal_23653 ;
    wire new_AGEMA_signal_23654 ;
    wire new_AGEMA_signal_23655 ;
    wire new_AGEMA_signal_23656 ;
    wire new_AGEMA_signal_23657 ;
    wire new_AGEMA_signal_23658 ;
    wire new_AGEMA_signal_23659 ;
    wire new_AGEMA_signal_23660 ;
    wire new_AGEMA_signal_23661 ;
    wire new_AGEMA_signal_23662 ;
    wire new_AGEMA_signal_23663 ;
    wire new_AGEMA_signal_23664 ;
    wire new_AGEMA_signal_23665 ;
    wire new_AGEMA_signal_23666 ;
    wire new_AGEMA_signal_23667 ;
    wire new_AGEMA_signal_23668 ;
    wire new_AGEMA_signal_23669 ;
    wire new_AGEMA_signal_23670 ;
    wire new_AGEMA_signal_23671 ;
    wire new_AGEMA_signal_23672 ;
    wire new_AGEMA_signal_23673 ;
    wire new_AGEMA_signal_23674 ;
    wire new_AGEMA_signal_23675 ;
    wire new_AGEMA_signal_23676 ;
    wire new_AGEMA_signal_23677 ;
    wire new_AGEMA_signal_23678 ;
    wire new_AGEMA_signal_23679 ;
    wire new_AGEMA_signal_23680 ;
    wire new_AGEMA_signal_23681 ;
    wire new_AGEMA_signal_23682 ;
    wire new_AGEMA_signal_23683 ;
    wire new_AGEMA_signal_23684 ;
    wire new_AGEMA_signal_23685 ;
    wire new_AGEMA_signal_23686 ;
    wire new_AGEMA_signal_23687 ;
    wire new_AGEMA_signal_23688 ;
    wire new_AGEMA_signal_23689 ;
    wire new_AGEMA_signal_23690 ;
    wire new_AGEMA_signal_23691 ;
    wire new_AGEMA_signal_23692 ;
    wire new_AGEMA_signal_23693 ;
    wire new_AGEMA_signal_23694 ;
    wire new_AGEMA_signal_23695 ;
    wire new_AGEMA_signal_23696 ;
    wire new_AGEMA_signal_23697 ;
    wire new_AGEMA_signal_23698 ;
    wire new_AGEMA_signal_23699 ;
    wire new_AGEMA_signal_23700 ;
    wire new_AGEMA_signal_23701 ;
    wire new_AGEMA_signal_23702 ;
    wire new_AGEMA_signal_23703 ;
    wire new_AGEMA_signal_23704 ;
    wire new_AGEMA_signal_23705 ;
    wire new_AGEMA_signal_23706 ;
    wire new_AGEMA_signal_23707 ;
    wire new_AGEMA_signal_23708 ;
    wire new_AGEMA_signal_23709 ;
    wire new_AGEMA_signal_23710 ;
    wire new_AGEMA_signal_23711 ;
    wire new_AGEMA_signal_23712 ;
    wire new_AGEMA_signal_23713 ;
    wire new_AGEMA_signal_23714 ;
    wire new_AGEMA_signal_23715 ;
    wire new_AGEMA_signal_23716 ;
    wire new_AGEMA_signal_23717 ;
    wire new_AGEMA_signal_23718 ;
    wire new_AGEMA_signal_23719 ;
    wire new_AGEMA_signal_23720 ;
    wire new_AGEMA_signal_23721 ;
    wire new_AGEMA_signal_23722 ;
    wire new_AGEMA_signal_23723 ;
    wire new_AGEMA_signal_23724 ;
    wire new_AGEMA_signal_23725 ;
    wire new_AGEMA_signal_23726 ;
    wire new_AGEMA_signal_23727 ;
    wire new_AGEMA_signal_23728 ;
    wire new_AGEMA_signal_23729 ;
    wire new_AGEMA_signal_23730 ;
    wire new_AGEMA_signal_23731 ;
    wire new_AGEMA_signal_23732 ;
    wire new_AGEMA_signal_23733 ;
    wire new_AGEMA_signal_23734 ;
    wire new_AGEMA_signal_23735 ;
    wire new_AGEMA_signal_23736 ;
    wire new_AGEMA_signal_23737 ;
    wire new_AGEMA_signal_23738 ;
    wire new_AGEMA_signal_23739 ;
    wire new_AGEMA_signal_23740 ;
    wire new_AGEMA_signal_23741 ;
    wire new_AGEMA_signal_23742 ;
    wire new_AGEMA_signal_23743 ;
    wire new_AGEMA_signal_23744 ;
    wire new_AGEMA_signal_23745 ;
    wire new_AGEMA_signal_23746 ;
    wire new_AGEMA_signal_23747 ;
    wire new_AGEMA_signal_23748 ;
    wire new_AGEMA_signal_23749 ;
    wire new_AGEMA_signal_23750 ;
    wire new_AGEMA_signal_23751 ;
    wire new_AGEMA_signal_23752 ;
    wire new_AGEMA_signal_23753 ;
    wire new_AGEMA_signal_23754 ;
    wire new_AGEMA_signal_23755 ;
    wire new_AGEMA_signal_23756 ;
    wire new_AGEMA_signal_23757 ;
    wire new_AGEMA_signal_23758 ;
    wire new_AGEMA_signal_23759 ;
    wire new_AGEMA_signal_23760 ;
    wire new_AGEMA_signal_23761 ;
    wire new_AGEMA_signal_23762 ;
    wire new_AGEMA_signal_23763 ;
    wire new_AGEMA_signal_23764 ;
    wire new_AGEMA_signal_23765 ;
    wire new_AGEMA_signal_23766 ;
    wire new_AGEMA_signal_23767 ;
    wire new_AGEMA_signal_23768 ;
    wire new_AGEMA_signal_23769 ;
    wire new_AGEMA_signal_23770 ;
    wire new_AGEMA_signal_23771 ;
    wire new_AGEMA_signal_23772 ;
    wire new_AGEMA_signal_23773 ;
    wire new_AGEMA_signal_23774 ;
    wire new_AGEMA_signal_23775 ;
    wire new_AGEMA_signal_23776 ;
    wire new_AGEMA_signal_23777 ;
    wire new_AGEMA_signal_23778 ;
    wire new_AGEMA_signal_23779 ;
    wire new_AGEMA_signal_23780 ;
    wire new_AGEMA_signal_23781 ;
    wire new_AGEMA_signal_23782 ;
    wire new_AGEMA_signal_23783 ;
    wire new_AGEMA_signal_23784 ;
    wire new_AGEMA_signal_23785 ;
    wire new_AGEMA_signal_23786 ;
    wire new_AGEMA_signal_23787 ;
    wire new_AGEMA_signal_23788 ;
    wire new_AGEMA_signal_23789 ;
    wire new_AGEMA_signal_23790 ;
    wire new_AGEMA_signal_23791 ;
    wire new_AGEMA_signal_23792 ;
    wire new_AGEMA_signal_23793 ;
    wire new_AGEMA_signal_23794 ;
    wire new_AGEMA_signal_23795 ;
    wire new_AGEMA_signal_23796 ;
    wire new_AGEMA_signal_23797 ;
    wire new_AGEMA_signal_23798 ;
    wire new_AGEMA_signal_23799 ;
    wire new_AGEMA_signal_23800 ;
    wire new_AGEMA_signal_23801 ;
    wire new_AGEMA_signal_23802 ;
    wire new_AGEMA_signal_23803 ;
    wire new_AGEMA_signal_23804 ;
    wire new_AGEMA_signal_23805 ;
    wire new_AGEMA_signal_23806 ;
    wire new_AGEMA_signal_23807 ;
    wire new_AGEMA_signal_23808 ;
    wire new_AGEMA_signal_23809 ;
    wire new_AGEMA_signal_23810 ;
    wire new_AGEMA_signal_23811 ;
    wire new_AGEMA_signal_23812 ;
    wire new_AGEMA_signal_23813 ;
    wire new_AGEMA_signal_23814 ;
    wire new_AGEMA_signal_23815 ;
    wire new_AGEMA_signal_23816 ;
    wire new_AGEMA_signal_23817 ;
    wire new_AGEMA_signal_23818 ;
    wire new_AGEMA_signal_23819 ;
    wire new_AGEMA_signal_23820 ;
    wire new_AGEMA_signal_23821 ;
    wire new_AGEMA_signal_23822 ;
    wire new_AGEMA_signal_23823 ;
    wire new_AGEMA_signal_23824 ;
    wire new_AGEMA_signal_23825 ;
    wire new_AGEMA_signal_23826 ;
    wire new_AGEMA_signal_23827 ;
    wire new_AGEMA_signal_23828 ;
    wire new_AGEMA_signal_23829 ;
    wire new_AGEMA_signal_23830 ;
    wire new_AGEMA_signal_23831 ;
    wire new_AGEMA_signal_23832 ;
    wire new_AGEMA_signal_23833 ;
    wire new_AGEMA_signal_23834 ;
    wire new_AGEMA_signal_23835 ;
    wire new_AGEMA_signal_23836 ;
    wire new_AGEMA_signal_23837 ;
    wire new_AGEMA_signal_23838 ;
    wire new_AGEMA_signal_23839 ;
    wire new_AGEMA_signal_23840 ;
    wire new_AGEMA_signal_23841 ;
    wire new_AGEMA_signal_23842 ;
    wire new_AGEMA_signal_23843 ;
    wire new_AGEMA_signal_23844 ;
    wire new_AGEMA_signal_23845 ;
    wire new_AGEMA_signal_23846 ;
    wire new_AGEMA_signal_23847 ;
    wire new_AGEMA_signal_23848 ;
    wire new_AGEMA_signal_23849 ;
    wire new_AGEMA_signal_23850 ;
    wire new_AGEMA_signal_23851 ;
    wire new_AGEMA_signal_23852 ;
    wire new_AGEMA_signal_23853 ;
    wire new_AGEMA_signal_23854 ;
    wire new_AGEMA_signal_23855 ;
    wire new_AGEMA_signal_23856 ;
    wire new_AGEMA_signal_23857 ;
    wire new_AGEMA_signal_23858 ;
    wire new_AGEMA_signal_23859 ;
    wire new_AGEMA_signal_23860 ;
    wire new_AGEMA_signal_23861 ;
    wire new_AGEMA_signal_23862 ;
    wire new_AGEMA_signal_23863 ;
    wire new_AGEMA_signal_23864 ;
    wire new_AGEMA_signal_23865 ;
    wire new_AGEMA_signal_23866 ;
    wire new_AGEMA_signal_23867 ;
    wire new_AGEMA_signal_23868 ;
    wire new_AGEMA_signal_23869 ;
    wire new_AGEMA_signal_23870 ;
    wire new_AGEMA_signal_23871 ;
    wire new_AGEMA_signal_23872 ;
    wire new_AGEMA_signal_23873 ;
    wire new_AGEMA_signal_23874 ;
    wire new_AGEMA_signal_23875 ;
    wire new_AGEMA_signal_23876 ;
    wire new_AGEMA_signal_23877 ;
    wire new_AGEMA_signal_23878 ;
    wire new_AGEMA_signal_23879 ;
    wire new_AGEMA_signal_23880 ;
    wire new_AGEMA_signal_23881 ;
    wire new_AGEMA_signal_23882 ;
    wire new_AGEMA_signal_23883 ;
    wire new_AGEMA_signal_23884 ;
    wire new_AGEMA_signal_23885 ;
    wire new_AGEMA_signal_23886 ;
    wire new_AGEMA_signal_23887 ;
    wire new_AGEMA_signal_23888 ;
    wire new_AGEMA_signal_23889 ;
    wire new_AGEMA_signal_23890 ;
    wire new_AGEMA_signal_23891 ;
    wire new_AGEMA_signal_23892 ;
    wire new_AGEMA_signal_23893 ;
    wire new_AGEMA_signal_23894 ;
    wire new_AGEMA_signal_23895 ;
    wire new_AGEMA_signal_23896 ;
    wire new_AGEMA_signal_23897 ;
    wire new_AGEMA_signal_23898 ;
    wire new_AGEMA_signal_23899 ;
    wire new_AGEMA_signal_23900 ;
    wire new_AGEMA_signal_23901 ;
    wire new_AGEMA_signal_23902 ;
    wire new_AGEMA_signal_23903 ;
    wire new_AGEMA_signal_23904 ;
    wire new_AGEMA_signal_23905 ;
    wire new_AGEMA_signal_23906 ;
    wire new_AGEMA_signal_23907 ;
    wire new_AGEMA_signal_23908 ;
    wire new_AGEMA_signal_23909 ;
    wire new_AGEMA_signal_23910 ;
    wire new_AGEMA_signal_23911 ;
    wire new_AGEMA_signal_23912 ;
    wire new_AGEMA_signal_23913 ;
    wire new_AGEMA_signal_23914 ;
    wire new_AGEMA_signal_23915 ;
    wire new_AGEMA_signal_23916 ;
    wire new_AGEMA_signal_23917 ;
    wire new_AGEMA_signal_23918 ;
    wire new_AGEMA_signal_23919 ;
    wire new_AGEMA_signal_23920 ;
    wire new_AGEMA_signal_23921 ;
    wire new_AGEMA_signal_23922 ;
    wire new_AGEMA_signal_23923 ;
    wire new_AGEMA_signal_23924 ;
    wire new_AGEMA_signal_23925 ;
    wire new_AGEMA_signal_23926 ;
    wire new_AGEMA_signal_23927 ;
    wire new_AGEMA_signal_23928 ;
    wire new_AGEMA_signal_23929 ;
    wire new_AGEMA_signal_23930 ;
    wire new_AGEMA_signal_23931 ;
    wire new_AGEMA_signal_23932 ;
    wire new_AGEMA_signal_23933 ;
    wire new_AGEMA_signal_23934 ;
    wire new_AGEMA_signal_23935 ;
    wire new_AGEMA_signal_23936 ;
    wire new_AGEMA_signal_23937 ;
    wire new_AGEMA_signal_23938 ;
    wire new_AGEMA_signal_23939 ;
    wire new_AGEMA_signal_23940 ;
    wire new_AGEMA_signal_23941 ;
    wire new_AGEMA_signal_23942 ;
    wire new_AGEMA_signal_23943 ;
    wire new_AGEMA_signal_23944 ;
    wire new_AGEMA_signal_23945 ;
    wire new_AGEMA_signal_23946 ;
    wire new_AGEMA_signal_23947 ;
    wire new_AGEMA_signal_23948 ;
    wire new_AGEMA_signal_23949 ;
    wire new_AGEMA_signal_23950 ;
    wire new_AGEMA_signal_23951 ;
    wire new_AGEMA_signal_23952 ;
    wire new_AGEMA_signal_23953 ;
    wire new_AGEMA_signal_23954 ;
    wire new_AGEMA_signal_23955 ;
    wire new_AGEMA_signal_23956 ;
    wire new_AGEMA_signal_23957 ;
    wire new_AGEMA_signal_23958 ;
    wire new_AGEMA_signal_23959 ;
    wire new_AGEMA_signal_23960 ;
    wire new_AGEMA_signal_23961 ;
    wire new_AGEMA_signal_23962 ;
    wire new_AGEMA_signal_23963 ;
    wire new_AGEMA_signal_23964 ;
    wire new_AGEMA_signal_23965 ;
    wire new_AGEMA_signal_23966 ;
    wire new_AGEMA_signal_23967 ;
    wire new_AGEMA_signal_23968 ;
    wire new_AGEMA_signal_23969 ;
    wire new_AGEMA_signal_23970 ;
    wire new_AGEMA_signal_23971 ;
    wire new_AGEMA_signal_23972 ;
    wire new_AGEMA_signal_23973 ;
    wire new_AGEMA_signal_23974 ;
    wire new_AGEMA_signal_23975 ;
    wire new_AGEMA_signal_23976 ;
    wire new_AGEMA_signal_23977 ;
    wire new_AGEMA_signal_23978 ;
    wire new_AGEMA_signal_23979 ;
    wire new_AGEMA_signal_23980 ;
    wire new_AGEMA_signal_23981 ;
    wire new_AGEMA_signal_23982 ;
    wire new_AGEMA_signal_23983 ;
    wire new_AGEMA_signal_23984 ;
    wire new_AGEMA_signal_23985 ;
    wire new_AGEMA_signal_23986 ;
    wire new_AGEMA_signal_23987 ;
    wire new_AGEMA_signal_23988 ;
    wire new_AGEMA_signal_23989 ;
    wire new_AGEMA_signal_23990 ;
    wire new_AGEMA_signal_23991 ;
    wire new_AGEMA_signal_23992 ;
    wire new_AGEMA_signal_23993 ;
    wire new_AGEMA_signal_23994 ;
    wire new_AGEMA_signal_23995 ;
    wire new_AGEMA_signal_23996 ;
    wire new_AGEMA_signal_23997 ;
    wire new_AGEMA_signal_23998 ;
    wire new_AGEMA_signal_23999 ;
    wire new_AGEMA_signal_24000 ;
    wire new_AGEMA_signal_24001 ;
    wire new_AGEMA_signal_24002 ;
    wire new_AGEMA_signal_24003 ;
    wire new_AGEMA_signal_24004 ;
    wire new_AGEMA_signal_24005 ;
    wire new_AGEMA_signal_24006 ;
    wire new_AGEMA_signal_24007 ;
    wire new_AGEMA_signal_24008 ;
    wire new_AGEMA_signal_24009 ;
    wire new_AGEMA_signal_24010 ;
    wire new_AGEMA_signal_24011 ;
    wire new_AGEMA_signal_24012 ;
    wire new_AGEMA_signal_24013 ;
    wire new_AGEMA_signal_24014 ;
    wire new_AGEMA_signal_24015 ;
    wire new_AGEMA_signal_24016 ;
    wire new_AGEMA_signal_24017 ;
    wire new_AGEMA_signal_24018 ;
    wire new_AGEMA_signal_24019 ;
    wire new_AGEMA_signal_24020 ;
    wire new_AGEMA_signal_24021 ;
    wire new_AGEMA_signal_24022 ;
    wire new_AGEMA_signal_24023 ;
    wire new_AGEMA_signal_24024 ;
    wire new_AGEMA_signal_24025 ;
    wire new_AGEMA_signal_24026 ;
    wire new_AGEMA_signal_24027 ;
    wire new_AGEMA_signal_24028 ;
    wire new_AGEMA_signal_24029 ;
    wire new_AGEMA_signal_24030 ;
    wire new_AGEMA_signal_24031 ;
    wire new_AGEMA_signal_24032 ;
    wire new_AGEMA_signal_24033 ;
    wire new_AGEMA_signal_24034 ;
    wire new_AGEMA_signal_24035 ;
    wire new_AGEMA_signal_24036 ;
    wire new_AGEMA_signal_24037 ;
    wire new_AGEMA_signal_24038 ;
    wire new_AGEMA_signal_24039 ;
    wire new_AGEMA_signal_24040 ;
    wire new_AGEMA_signal_24041 ;
    wire new_AGEMA_signal_24042 ;
    wire new_AGEMA_signal_24043 ;
    wire new_AGEMA_signal_24044 ;
    wire new_AGEMA_signal_24045 ;
    wire new_AGEMA_signal_24046 ;
    wire new_AGEMA_signal_24047 ;
    wire new_AGEMA_signal_24048 ;
    wire new_AGEMA_signal_24049 ;
    wire new_AGEMA_signal_24050 ;
    wire new_AGEMA_signal_24051 ;
    wire new_AGEMA_signal_24052 ;
    wire new_AGEMA_signal_24053 ;
    wire new_AGEMA_signal_24054 ;
    wire new_AGEMA_signal_24055 ;
    wire new_AGEMA_signal_24056 ;
    wire new_AGEMA_signal_24057 ;
    wire new_AGEMA_signal_24058 ;
    wire new_AGEMA_signal_24059 ;
    wire new_AGEMA_signal_24060 ;
    wire new_AGEMA_signal_24061 ;
    wire new_AGEMA_signal_24062 ;
    wire new_AGEMA_signal_24063 ;
    wire new_AGEMA_signal_24064 ;
    wire new_AGEMA_signal_24065 ;
    wire new_AGEMA_signal_24066 ;
    wire new_AGEMA_signal_24067 ;
    wire new_AGEMA_signal_24068 ;
    wire new_AGEMA_signal_24069 ;
    wire new_AGEMA_signal_24070 ;
    wire new_AGEMA_signal_24071 ;
    wire new_AGEMA_signal_24072 ;
    wire new_AGEMA_signal_24073 ;
    wire new_AGEMA_signal_24074 ;
    wire new_AGEMA_signal_24075 ;
    wire new_AGEMA_signal_24076 ;
    wire new_AGEMA_signal_24077 ;
    wire new_AGEMA_signal_24078 ;
    wire new_AGEMA_signal_24079 ;
    wire new_AGEMA_signal_24080 ;
    wire new_AGEMA_signal_24081 ;
    wire new_AGEMA_signal_24082 ;
    wire new_AGEMA_signal_24083 ;
    wire new_AGEMA_signal_24084 ;
    wire new_AGEMA_signal_24085 ;
    wire new_AGEMA_signal_24086 ;
    wire new_AGEMA_signal_24087 ;
    wire new_AGEMA_signal_24088 ;
    wire new_AGEMA_signal_24089 ;
    wire new_AGEMA_signal_24090 ;
    wire new_AGEMA_signal_24091 ;
    wire new_AGEMA_signal_24092 ;
    wire new_AGEMA_signal_24093 ;
    wire new_AGEMA_signal_24094 ;
    wire new_AGEMA_signal_24095 ;
    wire new_AGEMA_signal_24096 ;
    wire new_AGEMA_signal_24097 ;
    wire new_AGEMA_signal_24098 ;
    wire new_AGEMA_signal_24099 ;
    wire new_AGEMA_signal_24100 ;
    wire new_AGEMA_signal_24101 ;
    wire new_AGEMA_signal_24102 ;
    wire new_AGEMA_signal_24103 ;
    wire new_AGEMA_signal_24104 ;
    wire new_AGEMA_signal_24105 ;
    wire new_AGEMA_signal_24106 ;
    wire new_AGEMA_signal_24107 ;
    wire new_AGEMA_signal_24108 ;
    wire new_AGEMA_signal_24109 ;
    wire new_AGEMA_signal_24110 ;
    wire new_AGEMA_signal_24111 ;
    wire new_AGEMA_signal_24112 ;
    wire new_AGEMA_signal_24113 ;
    wire new_AGEMA_signal_24114 ;
    wire new_AGEMA_signal_24115 ;
    wire new_AGEMA_signal_24116 ;
    wire new_AGEMA_signal_24117 ;
    wire new_AGEMA_signal_24118 ;
    wire new_AGEMA_signal_24119 ;
    wire new_AGEMA_signal_24120 ;
    wire new_AGEMA_signal_24121 ;
    wire new_AGEMA_signal_24122 ;
    wire new_AGEMA_signal_24123 ;
    wire new_AGEMA_signal_24124 ;
    wire new_AGEMA_signal_24125 ;
    wire new_AGEMA_signal_24126 ;
    wire new_AGEMA_signal_24127 ;
    wire new_AGEMA_signal_24128 ;
    wire new_AGEMA_signal_24129 ;
    wire new_AGEMA_signal_24130 ;
    wire new_AGEMA_signal_24131 ;
    wire new_AGEMA_signal_24132 ;
    wire new_AGEMA_signal_24133 ;
    wire new_AGEMA_signal_24134 ;
    wire new_AGEMA_signal_24135 ;
    wire new_AGEMA_signal_24136 ;
    wire new_AGEMA_signal_24137 ;
    wire new_AGEMA_signal_24138 ;
    wire new_AGEMA_signal_24139 ;
    wire new_AGEMA_signal_24140 ;
    wire new_AGEMA_signal_24141 ;
    wire new_AGEMA_signal_24142 ;
    wire new_AGEMA_signal_24143 ;
    wire new_AGEMA_signal_24144 ;
    wire new_AGEMA_signal_24145 ;
    wire new_AGEMA_signal_24146 ;
    wire new_AGEMA_signal_24147 ;
    wire new_AGEMA_signal_24148 ;
    wire new_AGEMA_signal_24149 ;
    wire new_AGEMA_signal_24150 ;
    wire new_AGEMA_signal_24151 ;
    wire new_AGEMA_signal_24152 ;
    wire new_AGEMA_signal_24153 ;
    wire new_AGEMA_signal_24154 ;
    wire new_AGEMA_signal_24155 ;
    wire new_AGEMA_signal_24156 ;
    wire new_AGEMA_signal_24157 ;
    wire new_AGEMA_signal_24158 ;
    wire new_AGEMA_signal_24159 ;
    wire new_AGEMA_signal_24160 ;
    wire new_AGEMA_signal_24161 ;
    wire new_AGEMA_signal_24162 ;
    wire new_AGEMA_signal_24163 ;
    wire new_AGEMA_signal_24164 ;
    wire new_AGEMA_signal_24165 ;
    wire new_AGEMA_signal_24166 ;
    wire new_AGEMA_signal_24167 ;
    wire new_AGEMA_signal_24168 ;
    wire new_AGEMA_signal_24169 ;
    wire new_AGEMA_signal_24170 ;
    wire new_AGEMA_signal_24171 ;
    wire new_AGEMA_signal_24172 ;
    wire new_AGEMA_signal_24173 ;
    wire new_AGEMA_signal_24174 ;
    wire new_AGEMA_signal_24175 ;
    wire new_AGEMA_signal_24176 ;
    wire new_AGEMA_signal_24177 ;
    wire new_AGEMA_signal_24178 ;
    wire new_AGEMA_signal_24179 ;
    wire new_AGEMA_signal_24180 ;
    wire new_AGEMA_signal_24181 ;
    wire new_AGEMA_signal_24182 ;
    wire new_AGEMA_signal_24183 ;
    wire new_AGEMA_signal_24184 ;
    wire new_AGEMA_signal_24185 ;
    wire new_AGEMA_signal_24186 ;
    wire new_AGEMA_signal_24187 ;
    wire new_AGEMA_signal_24188 ;
    wire new_AGEMA_signal_24189 ;
    wire new_AGEMA_signal_24190 ;
    wire new_AGEMA_signal_24191 ;
    wire new_AGEMA_signal_24192 ;
    wire new_AGEMA_signal_24193 ;
    wire new_AGEMA_signal_24194 ;
    wire new_AGEMA_signal_24195 ;
    wire new_AGEMA_signal_24196 ;
    wire new_AGEMA_signal_24197 ;
    wire new_AGEMA_signal_24198 ;
    wire new_AGEMA_signal_24199 ;
    wire new_AGEMA_signal_24200 ;
    wire new_AGEMA_signal_24201 ;
    wire new_AGEMA_signal_24202 ;
    wire new_AGEMA_signal_24203 ;
    wire new_AGEMA_signal_24204 ;
    wire new_AGEMA_signal_24205 ;
    wire new_AGEMA_signal_24206 ;
    wire new_AGEMA_signal_24207 ;
    wire new_AGEMA_signal_24208 ;
    wire new_AGEMA_signal_24209 ;
    wire new_AGEMA_signal_24210 ;
    wire new_AGEMA_signal_24211 ;
    wire new_AGEMA_signal_24212 ;
    wire new_AGEMA_signal_24213 ;
    wire new_AGEMA_signal_24214 ;
    wire new_AGEMA_signal_24215 ;
    wire new_AGEMA_signal_24216 ;
    wire new_AGEMA_signal_24217 ;
    wire new_AGEMA_signal_24218 ;
    wire new_AGEMA_signal_24219 ;
    wire new_AGEMA_signal_24220 ;
    wire new_AGEMA_signal_24221 ;
    wire new_AGEMA_signal_24222 ;
    wire new_AGEMA_signal_24223 ;
    wire new_AGEMA_signal_24224 ;
    wire new_AGEMA_signal_24225 ;
    wire new_AGEMA_signal_24226 ;
    wire new_AGEMA_signal_24227 ;
    wire new_AGEMA_signal_24228 ;
    wire new_AGEMA_signal_24229 ;
    wire new_AGEMA_signal_24230 ;
    wire new_AGEMA_signal_24231 ;
    wire new_AGEMA_signal_24232 ;
    wire new_AGEMA_signal_24233 ;
    wire new_AGEMA_signal_24234 ;
    wire new_AGEMA_signal_24235 ;
    wire new_AGEMA_signal_24236 ;
    wire new_AGEMA_signal_24237 ;
    wire new_AGEMA_signal_24238 ;
    wire new_AGEMA_signal_24239 ;
    wire new_AGEMA_signal_24240 ;
    wire new_AGEMA_signal_24241 ;
    wire new_AGEMA_signal_24242 ;
    wire new_AGEMA_signal_24243 ;
    wire new_AGEMA_signal_24244 ;
    wire new_AGEMA_signal_24245 ;
    wire new_AGEMA_signal_24246 ;
    wire new_AGEMA_signal_24247 ;
    wire new_AGEMA_signal_24248 ;
    wire new_AGEMA_signal_24249 ;
    wire new_AGEMA_signal_24250 ;
    wire new_AGEMA_signal_24251 ;
    wire new_AGEMA_signal_24252 ;
    wire new_AGEMA_signal_24253 ;
    wire new_AGEMA_signal_24254 ;
    wire new_AGEMA_signal_24255 ;
    wire new_AGEMA_signal_24256 ;
    wire new_AGEMA_signal_24257 ;
    wire new_AGEMA_signal_24258 ;
    wire new_AGEMA_signal_24259 ;
    wire new_AGEMA_signal_24260 ;
    wire new_AGEMA_signal_24261 ;
    wire new_AGEMA_signal_24262 ;
    wire new_AGEMA_signal_24263 ;
    wire new_AGEMA_signal_24264 ;
    wire new_AGEMA_signal_24265 ;
    wire new_AGEMA_signal_24266 ;
    wire new_AGEMA_signal_24267 ;
    wire new_AGEMA_signal_24268 ;
    wire new_AGEMA_signal_24269 ;
    wire new_AGEMA_signal_24270 ;
    wire new_AGEMA_signal_24271 ;
    wire new_AGEMA_signal_24272 ;
    wire new_AGEMA_signal_24273 ;
    wire new_AGEMA_signal_24274 ;
    wire new_AGEMA_signal_24275 ;
    wire new_AGEMA_signal_24276 ;
    wire new_AGEMA_signal_24277 ;
    wire new_AGEMA_signal_24278 ;
    wire new_AGEMA_signal_24279 ;
    wire new_AGEMA_signal_24280 ;
    wire new_AGEMA_signal_24281 ;
    wire new_AGEMA_signal_24282 ;
    wire new_AGEMA_signal_24283 ;
    wire new_AGEMA_signal_24284 ;
    wire new_AGEMA_signal_24285 ;
    wire new_AGEMA_signal_24286 ;
    wire new_AGEMA_signal_24287 ;
    wire new_AGEMA_signal_24288 ;
    wire new_AGEMA_signal_24289 ;
    wire new_AGEMA_signal_24290 ;
    wire new_AGEMA_signal_24291 ;
    wire new_AGEMA_signal_24292 ;
    wire new_AGEMA_signal_24293 ;
    wire new_AGEMA_signal_24294 ;
    wire new_AGEMA_signal_24295 ;
    wire new_AGEMA_signal_24296 ;
    wire new_AGEMA_signal_24297 ;
    wire new_AGEMA_signal_24298 ;
    wire new_AGEMA_signal_24299 ;
    wire new_AGEMA_signal_24300 ;
    wire new_AGEMA_signal_24301 ;
    wire new_AGEMA_signal_24302 ;
    wire new_AGEMA_signal_24303 ;
    wire new_AGEMA_signal_24304 ;
    wire new_AGEMA_signal_24305 ;
    wire new_AGEMA_signal_24306 ;
    wire new_AGEMA_signal_24307 ;
    wire new_AGEMA_signal_24308 ;
    wire new_AGEMA_signal_24309 ;
    wire new_AGEMA_signal_24310 ;
    wire new_AGEMA_signal_24311 ;
    wire new_AGEMA_signal_24312 ;
    wire new_AGEMA_signal_24313 ;
    wire new_AGEMA_signal_24314 ;
    wire new_AGEMA_signal_24315 ;
    wire new_AGEMA_signal_24316 ;
    wire new_AGEMA_signal_24317 ;
    wire new_AGEMA_signal_24318 ;
    wire new_AGEMA_signal_24319 ;
    wire new_AGEMA_signal_24320 ;
    wire new_AGEMA_signal_24321 ;
    wire new_AGEMA_signal_24322 ;
    wire new_AGEMA_signal_24323 ;
    wire new_AGEMA_signal_24324 ;
    wire new_AGEMA_signal_24325 ;
    wire new_AGEMA_signal_24326 ;
    wire new_AGEMA_signal_24327 ;
    wire new_AGEMA_signal_24328 ;
    wire new_AGEMA_signal_24329 ;
    wire new_AGEMA_signal_24330 ;
    wire new_AGEMA_signal_24331 ;
    wire new_AGEMA_signal_24332 ;
    wire new_AGEMA_signal_24333 ;
    wire new_AGEMA_signal_24334 ;
    wire new_AGEMA_signal_24335 ;
    wire new_AGEMA_signal_24336 ;
    wire new_AGEMA_signal_24337 ;
    wire new_AGEMA_signal_24338 ;
    wire new_AGEMA_signal_24339 ;
    wire new_AGEMA_signal_24340 ;
    wire new_AGEMA_signal_24341 ;
    wire new_AGEMA_signal_24342 ;
    wire new_AGEMA_signal_24343 ;
    wire new_AGEMA_signal_24344 ;
    wire new_AGEMA_signal_24345 ;
    wire new_AGEMA_signal_24346 ;
    wire new_AGEMA_signal_24347 ;
    wire new_AGEMA_signal_24348 ;
    wire new_AGEMA_signal_24349 ;
    wire new_AGEMA_signal_24350 ;
    wire new_AGEMA_signal_24351 ;
    wire new_AGEMA_signal_24352 ;
    wire new_AGEMA_signal_24353 ;
    wire new_AGEMA_signal_24354 ;
    wire new_AGEMA_signal_24355 ;
    wire new_AGEMA_signal_24356 ;
    wire new_AGEMA_signal_24357 ;
    wire new_AGEMA_signal_24358 ;
    wire new_AGEMA_signal_24359 ;
    wire new_AGEMA_signal_24360 ;
    wire new_AGEMA_signal_24361 ;
    wire new_AGEMA_signal_24362 ;
    wire new_AGEMA_signal_24363 ;
    wire new_AGEMA_signal_24364 ;
    wire new_AGEMA_signal_24365 ;
    wire new_AGEMA_signal_24366 ;
    wire new_AGEMA_signal_24367 ;
    wire new_AGEMA_signal_24368 ;
    wire new_AGEMA_signal_24369 ;
    wire new_AGEMA_signal_24370 ;
    wire new_AGEMA_signal_24371 ;
    wire new_AGEMA_signal_24372 ;
    wire new_AGEMA_signal_24373 ;
    wire new_AGEMA_signal_24374 ;
    wire new_AGEMA_signal_24375 ;
    wire new_AGEMA_signal_24376 ;
    wire new_AGEMA_signal_24377 ;
    wire new_AGEMA_signal_24378 ;
    wire new_AGEMA_signal_24379 ;
    wire new_AGEMA_signal_24380 ;
    wire new_AGEMA_signal_24381 ;
    wire new_AGEMA_signal_24382 ;
    wire new_AGEMA_signal_24383 ;
    wire new_AGEMA_signal_24384 ;
    wire new_AGEMA_signal_24385 ;
    wire new_AGEMA_signal_24386 ;
    wire new_AGEMA_signal_24387 ;
    wire new_AGEMA_signal_24388 ;
    wire new_AGEMA_signal_24389 ;
    wire new_AGEMA_signal_24390 ;
    wire new_AGEMA_signal_24391 ;
    wire new_AGEMA_signal_24392 ;
    wire new_AGEMA_signal_24393 ;
    wire new_AGEMA_signal_24394 ;
    wire new_AGEMA_signal_24395 ;
    wire new_AGEMA_signal_24396 ;
    wire new_AGEMA_signal_24397 ;
    wire new_AGEMA_signal_24398 ;
    wire new_AGEMA_signal_24399 ;
    wire new_AGEMA_signal_24400 ;
    wire new_AGEMA_signal_24401 ;
    wire new_AGEMA_signal_24402 ;
    wire new_AGEMA_signal_24403 ;
    wire new_AGEMA_signal_24404 ;
    wire new_AGEMA_signal_24405 ;
    wire new_AGEMA_signal_24406 ;
    wire new_AGEMA_signal_24407 ;
    wire new_AGEMA_signal_24408 ;
    wire new_AGEMA_signal_24409 ;
    wire new_AGEMA_signal_24410 ;
    wire new_AGEMA_signal_24411 ;
    wire new_AGEMA_signal_24412 ;
    wire new_AGEMA_signal_24413 ;
    wire new_AGEMA_signal_24414 ;
    wire new_AGEMA_signal_24415 ;
    wire new_AGEMA_signal_24416 ;
    wire new_AGEMA_signal_24417 ;
    wire new_AGEMA_signal_24418 ;
    wire new_AGEMA_signal_24419 ;
    wire new_AGEMA_signal_24420 ;
    wire new_AGEMA_signal_24421 ;
    wire new_AGEMA_signal_24422 ;
    wire new_AGEMA_signal_24423 ;
    wire new_AGEMA_signal_24424 ;
    wire new_AGEMA_signal_24425 ;
    wire new_AGEMA_signal_24426 ;
    wire new_AGEMA_signal_24427 ;
    wire new_AGEMA_signal_24428 ;
    wire new_AGEMA_signal_24429 ;
    wire new_AGEMA_signal_24430 ;
    wire new_AGEMA_signal_24431 ;
    wire new_AGEMA_signal_24432 ;
    wire new_AGEMA_signal_24433 ;
    wire new_AGEMA_signal_24434 ;
    wire new_AGEMA_signal_24435 ;
    wire new_AGEMA_signal_24436 ;
    wire new_AGEMA_signal_24437 ;
    wire new_AGEMA_signal_24438 ;
    wire new_AGEMA_signal_24439 ;
    wire new_AGEMA_signal_24440 ;
    wire new_AGEMA_signal_24441 ;
    wire new_AGEMA_signal_24442 ;
    wire new_AGEMA_signal_24443 ;
    wire new_AGEMA_signal_24444 ;
    wire new_AGEMA_signal_24445 ;
    wire new_AGEMA_signal_24446 ;
    wire new_AGEMA_signal_24447 ;
    wire new_AGEMA_signal_24448 ;
    wire new_AGEMA_signal_24449 ;
    wire new_AGEMA_signal_24450 ;
    wire new_AGEMA_signal_24451 ;
    wire new_AGEMA_signal_24452 ;
    wire new_AGEMA_signal_24453 ;
    wire new_AGEMA_signal_24454 ;
    wire new_AGEMA_signal_24455 ;
    wire new_AGEMA_signal_24456 ;
    wire new_AGEMA_signal_24457 ;
    wire new_AGEMA_signal_24458 ;
    wire new_AGEMA_signal_24459 ;
    wire new_AGEMA_signal_24460 ;
    wire new_AGEMA_signal_24461 ;
    wire new_AGEMA_signal_24462 ;
    wire new_AGEMA_signal_24463 ;
    wire new_AGEMA_signal_24464 ;
    wire new_AGEMA_signal_24465 ;
    wire new_AGEMA_signal_24466 ;
    wire new_AGEMA_signal_24467 ;
    wire new_AGEMA_signal_24468 ;
    wire new_AGEMA_signal_24469 ;
    wire new_AGEMA_signal_24470 ;
    wire new_AGEMA_signal_24471 ;
    wire new_AGEMA_signal_24472 ;
    wire new_AGEMA_signal_24473 ;
    wire new_AGEMA_signal_24474 ;
    wire new_AGEMA_signal_24475 ;
    wire new_AGEMA_signal_24476 ;
    wire new_AGEMA_signal_24477 ;
    wire new_AGEMA_signal_24478 ;
    wire new_AGEMA_signal_24479 ;
    wire new_AGEMA_signal_24480 ;
    wire new_AGEMA_signal_24481 ;
    wire new_AGEMA_signal_24482 ;
    wire new_AGEMA_signal_24483 ;
    wire new_AGEMA_signal_24484 ;
    wire new_AGEMA_signal_24485 ;
    wire new_AGEMA_signal_24486 ;
    wire new_AGEMA_signal_24487 ;
    wire new_AGEMA_signal_24488 ;
    wire new_AGEMA_signal_24489 ;
    wire new_AGEMA_signal_24490 ;
    wire new_AGEMA_signal_24491 ;
    wire new_AGEMA_signal_24492 ;
    wire new_AGEMA_signal_24493 ;
    wire new_AGEMA_signal_24494 ;
    wire new_AGEMA_signal_24495 ;
    wire new_AGEMA_signal_24496 ;
    wire new_AGEMA_signal_24497 ;
    wire new_AGEMA_signal_24498 ;
    wire new_AGEMA_signal_24499 ;
    wire new_AGEMA_signal_24500 ;
    wire new_AGEMA_signal_24501 ;
    wire new_AGEMA_signal_24502 ;
    wire new_AGEMA_signal_24503 ;
    wire new_AGEMA_signal_24504 ;
    wire new_AGEMA_signal_24505 ;
    wire new_AGEMA_signal_24506 ;
    wire new_AGEMA_signal_24507 ;
    wire new_AGEMA_signal_24508 ;
    wire new_AGEMA_signal_24509 ;
    wire new_AGEMA_signal_24510 ;
    wire new_AGEMA_signal_24511 ;
    wire new_AGEMA_signal_24512 ;
    wire new_AGEMA_signal_24513 ;
    wire new_AGEMA_signal_24514 ;
    wire new_AGEMA_signal_24515 ;
    wire new_AGEMA_signal_24516 ;
    wire new_AGEMA_signal_24517 ;
    wire new_AGEMA_signal_24518 ;
    wire new_AGEMA_signal_24519 ;
    wire new_AGEMA_signal_24520 ;
    wire new_AGEMA_signal_24521 ;
    wire new_AGEMA_signal_24522 ;
    wire new_AGEMA_signal_24523 ;
    wire new_AGEMA_signal_24524 ;
    wire new_AGEMA_signal_24525 ;
    wire new_AGEMA_signal_24526 ;
    wire new_AGEMA_signal_24527 ;
    wire new_AGEMA_signal_24528 ;
    wire new_AGEMA_signal_24529 ;
    wire new_AGEMA_signal_24530 ;
    wire new_AGEMA_signal_24531 ;
    wire new_AGEMA_signal_24532 ;
    wire new_AGEMA_signal_24533 ;
    wire new_AGEMA_signal_24534 ;
    wire new_AGEMA_signal_24535 ;
    wire new_AGEMA_signal_24536 ;
    wire new_AGEMA_signal_24537 ;
    wire new_AGEMA_signal_24538 ;
    wire new_AGEMA_signal_24539 ;
    wire new_AGEMA_signal_24540 ;
    wire new_AGEMA_signal_24541 ;
    wire new_AGEMA_signal_24542 ;
    wire new_AGEMA_signal_24543 ;
    wire new_AGEMA_signal_24544 ;
    wire new_AGEMA_signal_24545 ;
    wire new_AGEMA_signal_24546 ;
    wire new_AGEMA_signal_24547 ;
    wire new_AGEMA_signal_24548 ;
    wire new_AGEMA_signal_24549 ;
    wire new_AGEMA_signal_24550 ;
    wire new_AGEMA_signal_24551 ;
    wire new_AGEMA_signal_24552 ;
    wire new_AGEMA_signal_24553 ;
    wire new_AGEMA_signal_24554 ;
    wire new_AGEMA_signal_24555 ;
    wire new_AGEMA_signal_24556 ;
    wire new_AGEMA_signal_24557 ;
    wire new_AGEMA_signal_24558 ;
    wire new_AGEMA_signal_24559 ;
    wire new_AGEMA_signal_24560 ;
    wire new_AGEMA_signal_24561 ;
    wire new_AGEMA_signal_24562 ;
    wire new_AGEMA_signal_24563 ;
    wire new_AGEMA_signal_24564 ;
    wire new_AGEMA_signal_24565 ;
    wire new_AGEMA_signal_24566 ;
    wire new_AGEMA_signal_24567 ;
    wire new_AGEMA_signal_24568 ;
    wire new_AGEMA_signal_24569 ;
    wire new_AGEMA_signal_24570 ;
    wire new_AGEMA_signal_24571 ;
    wire new_AGEMA_signal_24572 ;
    wire new_AGEMA_signal_24573 ;
    wire new_AGEMA_signal_24574 ;
    wire new_AGEMA_signal_24575 ;
    wire new_AGEMA_signal_24576 ;
    wire new_AGEMA_signal_24577 ;
    wire new_AGEMA_signal_24578 ;
    wire new_AGEMA_signal_24579 ;
    wire new_AGEMA_signal_24580 ;
    wire new_AGEMA_signal_24581 ;
    wire new_AGEMA_signal_24582 ;
    wire new_AGEMA_signal_24583 ;
    wire new_AGEMA_signal_24584 ;
    wire new_AGEMA_signal_24585 ;
    wire new_AGEMA_signal_24586 ;
    wire new_AGEMA_signal_24587 ;
    wire new_AGEMA_signal_24588 ;
    wire new_AGEMA_signal_24589 ;
    wire new_AGEMA_signal_24590 ;
    wire new_AGEMA_signal_24591 ;
    wire new_AGEMA_signal_24592 ;
    wire new_AGEMA_signal_24593 ;
    wire new_AGEMA_signal_24594 ;
    wire new_AGEMA_signal_24595 ;
    wire new_AGEMA_signal_24596 ;
    wire new_AGEMA_signal_24597 ;
    wire new_AGEMA_signal_24598 ;
    wire new_AGEMA_signal_24599 ;
    wire new_AGEMA_signal_24600 ;
    wire new_AGEMA_signal_24601 ;
    wire new_AGEMA_signal_24602 ;
    wire new_AGEMA_signal_24603 ;
    wire new_AGEMA_signal_24604 ;
    wire new_AGEMA_signal_24605 ;
    wire new_AGEMA_signal_24606 ;
    wire new_AGEMA_signal_24607 ;
    wire new_AGEMA_signal_24608 ;
    wire new_AGEMA_signal_24609 ;
    wire new_AGEMA_signal_24610 ;
    wire new_AGEMA_signal_24611 ;
    wire new_AGEMA_signal_24612 ;
    wire new_AGEMA_signal_24613 ;
    wire new_AGEMA_signal_24614 ;
    wire new_AGEMA_signal_24615 ;
    wire new_AGEMA_signal_24616 ;
    wire new_AGEMA_signal_24617 ;
    wire new_AGEMA_signal_24618 ;
    wire new_AGEMA_signal_24619 ;
    wire new_AGEMA_signal_24620 ;
    wire new_AGEMA_signal_24621 ;
    wire new_AGEMA_signal_24622 ;
    wire new_AGEMA_signal_24623 ;
    wire new_AGEMA_signal_24624 ;
    wire new_AGEMA_signal_24625 ;
    wire new_AGEMA_signal_24626 ;
    wire new_AGEMA_signal_24627 ;
    wire new_AGEMA_signal_24628 ;
    wire new_AGEMA_signal_24629 ;
    wire new_AGEMA_signal_24630 ;
    wire new_AGEMA_signal_24631 ;
    wire new_AGEMA_signal_24632 ;
    wire new_AGEMA_signal_24633 ;
    wire new_AGEMA_signal_24634 ;
    wire new_AGEMA_signal_24635 ;
    wire new_AGEMA_signal_24636 ;
    wire new_AGEMA_signal_24637 ;
    wire new_AGEMA_signal_24638 ;
    wire new_AGEMA_signal_24639 ;
    wire new_AGEMA_signal_24640 ;
    wire new_AGEMA_signal_24641 ;
    wire new_AGEMA_signal_24642 ;
    wire new_AGEMA_signal_24643 ;
    wire new_AGEMA_signal_24644 ;
    wire new_AGEMA_signal_24645 ;
    wire new_AGEMA_signal_24646 ;
    wire new_AGEMA_signal_24647 ;
    wire new_AGEMA_signal_24648 ;
    wire new_AGEMA_signal_24649 ;
    wire new_AGEMA_signal_24650 ;
    wire new_AGEMA_signal_24651 ;
    wire new_AGEMA_signal_24652 ;
    wire new_AGEMA_signal_24653 ;
    wire new_AGEMA_signal_24654 ;
    wire new_AGEMA_signal_24655 ;
    wire new_AGEMA_signal_24656 ;
    wire new_AGEMA_signal_24657 ;
    wire new_AGEMA_signal_24658 ;
    wire new_AGEMA_signal_24659 ;
    wire new_AGEMA_signal_24660 ;
    wire new_AGEMA_signal_24661 ;
    wire new_AGEMA_signal_24662 ;
    wire new_AGEMA_signal_24663 ;
    wire new_AGEMA_signal_24664 ;
    wire new_AGEMA_signal_24665 ;
    wire new_AGEMA_signal_24666 ;
    wire new_AGEMA_signal_24667 ;
    wire new_AGEMA_signal_24668 ;
    wire new_AGEMA_signal_24669 ;
    wire new_AGEMA_signal_24670 ;
    wire new_AGEMA_signal_24671 ;
    wire new_AGEMA_signal_24672 ;
    wire new_AGEMA_signal_24673 ;
    wire new_AGEMA_signal_24674 ;
    wire new_AGEMA_signal_24675 ;
    wire new_AGEMA_signal_24676 ;
    wire new_AGEMA_signal_24677 ;
    wire new_AGEMA_signal_24678 ;
    wire new_AGEMA_signal_24679 ;
    wire new_AGEMA_signal_24680 ;
    wire new_AGEMA_signal_24681 ;
    wire new_AGEMA_signal_24682 ;
    wire new_AGEMA_signal_24683 ;
    wire new_AGEMA_signal_24684 ;
    wire new_AGEMA_signal_24685 ;
    wire new_AGEMA_signal_24686 ;
    wire new_AGEMA_signal_24687 ;
    wire new_AGEMA_signal_24688 ;
    wire new_AGEMA_signal_24689 ;
    wire new_AGEMA_signal_24690 ;
    wire new_AGEMA_signal_24691 ;
    wire new_AGEMA_signal_24692 ;
    wire new_AGEMA_signal_24693 ;
    wire new_AGEMA_signal_24694 ;
    wire new_AGEMA_signal_24695 ;
    wire new_AGEMA_signal_24696 ;
    wire new_AGEMA_signal_24697 ;
    wire new_AGEMA_signal_24698 ;
    wire new_AGEMA_signal_24699 ;
    wire new_AGEMA_signal_24700 ;
    wire new_AGEMA_signal_24701 ;
    wire new_AGEMA_signal_24702 ;
    wire new_AGEMA_signal_24703 ;
    wire new_AGEMA_signal_24704 ;
    wire new_AGEMA_signal_24705 ;
    wire new_AGEMA_signal_24706 ;
    wire new_AGEMA_signal_24707 ;
    wire new_AGEMA_signal_24708 ;
    wire new_AGEMA_signal_24709 ;
    wire new_AGEMA_signal_24710 ;
    wire new_AGEMA_signal_24711 ;
    wire new_AGEMA_signal_24712 ;
    wire new_AGEMA_signal_24713 ;
    wire new_AGEMA_signal_24714 ;
    wire new_AGEMA_signal_24715 ;
    wire new_AGEMA_signal_24716 ;
    wire new_AGEMA_signal_24717 ;
    wire new_AGEMA_signal_24718 ;
    wire new_AGEMA_signal_24719 ;
    wire new_AGEMA_signal_24720 ;
    wire new_AGEMA_signal_24721 ;
    wire new_AGEMA_signal_24722 ;
    wire new_AGEMA_signal_24723 ;
    wire new_AGEMA_signal_24724 ;
    wire new_AGEMA_signal_24725 ;
    wire new_AGEMA_signal_24726 ;
    wire new_AGEMA_signal_24727 ;
    wire new_AGEMA_signal_24728 ;
    wire new_AGEMA_signal_24729 ;
    wire new_AGEMA_signal_24730 ;
    wire new_AGEMA_signal_24731 ;
    wire new_AGEMA_signal_24732 ;
    wire new_AGEMA_signal_24733 ;
    wire new_AGEMA_signal_24734 ;
    wire new_AGEMA_signal_24735 ;
    wire new_AGEMA_signal_24736 ;
    wire new_AGEMA_signal_24737 ;
    wire new_AGEMA_signal_24738 ;
    wire new_AGEMA_signal_24739 ;
    wire new_AGEMA_signal_24740 ;
    wire new_AGEMA_signal_24741 ;
    wire new_AGEMA_signal_24742 ;
    wire new_AGEMA_signal_24743 ;
    wire new_AGEMA_signal_24744 ;
    wire new_AGEMA_signal_24745 ;
    wire new_AGEMA_signal_24746 ;
    wire new_AGEMA_signal_24747 ;
    wire new_AGEMA_signal_24748 ;
    wire new_AGEMA_signal_24749 ;
    wire new_AGEMA_signal_24750 ;
    wire new_AGEMA_signal_24751 ;
    wire new_AGEMA_signal_24752 ;
    wire new_AGEMA_signal_24753 ;
    wire new_AGEMA_signal_24754 ;
    wire new_AGEMA_signal_24755 ;
    wire new_AGEMA_signal_24756 ;
    wire new_AGEMA_signal_24757 ;
    wire new_AGEMA_signal_24758 ;
    wire new_AGEMA_signal_24759 ;
    wire new_AGEMA_signal_24760 ;
    wire new_AGEMA_signal_24761 ;
    wire new_AGEMA_signal_24762 ;
    wire new_AGEMA_signal_24763 ;
    wire new_AGEMA_signal_24764 ;
    wire new_AGEMA_signal_24765 ;
    wire new_AGEMA_signal_24766 ;
    wire new_AGEMA_signal_24767 ;
    wire new_AGEMA_signal_24768 ;
    wire new_AGEMA_signal_24769 ;
    wire new_AGEMA_signal_24770 ;
    wire new_AGEMA_signal_24771 ;
    wire new_AGEMA_signal_24772 ;
    wire new_AGEMA_signal_24773 ;
    wire new_AGEMA_signal_24774 ;
    wire new_AGEMA_signal_24775 ;
    wire new_AGEMA_signal_24776 ;
    wire new_AGEMA_signal_24777 ;
    wire new_AGEMA_signal_24778 ;
    wire new_AGEMA_signal_24779 ;
    wire new_AGEMA_signal_24780 ;
    wire new_AGEMA_signal_24781 ;
    wire new_AGEMA_signal_24782 ;
    wire new_AGEMA_signal_24783 ;
    wire new_AGEMA_signal_24784 ;
    wire new_AGEMA_signal_24785 ;
    wire new_AGEMA_signal_24786 ;
    wire new_AGEMA_signal_24787 ;
    wire new_AGEMA_signal_24788 ;
    wire new_AGEMA_signal_24789 ;
    wire new_AGEMA_signal_24790 ;
    wire new_AGEMA_signal_24791 ;
    wire new_AGEMA_signal_24792 ;
    wire new_AGEMA_signal_24793 ;
    wire new_AGEMA_signal_24794 ;
    wire new_AGEMA_signal_24795 ;
    wire new_AGEMA_signal_24796 ;
    wire new_AGEMA_signal_24797 ;
    wire new_AGEMA_signal_24798 ;
    wire new_AGEMA_signal_24799 ;
    wire new_AGEMA_signal_24800 ;
    wire new_AGEMA_signal_24801 ;
    wire new_AGEMA_signal_24802 ;
    wire new_AGEMA_signal_24803 ;
    wire new_AGEMA_signal_24804 ;
    wire new_AGEMA_signal_24805 ;
    wire new_AGEMA_signal_24806 ;
    wire new_AGEMA_signal_24807 ;
    wire new_AGEMA_signal_24808 ;
    wire new_AGEMA_signal_24809 ;
    wire new_AGEMA_signal_24810 ;
    wire new_AGEMA_signal_24811 ;
    wire new_AGEMA_signal_24812 ;
    wire new_AGEMA_signal_24813 ;
    wire new_AGEMA_signal_24814 ;
    wire new_AGEMA_signal_24815 ;
    wire new_AGEMA_signal_24816 ;
    wire new_AGEMA_signal_24817 ;
    wire new_AGEMA_signal_24818 ;
    wire new_AGEMA_signal_24819 ;
    wire new_AGEMA_signal_24820 ;
    wire new_AGEMA_signal_24821 ;
    wire new_AGEMA_signal_24822 ;
    wire new_AGEMA_signal_24823 ;
    wire new_AGEMA_signal_24824 ;
    wire new_AGEMA_signal_24825 ;
    wire new_AGEMA_signal_24826 ;
    wire new_AGEMA_signal_24827 ;
    wire new_AGEMA_signal_24828 ;
    wire new_AGEMA_signal_24829 ;
    wire new_AGEMA_signal_24830 ;
    wire new_AGEMA_signal_24831 ;
    wire new_AGEMA_signal_24832 ;
    wire new_AGEMA_signal_24833 ;
    wire new_AGEMA_signal_24834 ;
    wire new_AGEMA_signal_24835 ;
    wire new_AGEMA_signal_24836 ;
    wire new_AGEMA_signal_24837 ;
    wire new_AGEMA_signal_24838 ;
    wire new_AGEMA_signal_24839 ;
    wire new_AGEMA_signal_24840 ;
    wire new_AGEMA_signal_24841 ;
    wire new_AGEMA_signal_24842 ;
    wire new_AGEMA_signal_24843 ;
    wire new_AGEMA_signal_24844 ;
    wire new_AGEMA_signal_24845 ;
    wire new_AGEMA_signal_24846 ;
    wire new_AGEMA_signal_24847 ;
    wire new_AGEMA_signal_24848 ;
    wire new_AGEMA_signal_24849 ;
    wire new_AGEMA_signal_24850 ;
    wire new_AGEMA_signal_24851 ;
    wire new_AGEMA_signal_24852 ;
    wire new_AGEMA_signal_24853 ;
    wire new_AGEMA_signal_24854 ;
    wire new_AGEMA_signal_24855 ;
    wire new_AGEMA_signal_24856 ;
    wire new_AGEMA_signal_24857 ;
    wire new_AGEMA_signal_24858 ;
    wire new_AGEMA_signal_24859 ;
    wire new_AGEMA_signal_24860 ;
    wire new_AGEMA_signal_24861 ;
    wire new_AGEMA_signal_24862 ;
    wire new_AGEMA_signal_24863 ;
    wire new_AGEMA_signal_24864 ;
    wire new_AGEMA_signal_24865 ;
    wire new_AGEMA_signal_24866 ;
    wire new_AGEMA_signal_24867 ;
    wire new_AGEMA_signal_24868 ;
    wire new_AGEMA_signal_24869 ;
    wire new_AGEMA_signal_24870 ;
    wire new_AGEMA_signal_24871 ;
    wire new_AGEMA_signal_24872 ;
    wire new_AGEMA_signal_24873 ;
    wire new_AGEMA_signal_24874 ;
    wire new_AGEMA_signal_24875 ;
    wire new_AGEMA_signal_24876 ;
    wire new_AGEMA_signal_24877 ;
    wire new_AGEMA_signal_24878 ;
    wire new_AGEMA_signal_24879 ;
    wire new_AGEMA_signal_24880 ;
    wire new_AGEMA_signal_24881 ;
    wire new_AGEMA_signal_24882 ;
    wire new_AGEMA_signal_24883 ;
    wire new_AGEMA_signal_24884 ;
    wire new_AGEMA_signal_24885 ;
    wire new_AGEMA_signal_24886 ;
    wire new_AGEMA_signal_24887 ;
    wire new_AGEMA_signal_24888 ;
    wire new_AGEMA_signal_24889 ;
    wire new_AGEMA_signal_24890 ;
    wire new_AGEMA_signal_24891 ;
    wire new_AGEMA_signal_24892 ;
    wire new_AGEMA_signal_24893 ;
    wire new_AGEMA_signal_24894 ;
    wire new_AGEMA_signal_24895 ;
    wire new_AGEMA_signal_24896 ;
    wire new_AGEMA_signal_24897 ;
    wire new_AGEMA_signal_24898 ;
    wire new_AGEMA_signal_24899 ;
    wire new_AGEMA_signal_24900 ;
    wire new_AGEMA_signal_24901 ;
    wire new_AGEMA_signal_24902 ;
    wire new_AGEMA_signal_24903 ;
    wire new_AGEMA_signal_24904 ;
    wire new_AGEMA_signal_24905 ;
    wire new_AGEMA_signal_24906 ;
    wire new_AGEMA_signal_24907 ;
    wire new_AGEMA_signal_24908 ;
    wire new_AGEMA_signal_24909 ;
    wire new_AGEMA_signal_24910 ;
    wire new_AGEMA_signal_24911 ;
    wire new_AGEMA_signal_24912 ;
    wire new_AGEMA_signal_24913 ;
    wire new_AGEMA_signal_24914 ;
    wire new_AGEMA_signal_24915 ;
    wire new_AGEMA_signal_24916 ;
    wire new_AGEMA_signal_24917 ;
    wire new_AGEMA_signal_24918 ;
    wire new_AGEMA_signal_24919 ;
    wire new_AGEMA_signal_24920 ;
    wire new_AGEMA_signal_24921 ;
    wire new_AGEMA_signal_24922 ;
    wire new_AGEMA_signal_24923 ;
    wire new_AGEMA_signal_24924 ;
    wire new_AGEMA_signal_24925 ;
    wire new_AGEMA_signal_24926 ;
    wire new_AGEMA_signal_24927 ;
    wire new_AGEMA_signal_24928 ;
    wire new_AGEMA_signal_24929 ;
    wire new_AGEMA_signal_24930 ;
    wire new_AGEMA_signal_24931 ;
    wire new_AGEMA_signal_24932 ;
    wire new_AGEMA_signal_24933 ;
    wire new_AGEMA_signal_24934 ;
    wire new_AGEMA_signal_24935 ;
    wire new_AGEMA_signal_24936 ;
    wire new_AGEMA_signal_24937 ;
    wire new_AGEMA_signal_24938 ;
    wire new_AGEMA_signal_24939 ;
    wire new_AGEMA_signal_24940 ;
    wire new_AGEMA_signal_24941 ;
    wire new_AGEMA_signal_24942 ;
    wire new_AGEMA_signal_24943 ;
    wire new_AGEMA_signal_24944 ;
    wire new_AGEMA_signal_24945 ;
    wire new_AGEMA_signal_24946 ;
    wire new_AGEMA_signal_24947 ;
    wire new_AGEMA_signal_24948 ;
    wire new_AGEMA_signal_24949 ;
    wire new_AGEMA_signal_24950 ;
    wire new_AGEMA_signal_24951 ;
    wire new_AGEMA_signal_24952 ;
    wire new_AGEMA_signal_24953 ;
    wire new_AGEMA_signal_24954 ;
    wire new_AGEMA_signal_24955 ;
    wire new_AGEMA_signal_24956 ;
    wire new_AGEMA_signal_24957 ;
    wire new_AGEMA_signal_24958 ;
    wire new_AGEMA_signal_24959 ;
    wire new_AGEMA_signal_24960 ;
    wire new_AGEMA_signal_24961 ;
    wire new_AGEMA_signal_24962 ;
    wire new_AGEMA_signal_24963 ;
    wire new_AGEMA_signal_24964 ;
    wire new_AGEMA_signal_24965 ;
    wire new_AGEMA_signal_24966 ;
    wire new_AGEMA_signal_24967 ;
    wire new_AGEMA_signal_24968 ;
    wire new_AGEMA_signal_24969 ;
    wire new_AGEMA_signal_24970 ;
    wire new_AGEMA_signal_24971 ;
    wire new_AGEMA_signal_24972 ;
    wire new_AGEMA_signal_24973 ;
    wire new_AGEMA_signal_24974 ;
    wire new_AGEMA_signal_24975 ;
    wire new_AGEMA_signal_24976 ;
    wire new_AGEMA_signal_24977 ;
    wire new_AGEMA_signal_24978 ;
    wire new_AGEMA_signal_24979 ;
    wire new_AGEMA_signal_24980 ;
    wire new_AGEMA_signal_24981 ;
    wire new_AGEMA_signal_24982 ;
    wire new_AGEMA_signal_24983 ;
    wire new_AGEMA_signal_24984 ;
    wire new_AGEMA_signal_24985 ;
    wire new_AGEMA_signal_24986 ;
    wire new_AGEMA_signal_24987 ;
    wire new_AGEMA_signal_24988 ;
    wire new_AGEMA_signal_24989 ;
    wire new_AGEMA_signal_24990 ;
    wire new_AGEMA_signal_24991 ;
    wire new_AGEMA_signal_24992 ;
    wire new_AGEMA_signal_24993 ;
    wire new_AGEMA_signal_24994 ;
    wire new_AGEMA_signal_24995 ;
    wire new_AGEMA_signal_24996 ;
    wire new_AGEMA_signal_24997 ;
    wire new_AGEMA_signal_24998 ;
    wire new_AGEMA_signal_24999 ;
    wire new_AGEMA_signal_25000 ;
    wire new_AGEMA_signal_25001 ;
    wire new_AGEMA_signal_25002 ;
    wire new_AGEMA_signal_25003 ;
    wire new_AGEMA_signal_25004 ;
    wire new_AGEMA_signal_25005 ;
    wire new_AGEMA_signal_25006 ;
    wire new_AGEMA_signal_25007 ;
    wire new_AGEMA_signal_25008 ;
    wire new_AGEMA_signal_25009 ;
    wire new_AGEMA_signal_25010 ;
    wire new_AGEMA_signal_25011 ;
    wire new_AGEMA_signal_25012 ;
    wire new_AGEMA_signal_25013 ;
    wire new_AGEMA_signal_25014 ;
    wire new_AGEMA_signal_25015 ;
    wire new_AGEMA_signal_25016 ;
    wire new_AGEMA_signal_25017 ;
    wire new_AGEMA_signal_25018 ;
    wire new_AGEMA_signal_25019 ;
    wire new_AGEMA_signal_25020 ;
    wire new_AGEMA_signal_25021 ;
    wire new_AGEMA_signal_25022 ;
    wire new_AGEMA_signal_25023 ;
    wire new_AGEMA_signal_25024 ;
    wire new_AGEMA_signal_25025 ;
    wire new_AGEMA_signal_25026 ;
    wire new_AGEMA_signal_25027 ;
    wire new_AGEMA_signal_25028 ;
    wire new_AGEMA_signal_25029 ;
    wire new_AGEMA_signal_25030 ;
    wire new_AGEMA_signal_25031 ;
    wire new_AGEMA_signal_25032 ;
    wire new_AGEMA_signal_25033 ;
    wire new_AGEMA_signal_25034 ;
    wire new_AGEMA_signal_25035 ;
    wire new_AGEMA_signal_25036 ;
    wire new_AGEMA_signal_25037 ;
    wire new_AGEMA_signal_25038 ;
    wire new_AGEMA_signal_25039 ;
    wire new_AGEMA_signal_25040 ;
    wire new_AGEMA_signal_25041 ;
    wire new_AGEMA_signal_25042 ;
    wire new_AGEMA_signal_25043 ;
    wire new_AGEMA_signal_25044 ;
    wire new_AGEMA_signal_25045 ;
    wire new_AGEMA_signal_25046 ;
    wire new_AGEMA_signal_25047 ;
    wire new_AGEMA_signal_25048 ;
    wire new_AGEMA_signal_25049 ;
    wire new_AGEMA_signal_25050 ;
    wire new_AGEMA_signal_25051 ;
    wire new_AGEMA_signal_25052 ;
    wire new_AGEMA_signal_25053 ;
    wire new_AGEMA_signal_25054 ;
    wire new_AGEMA_signal_25055 ;
    wire new_AGEMA_signal_25056 ;
    wire new_AGEMA_signal_25057 ;
    wire new_AGEMA_signal_25058 ;
    wire new_AGEMA_signal_25059 ;
    wire new_AGEMA_signal_25060 ;
    wire new_AGEMA_signal_25061 ;
    wire new_AGEMA_signal_25062 ;
    wire new_AGEMA_signal_25063 ;
    wire new_AGEMA_signal_25064 ;
    wire new_AGEMA_signal_25065 ;
    wire new_AGEMA_signal_25066 ;
    wire new_AGEMA_signal_25067 ;
    wire new_AGEMA_signal_25068 ;
    wire new_AGEMA_signal_25069 ;
    wire new_AGEMA_signal_25070 ;
    wire new_AGEMA_signal_25071 ;
    wire new_AGEMA_signal_25072 ;
    wire new_AGEMA_signal_25073 ;
    wire new_AGEMA_signal_25074 ;
    wire new_AGEMA_signal_25075 ;
    wire new_AGEMA_signal_25076 ;
    wire new_AGEMA_signal_25077 ;
    wire new_AGEMA_signal_25078 ;
    wire new_AGEMA_signal_25079 ;
    wire new_AGEMA_signal_25080 ;
    wire new_AGEMA_signal_25081 ;
    wire new_AGEMA_signal_25082 ;
    wire new_AGEMA_signal_25083 ;
    wire new_AGEMA_signal_25084 ;
    wire new_AGEMA_signal_25085 ;
    wire new_AGEMA_signal_25086 ;
    wire new_AGEMA_signal_25087 ;
    wire new_AGEMA_signal_25088 ;
    wire new_AGEMA_signal_25089 ;
    wire new_AGEMA_signal_25090 ;
    wire new_AGEMA_signal_25091 ;
    wire new_AGEMA_signal_25092 ;
    wire new_AGEMA_signal_25093 ;
    wire new_AGEMA_signal_25094 ;
    wire new_AGEMA_signal_25095 ;
    wire new_AGEMA_signal_25096 ;
    wire new_AGEMA_signal_25097 ;
    wire new_AGEMA_signal_25098 ;
    wire new_AGEMA_signal_25099 ;
    wire new_AGEMA_signal_25100 ;
    wire new_AGEMA_signal_25101 ;
    wire new_AGEMA_signal_25102 ;
    wire new_AGEMA_signal_25103 ;
    wire new_AGEMA_signal_25104 ;
    wire new_AGEMA_signal_25105 ;
    wire new_AGEMA_signal_25106 ;
    wire new_AGEMA_signal_25107 ;
    wire new_AGEMA_signal_25108 ;
    wire new_AGEMA_signal_25109 ;
    wire new_AGEMA_signal_25110 ;
    wire new_AGEMA_signal_25111 ;
    wire new_AGEMA_signal_25112 ;
    wire new_AGEMA_signal_25113 ;
    wire new_AGEMA_signal_25114 ;
    wire new_AGEMA_signal_25115 ;
    wire new_AGEMA_signal_25116 ;
    wire new_AGEMA_signal_25117 ;
    wire new_AGEMA_signal_25118 ;
    wire new_AGEMA_signal_25119 ;
    wire new_AGEMA_signal_25120 ;
    wire new_AGEMA_signal_25121 ;
    wire new_AGEMA_signal_25122 ;
    wire new_AGEMA_signal_25123 ;
    wire new_AGEMA_signal_25124 ;
    wire new_AGEMA_signal_25125 ;
    wire new_AGEMA_signal_25126 ;
    wire new_AGEMA_signal_25127 ;
    wire new_AGEMA_signal_25128 ;
    wire new_AGEMA_signal_25129 ;
    wire new_AGEMA_signal_25130 ;
    wire new_AGEMA_signal_25131 ;
    wire new_AGEMA_signal_25132 ;
    wire new_AGEMA_signal_25133 ;
    wire new_AGEMA_signal_25134 ;
    wire new_AGEMA_signal_25135 ;
    wire new_AGEMA_signal_25136 ;
    wire new_AGEMA_signal_25137 ;
    wire new_AGEMA_signal_25138 ;
    wire new_AGEMA_signal_25139 ;
    wire new_AGEMA_signal_25140 ;
    wire new_AGEMA_signal_25141 ;
    wire new_AGEMA_signal_25142 ;
    wire new_AGEMA_signal_25143 ;
    wire new_AGEMA_signal_25144 ;
    wire new_AGEMA_signal_25145 ;
    wire new_AGEMA_signal_25146 ;
    wire new_AGEMA_signal_25147 ;
    wire new_AGEMA_signal_25148 ;
    wire new_AGEMA_signal_25149 ;
    wire new_AGEMA_signal_25150 ;
    wire new_AGEMA_signal_25151 ;
    wire new_AGEMA_signal_25152 ;
    wire new_AGEMA_signal_25153 ;
    wire new_AGEMA_signal_25154 ;
    wire new_AGEMA_signal_25155 ;
    wire new_AGEMA_signal_25156 ;
    wire new_AGEMA_signal_25157 ;
    wire new_AGEMA_signal_25158 ;
    wire new_AGEMA_signal_25159 ;
    wire new_AGEMA_signal_25160 ;
    wire new_AGEMA_signal_25161 ;
    wire new_AGEMA_signal_25162 ;
    wire new_AGEMA_signal_25163 ;
    wire new_AGEMA_signal_25164 ;
    wire new_AGEMA_signal_25165 ;
    wire new_AGEMA_signal_25166 ;
    wire new_AGEMA_signal_25167 ;
    wire new_AGEMA_signal_25168 ;
    wire new_AGEMA_signal_25169 ;
    wire new_AGEMA_signal_25170 ;
    wire new_AGEMA_signal_25171 ;
    wire new_AGEMA_signal_25172 ;
    wire new_AGEMA_signal_25173 ;
    wire new_AGEMA_signal_25174 ;
    wire new_AGEMA_signal_25175 ;
    wire new_AGEMA_signal_25176 ;
    wire new_AGEMA_signal_25177 ;
    wire new_AGEMA_signal_25178 ;
    wire new_AGEMA_signal_25179 ;
    wire new_AGEMA_signal_25180 ;
    wire new_AGEMA_signal_25181 ;
    wire new_AGEMA_signal_25182 ;
    wire new_AGEMA_signal_25183 ;
    wire new_AGEMA_signal_25184 ;
    wire new_AGEMA_signal_25185 ;
    wire new_AGEMA_signal_25186 ;
    wire new_AGEMA_signal_25187 ;
    wire new_AGEMA_signal_25188 ;
    wire new_AGEMA_signal_25189 ;
    wire new_AGEMA_signal_25190 ;
    wire new_AGEMA_signal_25191 ;
    wire new_AGEMA_signal_25192 ;
    wire new_AGEMA_signal_25193 ;
    wire new_AGEMA_signal_25194 ;
    wire new_AGEMA_signal_25195 ;
    wire new_AGEMA_signal_25196 ;
    wire new_AGEMA_signal_25197 ;
    wire new_AGEMA_signal_25198 ;
    wire new_AGEMA_signal_25199 ;
    wire new_AGEMA_signal_25200 ;
    wire new_AGEMA_signal_25201 ;
    wire new_AGEMA_signal_25202 ;
    wire new_AGEMA_signal_25203 ;
    wire new_AGEMA_signal_25204 ;
    wire new_AGEMA_signal_25205 ;
    wire new_AGEMA_signal_25206 ;
    wire new_AGEMA_signal_25207 ;
    wire new_AGEMA_signal_25208 ;
    wire new_AGEMA_signal_25209 ;
    wire new_AGEMA_signal_25210 ;
    wire new_AGEMA_signal_25211 ;
    wire new_AGEMA_signal_25212 ;
    wire new_AGEMA_signal_25213 ;
    wire new_AGEMA_signal_25214 ;
    wire new_AGEMA_signal_25215 ;
    wire new_AGEMA_signal_25216 ;
    wire new_AGEMA_signal_25217 ;
    wire new_AGEMA_signal_25218 ;
    wire new_AGEMA_signal_25219 ;
    wire new_AGEMA_signal_25220 ;
    wire new_AGEMA_signal_25221 ;
    wire new_AGEMA_signal_25222 ;
    wire new_AGEMA_signal_25223 ;
    wire new_AGEMA_signal_25224 ;
    wire new_AGEMA_signal_25225 ;
    wire new_AGEMA_signal_25226 ;
    wire new_AGEMA_signal_25227 ;
    wire new_AGEMA_signal_25228 ;
    wire new_AGEMA_signal_25229 ;
    wire new_AGEMA_signal_25230 ;
    wire new_AGEMA_signal_25231 ;
    wire new_AGEMA_signal_25232 ;
    wire new_AGEMA_signal_25233 ;
    wire new_AGEMA_signal_25234 ;
    wire new_AGEMA_signal_25235 ;
    wire new_AGEMA_signal_25236 ;
    wire new_AGEMA_signal_25237 ;
    wire new_AGEMA_signal_25238 ;
    wire new_AGEMA_signal_25239 ;
    wire new_AGEMA_signal_25240 ;
    wire new_AGEMA_signal_25241 ;
    wire new_AGEMA_signal_25242 ;
    wire new_AGEMA_signal_25243 ;
    wire new_AGEMA_signal_25244 ;
    wire new_AGEMA_signal_25245 ;
    wire new_AGEMA_signal_25246 ;
    wire new_AGEMA_signal_25247 ;
    wire new_AGEMA_signal_25248 ;
    wire new_AGEMA_signal_25249 ;
    wire new_AGEMA_signal_25250 ;
    wire new_AGEMA_signal_25251 ;
    wire new_AGEMA_signal_25252 ;
    wire new_AGEMA_signal_25253 ;
    wire new_AGEMA_signal_25254 ;
    wire new_AGEMA_signal_25255 ;
    wire new_AGEMA_signal_25256 ;
    wire new_AGEMA_signal_25257 ;
    wire new_AGEMA_signal_25258 ;
    wire new_AGEMA_signal_25259 ;
    wire new_AGEMA_signal_25260 ;
    wire new_AGEMA_signal_25261 ;
    wire new_AGEMA_signal_25262 ;
    wire new_AGEMA_signal_25263 ;
    wire new_AGEMA_signal_25264 ;
    wire new_AGEMA_signal_25265 ;
    wire new_AGEMA_signal_25266 ;
    wire new_AGEMA_signal_25267 ;
    wire new_AGEMA_signal_25268 ;
    wire new_AGEMA_signal_25269 ;
    wire new_AGEMA_signal_25270 ;
    wire new_AGEMA_signal_25271 ;
    wire new_AGEMA_signal_25272 ;
    wire new_AGEMA_signal_25273 ;
    wire new_AGEMA_signal_25274 ;
    wire new_AGEMA_signal_25275 ;
    wire new_AGEMA_signal_25276 ;
    wire new_AGEMA_signal_25277 ;
    wire new_AGEMA_signal_25278 ;
    wire new_AGEMA_signal_25279 ;
    wire new_AGEMA_signal_25280 ;
    wire new_AGEMA_signal_25281 ;
    wire new_AGEMA_signal_25282 ;
    wire new_AGEMA_signal_25283 ;
    wire new_AGEMA_signal_25284 ;
    wire new_AGEMA_signal_25285 ;
    wire new_AGEMA_signal_25286 ;
    wire new_AGEMA_signal_25287 ;
    wire new_AGEMA_signal_25288 ;
    wire new_AGEMA_signal_25289 ;
    wire new_AGEMA_signal_25290 ;
    wire new_AGEMA_signal_25291 ;
    wire new_AGEMA_signal_25292 ;
    wire new_AGEMA_signal_25293 ;
    wire new_AGEMA_signal_25294 ;
    wire new_AGEMA_signal_25295 ;
    wire new_AGEMA_signal_25296 ;
    wire new_AGEMA_signal_25297 ;
    wire new_AGEMA_signal_25298 ;
    wire new_AGEMA_signal_25299 ;
    wire new_AGEMA_signal_25300 ;
    wire new_AGEMA_signal_25301 ;
    wire new_AGEMA_signal_25302 ;
    wire new_AGEMA_signal_25303 ;
    wire new_AGEMA_signal_25304 ;
    wire new_AGEMA_signal_25305 ;
    wire new_AGEMA_signal_25306 ;
    wire new_AGEMA_signal_25307 ;
    wire new_AGEMA_signal_25308 ;
    wire new_AGEMA_signal_25309 ;
    wire new_AGEMA_signal_25310 ;
    wire new_AGEMA_signal_25311 ;
    wire new_AGEMA_signal_25312 ;
    wire new_AGEMA_signal_25313 ;
    wire new_AGEMA_signal_25314 ;
    wire new_AGEMA_signal_25315 ;
    wire new_AGEMA_signal_25316 ;
    wire new_AGEMA_signal_25317 ;
    wire new_AGEMA_signal_25318 ;
    wire new_AGEMA_signal_25319 ;
    wire new_AGEMA_signal_25320 ;
    wire new_AGEMA_signal_25321 ;
    wire new_AGEMA_signal_25322 ;
    wire new_AGEMA_signal_25323 ;
    wire new_AGEMA_signal_25324 ;
    wire new_AGEMA_signal_25325 ;
    wire new_AGEMA_signal_25326 ;
    wire new_AGEMA_signal_25327 ;
    wire new_AGEMA_signal_25328 ;
    wire new_AGEMA_signal_25329 ;
    wire new_AGEMA_signal_25330 ;
    wire new_AGEMA_signal_25331 ;
    wire new_AGEMA_signal_25332 ;
    wire new_AGEMA_signal_25333 ;
    wire new_AGEMA_signal_25334 ;
    wire new_AGEMA_signal_25335 ;
    wire new_AGEMA_signal_25336 ;
    wire new_AGEMA_signal_25337 ;
    wire new_AGEMA_signal_25338 ;
    wire new_AGEMA_signal_25339 ;
    wire new_AGEMA_signal_25340 ;
    wire new_AGEMA_signal_25341 ;
    wire new_AGEMA_signal_25342 ;
    wire new_AGEMA_signal_25343 ;
    wire new_AGEMA_signal_25344 ;
    wire new_AGEMA_signal_25345 ;
    wire new_AGEMA_signal_25346 ;
    wire new_AGEMA_signal_25347 ;
    wire new_AGEMA_signal_25348 ;
    wire new_AGEMA_signal_25349 ;
    wire new_AGEMA_signal_25350 ;
    wire new_AGEMA_signal_25351 ;
    wire new_AGEMA_signal_25352 ;
    wire new_AGEMA_signal_25353 ;
    wire new_AGEMA_signal_25354 ;
    wire new_AGEMA_signal_25355 ;
    wire new_AGEMA_signal_25356 ;
    wire new_AGEMA_signal_25357 ;
    wire new_AGEMA_signal_25358 ;
    wire new_AGEMA_signal_25359 ;
    wire new_AGEMA_signal_25360 ;
    wire new_AGEMA_signal_25361 ;
    wire new_AGEMA_signal_25362 ;
    wire new_AGEMA_signal_25363 ;
    wire new_AGEMA_signal_25364 ;
    wire new_AGEMA_signal_25365 ;
    wire new_AGEMA_signal_25366 ;
    wire new_AGEMA_signal_25367 ;
    wire new_AGEMA_signal_25368 ;
    wire new_AGEMA_signal_25369 ;
    wire new_AGEMA_signal_25370 ;
    wire new_AGEMA_signal_25371 ;
    wire new_AGEMA_signal_25372 ;
    wire new_AGEMA_signal_25373 ;
    wire new_AGEMA_signal_25374 ;
    wire new_AGEMA_signal_25375 ;
    wire new_AGEMA_signal_25376 ;
    wire new_AGEMA_signal_25377 ;
    wire new_AGEMA_signal_25378 ;
    wire new_AGEMA_signal_25379 ;
    wire new_AGEMA_signal_25380 ;
    wire new_AGEMA_signal_25381 ;
    wire new_AGEMA_signal_25382 ;
    wire new_AGEMA_signal_25383 ;
    wire new_AGEMA_signal_25384 ;
    wire new_AGEMA_signal_25385 ;
    wire new_AGEMA_signal_25386 ;
    wire new_AGEMA_signal_25387 ;
    wire new_AGEMA_signal_25388 ;
    wire new_AGEMA_signal_25389 ;
    wire new_AGEMA_signal_25390 ;
    wire new_AGEMA_signal_25391 ;
    wire new_AGEMA_signal_25392 ;
    wire new_AGEMA_signal_25393 ;
    wire new_AGEMA_signal_25394 ;
    wire new_AGEMA_signal_25395 ;
    wire new_AGEMA_signal_25396 ;
    wire new_AGEMA_signal_25397 ;
    wire new_AGEMA_signal_25398 ;
    wire new_AGEMA_signal_25399 ;
    wire new_AGEMA_signal_25400 ;
    wire new_AGEMA_signal_25401 ;
    wire new_AGEMA_signal_25402 ;
    wire new_AGEMA_signal_25403 ;
    wire new_AGEMA_signal_25404 ;
    wire new_AGEMA_signal_25405 ;
    wire new_AGEMA_signal_25406 ;
    wire new_AGEMA_signal_25407 ;
    wire new_AGEMA_signal_25408 ;
    wire new_AGEMA_signal_25409 ;
    wire new_AGEMA_signal_25410 ;
    wire new_AGEMA_signal_25411 ;
    wire new_AGEMA_signal_25412 ;
    wire new_AGEMA_signal_25413 ;
    wire new_AGEMA_signal_25414 ;
    wire new_AGEMA_signal_25415 ;
    wire new_AGEMA_signal_25416 ;
    wire new_AGEMA_signal_25417 ;
    wire new_AGEMA_signal_25418 ;
    wire new_AGEMA_signal_25419 ;
    wire new_AGEMA_signal_25420 ;
    wire new_AGEMA_signal_25421 ;
    wire new_AGEMA_signal_25422 ;
    wire new_AGEMA_signal_25423 ;
    wire new_AGEMA_signal_25424 ;
    wire new_AGEMA_signal_25425 ;
    wire new_AGEMA_signal_25426 ;
    wire new_AGEMA_signal_25427 ;
    wire new_AGEMA_signal_25428 ;
    wire new_AGEMA_signal_25429 ;
    wire new_AGEMA_signal_25430 ;
    wire new_AGEMA_signal_25431 ;
    wire new_AGEMA_signal_25432 ;
    wire new_AGEMA_signal_25433 ;
    wire new_AGEMA_signal_25434 ;
    wire new_AGEMA_signal_25435 ;
    wire new_AGEMA_signal_25436 ;
    wire new_AGEMA_signal_25437 ;
    wire new_AGEMA_signal_25438 ;
    wire new_AGEMA_signal_25439 ;
    wire new_AGEMA_signal_25440 ;
    wire new_AGEMA_signal_25441 ;
    wire new_AGEMA_signal_25442 ;
    wire new_AGEMA_signal_25443 ;
    wire new_AGEMA_signal_25444 ;
    wire new_AGEMA_signal_25445 ;
    wire new_AGEMA_signal_25446 ;
    wire new_AGEMA_signal_25447 ;
    wire new_AGEMA_signal_25448 ;
    wire new_AGEMA_signal_25449 ;
    wire new_AGEMA_signal_25450 ;
    wire new_AGEMA_signal_25451 ;
    wire new_AGEMA_signal_25452 ;
    wire new_AGEMA_signal_25453 ;
    wire new_AGEMA_signal_25454 ;
    wire new_AGEMA_signal_25455 ;
    wire new_AGEMA_signal_25456 ;
    wire new_AGEMA_signal_25457 ;
    wire new_AGEMA_signal_25458 ;
    wire new_AGEMA_signal_25459 ;
    wire new_AGEMA_signal_25460 ;
    wire new_AGEMA_signal_25461 ;
    wire new_AGEMA_signal_25462 ;
    wire new_AGEMA_signal_25463 ;
    wire new_AGEMA_signal_25464 ;
    wire new_AGEMA_signal_25465 ;
    wire new_AGEMA_signal_25466 ;
    wire new_AGEMA_signal_25467 ;
    wire new_AGEMA_signal_25468 ;
    wire new_AGEMA_signal_25469 ;
    wire new_AGEMA_signal_25470 ;
    wire new_AGEMA_signal_25471 ;
    wire new_AGEMA_signal_25472 ;
    wire new_AGEMA_signal_25473 ;
    wire new_AGEMA_signal_25474 ;
    wire new_AGEMA_signal_25475 ;
    wire new_AGEMA_signal_25476 ;
    wire new_AGEMA_signal_25477 ;
    wire new_AGEMA_signal_25478 ;
    wire new_AGEMA_signal_25479 ;
    wire new_AGEMA_signal_25480 ;
    wire new_AGEMA_signal_25481 ;
    wire new_AGEMA_signal_25482 ;
    wire new_AGEMA_signal_25483 ;
    wire new_AGEMA_signal_25484 ;
    wire new_AGEMA_signal_25485 ;
    wire new_AGEMA_signal_25486 ;
    wire new_AGEMA_signal_25487 ;
    wire new_AGEMA_signal_25488 ;
    wire new_AGEMA_signal_25489 ;
    wire new_AGEMA_signal_25490 ;
    wire new_AGEMA_signal_25491 ;
    wire new_AGEMA_signal_25492 ;
    wire new_AGEMA_signal_25493 ;
    wire new_AGEMA_signal_25494 ;
    wire new_AGEMA_signal_25495 ;
    wire new_AGEMA_signal_25496 ;
    wire new_AGEMA_signal_25497 ;
    wire new_AGEMA_signal_25498 ;
    wire new_AGEMA_signal_25499 ;
    wire new_AGEMA_signal_25500 ;
    wire new_AGEMA_signal_25501 ;
    wire new_AGEMA_signal_25502 ;
    wire new_AGEMA_signal_25503 ;
    wire new_AGEMA_signal_25504 ;
    wire new_AGEMA_signal_25505 ;
    wire new_AGEMA_signal_25506 ;
    wire new_AGEMA_signal_25507 ;
    wire new_AGEMA_signal_25508 ;
    wire new_AGEMA_signal_25509 ;
    wire new_AGEMA_signal_25510 ;
    wire new_AGEMA_signal_25511 ;
    wire new_AGEMA_signal_25512 ;
    wire new_AGEMA_signal_25513 ;
    wire new_AGEMA_signal_25514 ;
    wire new_AGEMA_signal_25515 ;
    wire new_AGEMA_signal_25516 ;
    wire new_AGEMA_signal_25517 ;
    wire new_AGEMA_signal_25518 ;
    wire new_AGEMA_signal_25519 ;
    wire new_AGEMA_signal_25520 ;
    wire new_AGEMA_signal_25521 ;
    wire new_AGEMA_signal_25522 ;
    wire new_AGEMA_signal_25523 ;
    wire new_AGEMA_signal_25524 ;
    wire new_AGEMA_signal_25525 ;
    wire new_AGEMA_signal_25526 ;
    wire new_AGEMA_signal_25527 ;
    wire new_AGEMA_signal_25528 ;
    wire new_AGEMA_signal_25529 ;
    wire new_AGEMA_signal_25530 ;
    wire new_AGEMA_signal_25531 ;
    wire new_AGEMA_signal_25532 ;
    wire new_AGEMA_signal_25533 ;
    wire new_AGEMA_signal_25534 ;
    wire new_AGEMA_signal_25535 ;
    wire new_AGEMA_signal_25536 ;
    wire new_AGEMA_signal_25537 ;
    wire new_AGEMA_signal_25538 ;
    wire new_AGEMA_signal_25539 ;
    wire new_AGEMA_signal_25540 ;
    wire new_AGEMA_signal_25541 ;
    wire new_AGEMA_signal_25542 ;
    wire new_AGEMA_signal_25543 ;
    wire new_AGEMA_signal_25544 ;
    wire new_AGEMA_signal_25545 ;
    wire new_AGEMA_signal_25546 ;
    wire new_AGEMA_signal_25547 ;
    wire new_AGEMA_signal_25548 ;
    wire new_AGEMA_signal_25549 ;
    wire new_AGEMA_signal_25550 ;
    wire new_AGEMA_signal_25551 ;
    wire new_AGEMA_signal_25552 ;
    wire new_AGEMA_signal_25553 ;
    wire new_AGEMA_signal_25554 ;
    wire new_AGEMA_signal_25555 ;
    wire new_AGEMA_signal_25556 ;
    wire new_AGEMA_signal_25557 ;
    wire new_AGEMA_signal_25558 ;
    wire new_AGEMA_signal_25559 ;
    wire new_AGEMA_signal_25560 ;
    wire new_AGEMA_signal_25561 ;
    wire new_AGEMA_signal_25562 ;
    wire new_AGEMA_signal_25563 ;
    wire new_AGEMA_signal_25564 ;
    wire new_AGEMA_signal_25565 ;
    wire new_AGEMA_signal_25566 ;
    wire new_AGEMA_signal_25567 ;
    wire new_AGEMA_signal_25568 ;
    wire new_AGEMA_signal_25569 ;
    wire new_AGEMA_signal_25570 ;
    wire new_AGEMA_signal_25571 ;
    wire new_AGEMA_signal_25572 ;
    wire new_AGEMA_signal_25573 ;
    wire new_AGEMA_signal_25574 ;
    wire new_AGEMA_signal_25575 ;
    wire new_AGEMA_signal_25576 ;
    wire new_AGEMA_signal_25577 ;
    wire new_AGEMA_signal_25578 ;
    wire new_AGEMA_signal_25579 ;
    wire new_AGEMA_signal_25580 ;
    wire new_AGEMA_signal_25581 ;
    wire new_AGEMA_signal_25582 ;
    wire new_AGEMA_signal_25583 ;
    wire new_AGEMA_signal_25584 ;
    wire new_AGEMA_signal_25585 ;
    wire new_AGEMA_signal_25586 ;
    wire new_AGEMA_signal_25587 ;
    wire new_AGEMA_signal_25588 ;
    wire new_AGEMA_signal_25589 ;
    wire new_AGEMA_signal_25590 ;
    wire new_AGEMA_signal_25591 ;
    wire new_AGEMA_signal_25592 ;
    wire new_AGEMA_signal_25593 ;
    wire new_AGEMA_signal_25594 ;
    wire new_AGEMA_signal_25595 ;
    wire new_AGEMA_signal_25596 ;
    wire new_AGEMA_signal_25597 ;
    wire new_AGEMA_signal_25598 ;
    wire new_AGEMA_signal_25599 ;
    wire new_AGEMA_signal_25600 ;
    wire new_AGEMA_signal_25601 ;
    wire new_AGEMA_signal_25602 ;
    wire new_AGEMA_signal_25603 ;
    wire new_AGEMA_signal_25604 ;
    wire new_AGEMA_signal_25605 ;
    wire new_AGEMA_signal_25606 ;
    wire new_AGEMA_signal_25607 ;
    wire new_AGEMA_signal_25608 ;
    wire new_AGEMA_signal_25609 ;
    wire new_AGEMA_signal_25610 ;
    wire new_AGEMA_signal_25611 ;
    wire new_AGEMA_signal_25612 ;
    wire new_AGEMA_signal_25613 ;
    wire new_AGEMA_signal_25614 ;
    wire new_AGEMA_signal_25615 ;
    wire new_AGEMA_signal_25616 ;
    wire new_AGEMA_signal_25617 ;
    wire new_AGEMA_signal_25618 ;
    wire new_AGEMA_signal_25619 ;
    wire new_AGEMA_signal_25620 ;
    wire new_AGEMA_signal_25621 ;
    wire new_AGEMA_signal_25622 ;
    wire new_AGEMA_signal_25623 ;
    wire new_AGEMA_signal_25624 ;
    wire new_AGEMA_signal_25625 ;
    wire new_AGEMA_signal_25626 ;
    wire new_AGEMA_signal_25627 ;
    wire new_AGEMA_signal_25628 ;
    wire new_AGEMA_signal_25629 ;
    wire new_AGEMA_signal_25630 ;
    wire new_AGEMA_signal_25631 ;
    wire new_AGEMA_signal_25632 ;
    wire new_AGEMA_signal_25633 ;
    wire new_AGEMA_signal_25634 ;
    wire new_AGEMA_signal_25635 ;
    wire new_AGEMA_signal_25636 ;
    wire new_AGEMA_signal_25637 ;
    wire new_AGEMA_signal_25638 ;
    wire new_AGEMA_signal_25639 ;
    wire new_AGEMA_signal_25640 ;
    wire new_AGEMA_signal_25641 ;
    wire new_AGEMA_signal_25642 ;
    wire new_AGEMA_signal_25643 ;
    wire new_AGEMA_signal_25644 ;
    wire new_AGEMA_signal_25645 ;
    wire new_AGEMA_signal_25646 ;
    wire new_AGEMA_signal_25647 ;
    wire new_AGEMA_signal_25648 ;
    wire new_AGEMA_signal_25649 ;
    wire new_AGEMA_signal_25650 ;
    wire new_AGEMA_signal_25651 ;
    wire new_AGEMA_signal_25652 ;
    wire new_AGEMA_signal_25653 ;
    wire new_AGEMA_signal_25654 ;
    wire new_AGEMA_signal_25655 ;
    wire new_AGEMA_signal_25656 ;
    wire new_AGEMA_signal_25657 ;
    wire new_AGEMA_signal_25658 ;
    wire new_AGEMA_signal_25659 ;
    wire new_AGEMA_signal_25660 ;
    wire new_AGEMA_signal_25661 ;
    wire new_AGEMA_signal_25662 ;
    wire new_AGEMA_signal_25663 ;
    wire new_AGEMA_signal_25664 ;
    wire new_AGEMA_signal_25665 ;
    wire new_AGEMA_signal_25666 ;
    wire new_AGEMA_signal_25667 ;
    wire new_AGEMA_signal_25668 ;
    wire new_AGEMA_signal_25669 ;
    wire new_AGEMA_signal_25670 ;
    wire new_AGEMA_signal_25671 ;
    wire new_AGEMA_signal_25672 ;
    wire new_AGEMA_signal_25673 ;
    wire new_AGEMA_signal_25674 ;
    wire new_AGEMA_signal_25675 ;
    wire new_AGEMA_signal_25676 ;
    wire new_AGEMA_signal_25677 ;
    wire new_AGEMA_signal_25678 ;
    wire new_AGEMA_signal_25679 ;
    wire new_AGEMA_signal_25680 ;
    wire new_AGEMA_signal_25681 ;
    wire new_AGEMA_signal_25682 ;
    wire new_AGEMA_signal_25683 ;
    wire new_AGEMA_signal_25684 ;
    wire new_AGEMA_signal_25685 ;
    wire new_AGEMA_signal_25686 ;
    wire new_AGEMA_signal_25687 ;
    wire new_AGEMA_signal_25688 ;
    wire new_AGEMA_signal_25689 ;
    wire new_AGEMA_signal_25690 ;
    wire new_AGEMA_signal_25691 ;
    wire new_AGEMA_signal_25692 ;
    wire new_AGEMA_signal_25693 ;
    wire new_AGEMA_signal_25694 ;
    wire new_AGEMA_signal_25695 ;
    wire new_AGEMA_signal_25696 ;
    wire new_AGEMA_signal_25697 ;
    wire new_AGEMA_signal_25698 ;
    wire new_AGEMA_signal_25699 ;
    wire new_AGEMA_signal_25700 ;
    wire new_AGEMA_signal_25701 ;
    wire new_AGEMA_signal_25702 ;
    wire new_AGEMA_signal_25703 ;
    wire new_AGEMA_signal_25704 ;
    wire new_AGEMA_signal_25705 ;
    wire new_AGEMA_signal_25706 ;
    wire new_AGEMA_signal_25707 ;
    wire new_AGEMA_signal_25708 ;
    wire new_AGEMA_signal_25709 ;
    wire new_AGEMA_signal_25710 ;
    wire new_AGEMA_signal_25711 ;
    wire new_AGEMA_signal_25712 ;
    wire new_AGEMA_signal_25713 ;
    wire new_AGEMA_signal_25714 ;
    wire new_AGEMA_signal_25715 ;
    wire new_AGEMA_signal_25716 ;
    wire new_AGEMA_signal_25717 ;
    wire new_AGEMA_signal_25718 ;
    wire new_AGEMA_signal_25719 ;
    wire new_AGEMA_signal_25720 ;
    wire new_AGEMA_signal_25721 ;
    wire new_AGEMA_signal_25722 ;
    wire new_AGEMA_signal_25723 ;
    wire new_AGEMA_signal_25724 ;
    wire new_AGEMA_signal_25725 ;
    wire new_AGEMA_signal_25726 ;
    wire new_AGEMA_signal_25727 ;
    wire new_AGEMA_signal_25728 ;
    wire new_AGEMA_signal_25729 ;
    wire new_AGEMA_signal_25730 ;
    wire new_AGEMA_signal_25731 ;
    wire new_AGEMA_signal_25732 ;
    wire new_AGEMA_signal_25733 ;
    wire new_AGEMA_signal_25734 ;
    wire new_AGEMA_signal_25735 ;
    wire new_AGEMA_signal_25736 ;
    wire new_AGEMA_signal_25737 ;
    wire new_AGEMA_signal_25738 ;
    wire new_AGEMA_signal_25739 ;
    wire new_AGEMA_signal_25740 ;
    wire new_AGEMA_signal_25741 ;
    wire new_AGEMA_signal_25742 ;
    wire new_AGEMA_signal_25743 ;
    wire new_AGEMA_signal_25744 ;
    wire new_AGEMA_signal_25745 ;
    wire new_AGEMA_signal_25746 ;
    wire new_AGEMA_signal_25747 ;
    wire new_AGEMA_signal_25748 ;
    wire new_AGEMA_signal_25749 ;
    wire new_AGEMA_signal_25750 ;
    wire new_AGEMA_signal_25751 ;
    wire new_AGEMA_signal_25752 ;
    wire new_AGEMA_signal_25753 ;
    wire new_AGEMA_signal_25754 ;
    wire new_AGEMA_signal_25755 ;
    wire new_AGEMA_signal_25756 ;
    wire new_AGEMA_signal_25757 ;
    wire new_AGEMA_signal_25758 ;
    wire new_AGEMA_signal_25759 ;
    wire new_AGEMA_signal_25760 ;
    wire new_AGEMA_signal_25761 ;
    wire new_AGEMA_signal_25762 ;
    wire new_AGEMA_signal_25763 ;
    wire new_AGEMA_signal_25764 ;
    wire new_AGEMA_signal_25765 ;
    wire new_AGEMA_signal_25766 ;
    wire new_AGEMA_signal_25767 ;
    wire new_AGEMA_signal_25768 ;
    wire new_AGEMA_signal_25769 ;
    wire new_AGEMA_signal_25770 ;
    wire new_AGEMA_signal_25771 ;
    wire new_AGEMA_signal_25772 ;
    wire new_AGEMA_signal_25773 ;
    wire new_AGEMA_signal_25774 ;
    wire new_AGEMA_signal_25775 ;
    wire new_AGEMA_signal_25776 ;
    wire new_AGEMA_signal_25777 ;
    wire new_AGEMA_signal_25778 ;
    wire new_AGEMA_signal_25779 ;
    wire new_AGEMA_signal_25780 ;
    wire new_AGEMA_signal_25781 ;
    wire new_AGEMA_signal_25782 ;
    wire new_AGEMA_signal_25783 ;
    wire new_AGEMA_signal_25784 ;
    wire new_AGEMA_signal_25785 ;
    wire new_AGEMA_signal_25786 ;
    wire new_AGEMA_signal_25787 ;
    wire new_AGEMA_signal_25788 ;
    wire new_AGEMA_signal_25789 ;
    wire new_AGEMA_signal_25790 ;
    wire new_AGEMA_signal_25791 ;
    wire new_AGEMA_signal_25792 ;
    wire new_AGEMA_signal_25793 ;
    wire new_AGEMA_signal_25794 ;
    wire new_AGEMA_signal_25795 ;
    wire new_AGEMA_signal_25796 ;
    wire new_AGEMA_signal_25797 ;
    wire new_AGEMA_signal_25798 ;
    wire new_AGEMA_signal_25799 ;
    wire new_AGEMA_signal_25800 ;
    wire new_AGEMA_signal_25801 ;
    wire new_AGEMA_signal_25802 ;
    wire new_AGEMA_signal_25803 ;
    wire new_AGEMA_signal_25804 ;
    wire new_AGEMA_signal_25805 ;
    wire new_AGEMA_signal_25806 ;
    wire new_AGEMA_signal_25807 ;
    wire new_AGEMA_signal_25808 ;
    wire new_AGEMA_signal_25809 ;
    wire new_AGEMA_signal_25810 ;
    wire new_AGEMA_signal_25811 ;
    wire new_AGEMA_signal_25812 ;
    wire new_AGEMA_signal_25813 ;
    wire new_AGEMA_signal_25814 ;
    wire new_AGEMA_signal_25815 ;
    wire new_AGEMA_signal_25816 ;
    wire new_AGEMA_signal_25817 ;
    wire new_AGEMA_signal_25818 ;
    wire new_AGEMA_signal_25819 ;
    wire new_AGEMA_signal_25820 ;
    wire new_AGEMA_signal_25821 ;
    wire new_AGEMA_signal_25822 ;
    wire new_AGEMA_signal_25823 ;
    wire new_AGEMA_signal_25824 ;
    wire new_AGEMA_signal_25825 ;
    wire new_AGEMA_signal_25826 ;
    wire new_AGEMA_signal_25827 ;
    wire new_AGEMA_signal_25828 ;
    wire new_AGEMA_signal_25829 ;
    wire new_AGEMA_signal_25830 ;
    wire new_AGEMA_signal_25831 ;
    wire new_AGEMA_signal_25832 ;
    wire new_AGEMA_signal_25833 ;
    wire new_AGEMA_signal_25834 ;
    wire new_AGEMA_signal_25835 ;
    wire new_AGEMA_signal_25836 ;
    wire new_AGEMA_signal_25837 ;
    wire new_AGEMA_signal_25838 ;
    wire new_AGEMA_signal_25839 ;
    wire new_AGEMA_signal_25840 ;
    wire new_AGEMA_signal_25841 ;
    wire new_AGEMA_signal_25842 ;
    wire new_AGEMA_signal_25843 ;
    wire new_AGEMA_signal_25844 ;
    wire new_AGEMA_signal_25845 ;
    wire new_AGEMA_signal_25846 ;
    wire new_AGEMA_signal_25847 ;
    wire new_AGEMA_signal_25848 ;
    wire new_AGEMA_signal_25849 ;
    wire new_AGEMA_signal_25850 ;
    wire new_AGEMA_signal_25851 ;
    wire new_AGEMA_signal_25852 ;
    wire new_AGEMA_signal_25853 ;
    wire new_AGEMA_signal_25854 ;
    wire new_AGEMA_signal_25855 ;
    wire new_AGEMA_signal_25856 ;
    wire new_AGEMA_signal_25857 ;
    wire new_AGEMA_signal_25858 ;
    wire new_AGEMA_signal_25859 ;
    wire new_AGEMA_signal_25860 ;
    wire new_AGEMA_signal_25861 ;
    wire new_AGEMA_signal_25862 ;
    wire new_AGEMA_signal_25863 ;
    wire new_AGEMA_signal_25864 ;
    wire new_AGEMA_signal_25865 ;
    wire new_AGEMA_signal_25866 ;
    wire new_AGEMA_signal_25867 ;
    wire new_AGEMA_signal_25868 ;
    wire new_AGEMA_signal_25869 ;
    wire new_AGEMA_signal_25870 ;
    wire new_AGEMA_signal_25871 ;
    wire new_AGEMA_signal_25872 ;
    wire new_AGEMA_signal_25873 ;
    wire new_AGEMA_signal_25874 ;
    wire new_AGEMA_signal_25875 ;
    wire new_AGEMA_signal_25876 ;
    wire new_AGEMA_signal_25877 ;
    wire new_AGEMA_signal_25878 ;
    wire new_AGEMA_signal_25879 ;
    wire new_AGEMA_signal_25880 ;
    wire new_AGEMA_signal_25881 ;
    wire new_AGEMA_signal_25882 ;
    wire new_AGEMA_signal_25883 ;
    wire new_AGEMA_signal_25884 ;
    wire new_AGEMA_signal_25885 ;
    wire new_AGEMA_signal_25886 ;
    wire new_AGEMA_signal_25887 ;
    wire new_AGEMA_signal_25888 ;
    wire new_AGEMA_signal_25889 ;
    wire new_AGEMA_signal_25890 ;
    wire new_AGEMA_signal_25891 ;
    wire new_AGEMA_signal_25892 ;
    wire new_AGEMA_signal_25893 ;
    wire new_AGEMA_signal_25894 ;
    wire new_AGEMA_signal_25895 ;
    wire new_AGEMA_signal_25896 ;
    wire new_AGEMA_signal_25897 ;
    wire new_AGEMA_signal_25898 ;
    wire new_AGEMA_signal_25899 ;
    wire new_AGEMA_signal_25900 ;
    wire new_AGEMA_signal_25901 ;
    wire new_AGEMA_signal_25902 ;
    wire new_AGEMA_signal_25903 ;
    wire new_AGEMA_signal_25904 ;
    wire new_AGEMA_signal_25905 ;
    wire new_AGEMA_signal_25906 ;
    wire new_AGEMA_signal_25907 ;
    wire new_AGEMA_signal_25908 ;
    wire new_AGEMA_signal_25909 ;
    wire new_AGEMA_signal_25910 ;
    wire new_AGEMA_signal_25911 ;
    wire new_AGEMA_signal_25912 ;
    wire new_AGEMA_signal_25913 ;
    wire new_AGEMA_signal_25914 ;
    wire new_AGEMA_signal_25915 ;
    wire new_AGEMA_signal_25916 ;
    wire new_AGEMA_signal_25917 ;
    wire new_AGEMA_signal_25918 ;
    wire new_AGEMA_signal_25919 ;
    wire new_AGEMA_signal_25920 ;
    wire new_AGEMA_signal_25921 ;
    wire new_AGEMA_signal_25922 ;
    wire new_AGEMA_signal_25923 ;
    wire new_AGEMA_signal_25924 ;
    wire new_AGEMA_signal_25925 ;
    wire new_AGEMA_signal_25926 ;
    wire new_AGEMA_signal_25927 ;
    wire new_AGEMA_signal_25928 ;
    wire new_AGEMA_signal_25929 ;
    wire new_AGEMA_signal_25930 ;
    wire new_AGEMA_signal_25931 ;
    wire new_AGEMA_signal_25932 ;
    wire new_AGEMA_signal_25933 ;
    wire new_AGEMA_signal_25934 ;
    wire new_AGEMA_signal_25935 ;
    wire new_AGEMA_signal_25936 ;
    wire new_AGEMA_signal_25937 ;
    wire new_AGEMA_signal_25938 ;
    wire new_AGEMA_signal_25939 ;
    wire new_AGEMA_signal_25940 ;
    wire new_AGEMA_signal_25941 ;
    wire new_AGEMA_signal_25942 ;
    wire new_AGEMA_signal_25943 ;
    wire new_AGEMA_signal_25944 ;
    wire new_AGEMA_signal_25945 ;
    wire new_AGEMA_signal_25946 ;
    wire new_AGEMA_signal_25947 ;
    wire new_AGEMA_signal_25948 ;
    wire new_AGEMA_signal_25949 ;
    wire new_AGEMA_signal_25950 ;
    wire new_AGEMA_signal_25951 ;
    wire new_AGEMA_signal_25952 ;
    wire new_AGEMA_signal_25953 ;
    wire new_AGEMA_signal_25954 ;
    wire new_AGEMA_signal_25955 ;
    wire new_AGEMA_signal_25956 ;
    wire new_AGEMA_signal_25957 ;
    wire new_AGEMA_signal_25958 ;
    wire new_AGEMA_signal_25959 ;
    wire new_AGEMA_signal_25960 ;
    wire new_AGEMA_signal_25961 ;
    wire new_AGEMA_signal_25962 ;
    wire new_AGEMA_signal_25963 ;
    wire new_AGEMA_signal_25964 ;
    wire new_AGEMA_signal_25965 ;
    wire new_AGEMA_signal_25966 ;
    wire new_AGEMA_signal_25967 ;
    wire new_AGEMA_signal_25968 ;
    wire new_AGEMA_signal_25969 ;
    wire new_AGEMA_signal_25970 ;
    wire new_AGEMA_signal_25971 ;
    wire new_AGEMA_signal_25972 ;
    wire new_AGEMA_signal_25973 ;
    wire new_AGEMA_signal_25974 ;
    wire new_AGEMA_signal_25975 ;
    wire new_AGEMA_signal_25976 ;
    wire new_AGEMA_signal_25977 ;
    wire new_AGEMA_signal_25978 ;
    wire new_AGEMA_signal_25979 ;
    wire new_AGEMA_signal_25980 ;
    wire new_AGEMA_signal_25981 ;
    wire new_AGEMA_signal_25982 ;
    wire new_AGEMA_signal_25983 ;
    wire new_AGEMA_signal_25984 ;
    wire new_AGEMA_signal_25985 ;
    wire new_AGEMA_signal_25986 ;
    wire new_AGEMA_signal_25987 ;
    wire new_AGEMA_signal_25988 ;
    wire new_AGEMA_signal_25989 ;
    wire new_AGEMA_signal_25990 ;
    wire new_AGEMA_signal_25991 ;
    wire new_AGEMA_signal_25992 ;
    wire new_AGEMA_signal_25993 ;
    wire new_AGEMA_signal_25994 ;
    wire new_AGEMA_signal_25995 ;
    wire new_AGEMA_signal_25996 ;
    wire new_AGEMA_signal_25997 ;
    wire new_AGEMA_signal_25998 ;
    wire new_AGEMA_signal_25999 ;
    wire new_AGEMA_signal_26000 ;
    wire new_AGEMA_signal_26001 ;
    wire new_AGEMA_signal_26002 ;
    wire new_AGEMA_signal_26003 ;
    wire new_AGEMA_signal_26004 ;
    wire new_AGEMA_signal_26005 ;
    wire new_AGEMA_signal_26006 ;
    wire new_AGEMA_signal_26007 ;
    wire new_AGEMA_signal_26008 ;
    wire new_AGEMA_signal_26009 ;
    wire new_AGEMA_signal_26010 ;
    wire new_AGEMA_signal_26011 ;
    wire new_AGEMA_signal_26012 ;
    wire new_AGEMA_signal_26013 ;
    wire new_AGEMA_signal_26014 ;
    wire new_AGEMA_signal_26015 ;
    wire new_AGEMA_signal_26016 ;
    wire new_AGEMA_signal_26017 ;
    wire new_AGEMA_signal_26018 ;
    wire new_AGEMA_signal_26019 ;
    wire new_AGEMA_signal_26020 ;
    wire new_AGEMA_signal_26021 ;
    wire new_AGEMA_signal_26022 ;
    wire new_AGEMA_signal_26023 ;
    wire new_AGEMA_signal_26024 ;
    wire new_AGEMA_signal_26025 ;
    wire new_AGEMA_signal_26026 ;
    wire new_AGEMA_signal_26027 ;
    wire new_AGEMA_signal_26028 ;
    wire new_AGEMA_signal_26029 ;
    wire new_AGEMA_signal_26030 ;
    wire new_AGEMA_signal_26031 ;
    wire new_AGEMA_signal_26032 ;
    wire new_AGEMA_signal_26033 ;
    wire new_AGEMA_signal_26034 ;
    wire new_AGEMA_signal_26035 ;
    wire new_AGEMA_signal_26036 ;
    wire new_AGEMA_signal_26037 ;
    wire new_AGEMA_signal_26038 ;
    wire new_AGEMA_signal_26039 ;
    wire new_AGEMA_signal_26040 ;
    wire new_AGEMA_signal_26041 ;
    wire new_AGEMA_signal_26042 ;
    wire new_AGEMA_signal_26043 ;
    wire new_AGEMA_signal_26044 ;
    wire new_AGEMA_signal_26045 ;
    wire new_AGEMA_signal_26046 ;
    wire new_AGEMA_signal_26047 ;
    wire new_AGEMA_signal_26048 ;
    wire new_AGEMA_signal_26049 ;
    wire new_AGEMA_signal_26050 ;
    wire new_AGEMA_signal_26051 ;
    wire new_AGEMA_signal_26052 ;
    wire new_AGEMA_signal_26053 ;
    wire new_AGEMA_signal_26054 ;
    wire new_AGEMA_signal_26055 ;
    wire new_AGEMA_signal_26056 ;
    wire new_AGEMA_signal_26057 ;
    wire new_AGEMA_signal_26058 ;
    wire new_AGEMA_signal_26059 ;
    wire new_AGEMA_signal_26060 ;
    wire new_AGEMA_signal_26061 ;
    wire new_AGEMA_signal_26062 ;
    wire new_AGEMA_signal_26063 ;
    wire new_AGEMA_signal_26064 ;
    wire new_AGEMA_signal_26065 ;
    wire new_AGEMA_signal_26066 ;
    wire new_AGEMA_signal_26067 ;
    wire new_AGEMA_signal_26068 ;
    wire new_AGEMA_signal_26069 ;
    wire new_AGEMA_signal_26070 ;
    wire new_AGEMA_signal_26071 ;
    wire new_AGEMA_signal_26072 ;
    wire new_AGEMA_signal_26073 ;
    wire new_AGEMA_signal_26074 ;
    wire new_AGEMA_signal_26075 ;
    wire new_AGEMA_signal_26076 ;
    wire new_AGEMA_signal_26077 ;
    wire new_AGEMA_signal_26078 ;
    wire new_AGEMA_signal_26079 ;
    wire new_AGEMA_signal_26080 ;
    wire new_AGEMA_signal_26081 ;
    wire new_AGEMA_signal_26082 ;
    wire new_AGEMA_signal_26083 ;
    wire new_AGEMA_signal_26084 ;
    wire new_AGEMA_signal_26085 ;
    wire new_AGEMA_signal_26086 ;
    wire new_AGEMA_signal_26087 ;
    wire new_AGEMA_signal_26088 ;
    wire new_AGEMA_signal_26089 ;
    wire new_AGEMA_signal_26090 ;
    wire new_AGEMA_signal_26091 ;
    wire new_AGEMA_signal_26092 ;
    wire new_AGEMA_signal_26093 ;
    wire new_AGEMA_signal_26094 ;
    wire new_AGEMA_signal_26095 ;
    wire new_AGEMA_signal_26096 ;
    wire new_AGEMA_signal_26097 ;
    wire new_AGEMA_signal_26098 ;
    wire new_AGEMA_signal_26099 ;
    wire new_AGEMA_signal_26100 ;
    wire new_AGEMA_signal_26101 ;
    wire new_AGEMA_signal_26102 ;
    wire new_AGEMA_signal_26103 ;
    wire new_AGEMA_signal_26104 ;
    wire new_AGEMA_signal_26105 ;
    wire new_AGEMA_signal_26106 ;
    wire new_AGEMA_signal_26107 ;
    wire new_AGEMA_signal_26108 ;
    wire new_AGEMA_signal_26109 ;
    wire new_AGEMA_signal_26110 ;
    wire new_AGEMA_signal_26111 ;
    wire new_AGEMA_signal_26112 ;
    wire new_AGEMA_signal_26113 ;
    wire new_AGEMA_signal_26114 ;
    wire new_AGEMA_signal_26115 ;
    wire new_AGEMA_signal_26116 ;
    wire new_AGEMA_signal_26117 ;
    wire new_AGEMA_signal_26118 ;
    wire new_AGEMA_signal_26119 ;
    wire new_AGEMA_signal_26120 ;
    wire new_AGEMA_signal_26121 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) U1938 ( .a ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1939 ( .a ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1940 ( .a ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, new_AGEMA_signal_962, n2462}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1941 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1942 ( .a ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1944 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1945 ( .a ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, n2630}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1946 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_17702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_17704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( new_AGEMA_signal_17706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s3[4] ), .Q ( new_AGEMA_signal_17708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s4[4] ), .Q ( new_AGEMA_signal_17710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_17712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_17714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( new_AGEMA_signal_17716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( SI_s3[6] ), .Q ( new_AGEMA_signal_17718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( SI_s4[6] ), .Q ( new_AGEMA_signal_17720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_17722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_17724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( new_AGEMA_signal_17726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( SI_s3[7] ), .Q ( new_AGEMA_signal_17728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( SI_s4[7] ), .Q ( new_AGEMA_signal_17730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_17732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_17734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( new_AGEMA_signal_17736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( new_AGEMA_signal_17738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( SI_s4[0] ), .Q ( new_AGEMA_signal_17740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_17742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_17744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_17746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_17748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( SI_s4[1] ), .Q ( new_AGEMA_signal_17750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_17752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_17754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_17756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_17758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_17760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_17762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_17764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( new_AGEMA_signal_17766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( SI_s3[5] ), .Q ( new_AGEMA_signal_17768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( SI_s4[5] ), .Q ( new_AGEMA_signal_17770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_17772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( new_AGEMA_signal_962 ), .Q ( new_AGEMA_signal_17774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( new_AGEMA_signal_963 ), .Q ( new_AGEMA_signal_17776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_17778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( new_AGEMA_signal_965 ), .Q ( new_AGEMA_signal_17780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_17782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_17784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_17786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( new_AGEMA_signal_972 ), .Q ( new_AGEMA_signal_17788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( new_AGEMA_signal_973 ), .Q ( new_AGEMA_signal_17790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_17792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( new_AGEMA_signal_946 ), .Q ( new_AGEMA_signal_17794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_17796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( new_AGEMA_signal_948 ), .Q ( new_AGEMA_signal_17798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( new_AGEMA_signal_949 ), .Q ( new_AGEMA_signal_17800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_17802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( new_AGEMA_signal_1002 ), .Q ( new_AGEMA_signal_17804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_17806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_17808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_17810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_17812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( new_AGEMA_signal_978 ), .Q ( new_AGEMA_signal_17814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( new_AGEMA_signal_979 ), .Q ( new_AGEMA_signal_17816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( new_AGEMA_signal_980 ), .Q ( new_AGEMA_signal_17818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_17820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_17822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_17824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_17826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_17828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( SI_s4[3] ), .Q ( new_AGEMA_signal_17830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_17832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( new_AGEMA_signal_986 ), .Q ( new_AGEMA_signal_17834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_17836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_17838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_17840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_17842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( new_AGEMA_signal_954 ), .Q ( new_AGEMA_signal_17844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( new_AGEMA_signal_955 ), .Q ( new_AGEMA_signal_17846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( new_AGEMA_signal_956 ), .Q ( new_AGEMA_signal_17848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_17850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_19132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_19138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_19144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_19150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( SI_s4[2] ), .Q ( new_AGEMA_signal_19156 ) ) ;

    /* cells in depth 2 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1937 ( .ina ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}), .inb ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, n2624}), .b ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1947 ( .ina ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15]}), .outt ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1948 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, new_AGEMA_signal_962, n2462}), .inb ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1949 ( .ina ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45]}), .outt ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1950 ( .ina ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .b ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1952 ( .ina ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75]}), .outt ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}), .b ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2640}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1955 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, n2630}), .clk ( clk ), .rnd ({Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2699}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2699}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1957 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105]}), .outt ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}), .b ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1961 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1963 ( .ina ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135]}), .outt ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2317}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1965 ( .ina ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .inb ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .clk ( clk ), .rnd ({Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1969 ( .ina ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .inb ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165]}), .outt ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, n2073}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, n2073}), .b ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1971 ( .ina ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1972 ( .ina ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195]}), .outt ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}), .b ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1975 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .inb ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2723}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2723}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1978 ( .ina ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .inb ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225]}), .outt ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2541}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1984 ( .ina ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .inb ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, n2086}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1987 ( .ina ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .inb ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .clk ( clk ), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255]}), .outt ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2600}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1990 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, new_AGEMA_signal_962, n2462}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2538}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2538}), .b ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1995 ( .ina ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285]}), .outt ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2595}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2595}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1999 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, n2630}), .clk ( clk ), .rnd ({Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2753}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2753}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2577}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2004 ( .ina ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .inb ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315]}), .outt ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2400}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2008 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, n2785}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, n2785}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2013 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .inb ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345]}), .outt ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2609}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2609}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, new_AGEMA_signal_1334, n2724}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2017 ( .ina ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .clk ( clk ), .rnd ({Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2661}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2661}), .b ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2174}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2020 ( .ina ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375]}), .outt ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .b ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n2493}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2025 ( .ina ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2587}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .b ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2570}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2029 ( .ina ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405]}), .outt ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2035 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .outt ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .b ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2739}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2044 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, new_AGEMA_signal_962, n2462}), .inb ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}), .clk ( clk ), .rnd ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435]}), .outt ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2045 ( .ina ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .outt ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2052 ( .ina ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .clk ( clk ), .rnd ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465]}), .outt ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2452}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2068 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .outt ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2772}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2070 ( .ina ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495]}), .outt ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2400}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2313}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2089 ( .ina ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .inb ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .clk ( clk ), .rnd ({Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .outt ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2395}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2395}), .b ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2094 ( .ina ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525]}), .outt ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2779}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2096 ( .ina ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, n2630}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .clk ( clk ), .rnd ({Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .outt ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, n2624}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2097 ( .ina ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555]}), .outt ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2242}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2100 ( .ina ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .clk ( clk ), .rnd ({Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .outt ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2356}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2772}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2823}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2122 ( .ina ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585]}), .outt ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}), .b ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2828}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2133 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .outt ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2616}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2616}), .b ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, n2679}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2138 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, n2760}), .clk ( clk ), .rnd ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615]}), .outt ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2563}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2563}), .b ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2809}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}), .b ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2709}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2163 ( .ina ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}), .inb ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .clk ( clk ), .rnd ({Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .outt ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2401}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2211 ( .ina ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .inb ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645]}), .outt ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, n2061}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2232 ( .ina ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, n2796}), .inb ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .clk ( clk ), .rnd ({Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .outt ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2721}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2276 ( .ina ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .inb ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2765}), .clk ( clk ), .rnd ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675]}), .outt ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2298}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2401}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2118}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2307 ( .ina ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, n2630}), .clk ( clk ), .rnd ({Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .outt ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, new_AGEMA_signal_1226, n2346}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2341 ( .ina ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_981, new_AGEMA_signal_980, new_AGEMA_signal_979, new_AGEMA_signal_978, n2791}), .clk ( clk ), .rnd ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705]}), .outt ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2430}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2383 ( .ina ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .outt ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2712}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2402 ( .ina ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, n2813}), .clk ( clk ), .rnd ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735]}), .outt ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n2777}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2615 ( .ina ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, new_AGEMA_signal_962, n2462}), .clk ( clk ), .rnd ({Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .outt ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, n2463}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2627 ( .ina ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, new_AGEMA_signal_954, n2810}), .inb ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765]}), .outt ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( new_AGEMA_signal_17702 ), .Q ( new_AGEMA_signal_17703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( new_AGEMA_signal_17704 ), .Q ( new_AGEMA_signal_17705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( new_AGEMA_signal_17706 ), .Q ( new_AGEMA_signal_17707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( new_AGEMA_signal_17708 ), .Q ( new_AGEMA_signal_17709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( new_AGEMA_signal_17710 ), .Q ( new_AGEMA_signal_17711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_17712 ), .Q ( new_AGEMA_signal_17713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( new_AGEMA_signal_17714 ), .Q ( new_AGEMA_signal_17715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_17716 ), .Q ( new_AGEMA_signal_17717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_17718 ), .Q ( new_AGEMA_signal_17719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_17720 ), .Q ( new_AGEMA_signal_17721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_17722 ), .Q ( new_AGEMA_signal_17723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_17724 ), .Q ( new_AGEMA_signal_17725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( new_AGEMA_signal_17726 ), .Q ( new_AGEMA_signal_17727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_17728 ), .Q ( new_AGEMA_signal_17729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_17730 ), .Q ( new_AGEMA_signal_17731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_17732 ), .Q ( new_AGEMA_signal_17733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_17734 ), .Q ( new_AGEMA_signal_17735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_17736 ), .Q ( new_AGEMA_signal_17737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_17738 ), .Q ( new_AGEMA_signal_17739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_17740 ), .Q ( new_AGEMA_signal_17741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_17742 ), .Q ( new_AGEMA_signal_17743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_17744 ), .Q ( new_AGEMA_signal_17745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_17746 ), .Q ( new_AGEMA_signal_17747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_17748 ), .Q ( new_AGEMA_signal_17749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_17750 ), .Q ( new_AGEMA_signal_17751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_17752 ), .Q ( new_AGEMA_signal_17753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_17754 ), .Q ( new_AGEMA_signal_17755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_17756 ), .Q ( new_AGEMA_signal_17757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_17758 ), .Q ( new_AGEMA_signal_17759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_17760 ), .Q ( new_AGEMA_signal_17761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_17762 ), .Q ( new_AGEMA_signal_17763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_17764 ), .Q ( new_AGEMA_signal_17765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_17766 ), .Q ( new_AGEMA_signal_17767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_17768 ), .Q ( new_AGEMA_signal_17769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_17770 ), .Q ( new_AGEMA_signal_17771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_17772 ), .Q ( new_AGEMA_signal_17773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_17774 ), .Q ( new_AGEMA_signal_17775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_17776 ), .Q ( new_AGEMA_signal_17777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_17778 ), .Q ( new_AGEMA_signal_17779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_17780 ), .Q ( new_AGEMA_signal_17781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_17782 ), .Q ( new_AGEMA_signal_17783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_17784 ), .Q ( new_AGEMA_signal_17785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_17786 ), .Q ( new_AGEMA_signal_17787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_17788 ), .Q ( new_AGEMA_signal_17789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_17790 ), .Q ( new_AGEMA_signal_17791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_17792 ), .Q ( new_AGEMA_signal_17793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_17794 ), .Q ( new_AGEMA_signal_17795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_17796 ), .Q ( new_AGEMA_signal_17797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_17798 ), .Q ( new_AGEMA_signal_17799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_17800 ), .Q ( new_AGEMA_signal_17801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_17802 ), .Q ( new_AGEMA_signal_17803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_17804 ), .Q ( new_AGEMA_signal_17805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_17806 ), .Q ( new_AGEMA_signal_17807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_17808 ), .Q ( new_AGEMA_signal_17809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_17810 ), .Q ( new_AGEMA_signal_17811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_17812 ), .Q ( new_AGEMA_signal_17813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_17814 ), .Q ( new_AGEMA_signal_17815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_17816 ), .Q ( new_AGEMA_signal_17817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_17818 ), .Q ( new_AGEMA_signal_17819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_17820 ), .Q ( new_AGEMA_signal_17821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_17822 ), .Q ( new_AGEMA_signal_17823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_17824 ), .Q ( new_AGEMA_signal_17825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_17826 ), .Q ( new_AGEMA_signal_17827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_17828 ), .Q ( new_AGEMA_signal_17829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_17830 ), .Q ( new_AGEMA_signal_17831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_17832 ), .Q ( new_AGEMA_signal_17833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_17834 ), .Q ( new_AGEMA_signal_17835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_17836 ), .Q ( new_AGEMA_signal_17837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_17838 ), .Q ( new_AGEMA_signal_17839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_17840 ), .Q ( new_AGEMA_signal_17841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_17842 ), .Q ( new_AGEMA_signal_17843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_17844 ), .Q ( new_AGEMA_signal_17845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_17846 ), .Q ( new_AGEMA_signal_17847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_17848 ), .Q ( new_AGEMA_signal_17849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_17850 ), .Q ( new_AGEMA_signal_17851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_19132 ), .Q ( new_AGEMA_signal_19133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_19138 ), .Q ( new_AGEMA_signal_19139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_19144 ), .Q ( new_AGEMA_signal_19145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_19150 ), .Q ( new_AGEMA_signal_19151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_19156 ), .Q ( new_AGEMA_signal_19157 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_17852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( new_AGEMA_signal_1286 ), .Q ( new_AGEMA_signal_17854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( new_AGEMA_signal_1287 ), .Q ( new_AGEMA_signal_17856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( new_AGEMA_signal_1288 ), .Q ( new_AGEMA_signal_17858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( new_AGEMA_signal_1289 ), .Q ( new_AGEMA_signal_17860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( new_AGEMA_signal_17823 ), .Q ( new_AGEMA_signal_17862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( new_AGEMA_signal_17825 ), .Q ( new_AGEMA_signal_17864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( new_AGEMA_signal_17827 ), .Q ( new_AGEMA_signal_17866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( new_AGEMA_signal_17829 ), .Q ( new_AGEMA_signal_17868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( new_AGEMA_signal_17831 ), .Q ( new_AGEMA_signal_17870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( new_AGEMA_signal_17713 ), .Q ( new_AGEMA_signal_17872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( new_AGEMA_signal_17715 ), .Q ( new_AGEMA_signal_17874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( new_AGEMA_signal_17717 ), .Q ( new_AGEMA_signal_17876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( new_AGEMA_signal_17719 ), .Q ( new_AGEMA_signal_17878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( new_AGEMA_signal_17721 ), .Q ( new_AGEMA_signal_17880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_17882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( new_AGEMA_signal_1338 ), .Q ( new_AGEMA_signal_17884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( new_AGEMA_signal_1339 ), .Q ( new_AGEMA_signal_17886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( new_AGEMA_signal_1340 ), .Q ( new_AGEMA_signal_17888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( new_AGEMA_signal_1341 ), .Q ( new_AGEMA_signal_17890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( new_AGEMA_signal_17703 ), .Q ( new_AGEMA_signal_17892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( new_AGEMA_signal_17705 ), .Q ( new_AGEMA_signal_17894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_17707 ), .Q ( new_AGEMA_signal_17896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( new_AGEMA_signal_17709 ), .Q ( new_AGEMA_signal_17898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( new_AGEMA_signal_17711 ), .Q ( new_AGEMA_signal_17900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( new_AGEMA_signal_17733 ), .Q ( new_AGEMA_signal_17902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( new_AGEMA_signal_17735 ), .Q ( new_AGEMA_signal_17904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( new_AGEMA_signal_17737 ), .Q ( new_AGEMA_signal_17906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( new_AGEMA_signal_17739 ), .Q ( new_AGEMA_signal_17908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( new_AGEMA_signal_17741 ), .Q ( new_AGEMA_signal_17910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_17912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( new_AGEMA_signal_1350 ), .Q ( new_AGEMA_signal_17914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( new_AGEMA_signal_1351 ), .Q ( new_AGEMA_signal_17916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( new_AGEMA_signal_1352 ), .Q ( new_AGEMA_signal_17918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( new_AGEMA_signal_1353 ), .Q ( new_AGEMA_signal_17920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_17922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_1330 ), .Q ( new_AGEMA_signal_17924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( new_AGEMA_signal_1331 ), .Q ( new_AGEMA_signal_17926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( new_AGEMA_signal_1332 ), .Q ( new_AGEMA_signal_17928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( new_AGEMA_signal_1333 ), .Q ( new_AGEMA_signal_17930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_17932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_17934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_17936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_17938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( new_AGEMA_signal_1009 ), .Q ( new_AGEMA_signal_17940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_17942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_1146 ), .Q ( new_AGEMA_signal_17944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( new_AGEMA_signal_1147 ), .Q ( new_AGEMA_signal_17946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( new_AGEMA_signal_1148 ), .Q ( new_AGEMA_signal_17948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( new_AGEMA_signal_1149 ), .Q ( new_AGEMA_signal_17950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_17952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_17954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( new_AGEMA_signal_1103 ), .Q ( new_AGEMA_signal_17956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( new_AGEMA_signal_1104 ), .Q ( new_AGEMA_signal_17958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( new_AGEMA_signal_1105 ), .Q ( new_AGEMA_signal_17960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_17962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_17964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_17966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_17968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( new_AGEMA_signal_1033 ), .Q ( new_AGEMA_signal_17970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_17972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( new_AGEMA_signal_1406 ), .Q ( new_AGEMA_signal_17974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_1407 ), .Q ( new_AGEMA_signal_17976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( new_AGEMA_signal_1408 ), .Q ( new_AGEMA_signal_17978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_1409 ), .Q ( new_AGEMA_signal_17980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_17982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( new_AGEMA_signal_1010 ), .Q ( new_AGEMA_signal_17984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( new_AGEMA_signal_1011 ), .Q ( new_AGEMA_signal_17986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( new_AGEMA_signal_1012 ), .Q ( new_AGEMA_signal_17988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( new_AGEMA_signal_1013 ), .Q ( new_AGEMA_signal_17990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_17992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( new_AGEMA_signal_1314 ), .Q ( new_AGEMA_signal_17994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( new_AGEMA_signal_1315 ), .Q ( new_AGEMA_signal_17996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( new_AGEMA_signal_1316 ), .Q ( new_AGEMA_signal_17998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_1317 ), .Q ( new_AGEMA_signal_18000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_18002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_18004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( new_AGEMA_signal_1127 ), .Q ( new_AGEMA_signal_18006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( new_AGEMA_signal_1128 ), .Q ( new_AGEMA_signal_18008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( new_AGEMA_signal_1129 ), .Q ( new_AGEMA_signal_18010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_17743 ), .Q ( new_AGEMA_signal_18012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( new_AGEMA_signal_17745 ), .Q ( new_AGEMA_signal_18014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( new_AGEMA_signal_17747 ), .Q ( new_AGEMA_signal_18016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( new_AGEMA_signal_17749 ), .Q ( new_AGEMA_signal_18018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( new_AGEMA_signal_17751 ), .Q ( new_AGEMA_signal_18020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_18022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( new_AGEMA_signal_1106 ), .Q ( new_AGEMA_signal_18024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_18026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_18028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( new_AGEMA_signal_1109 ), .Q ( new_AGEMA_signal_18030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_18032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_18034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_1099 ), .Q ( new_AGEMA_signal_18036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( new_AGEMA_signal_1100 ), .Q ( new_AGEMA_signal_18038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( new_AGEMA_signal_1101 ), .Q ( new_AGEMA_signal_18040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_18042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_18044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_18046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_1448 ), .Q ( new_AGEMA_signal_18048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( new_AGEMA_signal_1449 ), .Q ( new_AGEMA_signal_18050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_18052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( new_AGEMA_signal_1122 ), .Q ( new_AGEMA_signal_18054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( new_AGEMA_signal_1123 ), .Q ( new_AGEMA_signal_18056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( new_AGEMA_signal_1124 ), .Q ( new_AGEMA_signal_18058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_1125 ), .Q ( new_AGEMA_signal_18060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_18062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( new_AGEMA_signal_1206 ), .Q ( new_AGEMA_signal_18064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( new_AGEMA_signal_1207 ), .Q ( new_AGEMA_signal_18066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( new_AGEMA_signal_1208 ), .Q ( new_AGEMA_signal_18068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_18070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_17803 ), .Q ( new_AGEMA_signal_18072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( new_AGEMA_signal_17805 ), .Q ( new_AGEMA_signal_18074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_17807 ), .Q ( new_AGEMA_signal_18076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( new_AGEMA_signal_17809 ), .Q ( new_AGEMA_signal_18078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( new_AGEMA_signal_17811 ), .Q ( new_AGEMA_signal_18080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( new_AGEMA_signal_17753 ), .Q ( new_AGEMA_signal_18082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_17755 ), .Q ( new_AGEMA_signal_18084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( new_AGEMA_signal_17757 ), .Q ( new_AGEMA_signal_18086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_17759 ), .Q ( new_AGEMA_signal_18088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( new_AGEMA_signal_17761 ), .Q ( new_AGEMA_signal_18090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_18092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_18094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_18096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_18098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_18100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_18102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( new_AGEMA_signal_1150 ), .Q ( new_AGEMA_signal_18104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( new_AGEMA_signal_1151 ), .Q ( new_AGEMA_signal_18106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_1152 ), .Q ( new_AGEMA_signal_18108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( new_AGEMA_signal_1153 ), .Q ( new_AGEMA_signal_18110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_18112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( new_AGEMA_signal_1202 ), .Q ( new_AGEMA_signal_18114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( new_AGEMA_signal_1203 ), .Q ( new_AGEMA_signal_18116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( new_AGEMA_signal_1204 ), .Q ( new_AGEMA_signal_18118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_1205 ), .Q ( new_AGEMA_signal_18120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_18122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( new_AGEMA_signal_1386 ), .Q ( new_AGEMA_signal_18124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( new_AGEMA_signal_1387 ), .Q ( new_AGEMA_signal_18126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( new_AGEMA_signal_1388 ), .Q ( new_AGEMA_signal_18128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( new_AGEMA_signal_1389 ), .Q ( new_AGEMA_signal_18130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_18132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( new_AGEMA_signal_1178 ), .Q ( new_AGEMA_signal_18134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( new_AGEMA_signal_1179 ), .Q ( new_AGEMA_signal_18136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( new_AGEMA_signal_1180 ), .Q ( new_AGEMA_signal_18138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( new_AGEMA_signal_1181 ), .Q ( new_AGEMA_signal_18140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_18142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_18144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_18146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_1076 ), .Q ( new_AGEMA_signal_18148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( new_AGEMA_signal_1077 ), .Q ( new_AGEMA_signal_18150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_18152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( new_AGEMA_signal_1090 ), .Q ( new_AGEMA_signal_18154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_18156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_18158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_1093 ), .Q ( new_AGEMA_signal_18160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_18162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( new_AGEMA_signal_1014 ), .Q ( new_AGEMA_signal_18164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( new_AGEMA_signal_1015 ), .Q ( new_AGEMA_signal_18166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_1016 ), .Q ( new_AGEMA_signal_18168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_18170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_18172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( new_AGEMA_signal_1198 ), .Q ( new_AGEMA_signal_18174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( new_AGEMA_signal_1199 ), .Q ( new_AGEMA_signal_18176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( new_AGEMA_signal_1200 ), .Q ( new_AGEMA_signal_18178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( new_AGEMA_signal_1201 ), .Q ( new_AGEMA_signal_18180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( new_AGEMA_signal_17813 ), .Q ( new_AGEMA_signal_18182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( new_AGEMA_signal_17815 ), .Q ( new_AGEMA_signal_18184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( new_AGEMA_signal_17817 ), .Q ( new_AGEMA_signal_18186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( new_AGEMA_signal_17819 ), .Q ( new_AGEMA_signal_18188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( new_AGEMA_signal_17821 ), .Q ( new_AGEMA_signal_18190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_18192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( new_AGEMA_signal_1078 ), .Q ( new_AGEMA_signal_18194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_18196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( new_AGEMA_signal_1080 ), .Q ( new_AGEMA_signal_18198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_18200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( new_AGEMA_signal_17833 ), .Q ( new_AGEMA_signal_18202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( new_AGEMA_signal_17835 ), .Q ( new_AGEMA_signal_18204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( new_AGEMA_signal_17837 ), .Q ( new_AGEMA_signal_18206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( new_AGEMA_signal_17839 ), .Q ( new_AGEMA_signal_18208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( new_AGEMA_signal_17841 ), .Q ( new_AGEMA_signal_18210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_18212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( new_AGEMA_signal_1118 ), .Q ( new_AGEMA_signal_18214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_18216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_18218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( new_AGEMA_signal_1121 ), .Q ( new_AGEMA_signal_18220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_18222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( new_AGEMA_signal_1334 ), .Q ( new_AGEMA_signal_18224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( new_AGEMA_signal_1335 ), .Q ( new_AGEMA_signal_18226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( new_AGEMA_signal_1336 ), .Q ( new_AGEMA_signal_18228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_1337 ), .Q ( new_AGEMA_signal_18230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_18232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_1082 ), .Q ( new_AGEMA_signal_18234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( new_AGEMA_signal_1083 ), .Q ( new_AGEMA_signal_18236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_18238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_18240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_18242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_1298 ), .Q ( new_AGEMA_signal_18244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( new_AGEMA_signal_1299 ), .Q ( new_AGEMA_signal_18246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( new_AGEMA_signal_1300 ), .Q ( new_AGEMA_signal_18248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_1301 ), .Q ( new_AGEMA_signal_18250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_18252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( new_AGEMA_signal_1134 ), .Q ( new_AGEMA_signal_18254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_1135 ), .Q ( new_AGEMA_signal_18256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_1136 ), .Q ( new_AGEMA_signal_18258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( new_AGEMA_signal_1137 ), .Q ( new_AGEMA_signal_18260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_18262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_1266 ), .Q ( new_AGEMA_signal_18264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( new_AGEMA_signal_1267 ), .Q ( new_AGEMA_signal_18266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_1268 ), .Q ( new_AGEMA_signal_18268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( new_AGEMA_signal_1269 ), .Q ( new_AGEMA_signal_18270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_18272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( new_AGEMA_signal_1270 ), .Q ( new_AGEMA_signal_18274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( new_AGEMA_signal_1271 ), .Q ( new_AGEMA_signal_18276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( new_AGEMA_signal_1272 ), .Q ( new_AGEMA_signal_18278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( new_AGEMA_signal_1273 ), .Q ( new_AGEMA_signal_18280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_18282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_1094 ), .Q ( new_AGEMA_signal_18284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( new_AGEMA_signal_1095 ), .Q ( new_AGEMA_signal_18286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_1096 ), .Q ( new_AGEMA_signal_18288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( new_AGEMA_signal_1097 ), .Q ( new_AGEMA_signal_18290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_18292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( new_AGEMA_signal_1242 ), .Q ( new_AGEMA_signal_18294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_1243 ), .Q ( new_AGEMA_signal_18296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_1244 ), .Q ( new_AGEMA_signal_18298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( new_AGEMA_signal_1245 ), .Q ( new_AGEMA_signal_18300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_18302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_1282 ), .Q ( new_AGEMA_signal_18304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_1283 ), .Q ( new_AGEMA_signal_18306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( new_AGEMA_signal_1284 ), .Q ( new_AGEMA_signal_18308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( new_AGEMA_signal_1285 ), .Q ( new_AGEMA_signal_18310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_18312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( new_AGEMA_signal_1138 ), .Q ( new_AGEMA_signal_18314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_1139 ), .Q ( new_AGEMA_signal_18316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( new_AGEMA_signal_1140 ), .Q ( new_AGEMA_signal_18318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( new_AGEMA_signal_1141 ), .Q ( new_AGEMA_signal_18320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_17773 ), .Q ( new_AGEMA_signal_18322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_17775 ), .Q ( new_AGEMA_signal_18324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( new_AGEMA_signal_17777 ), .Q ( new_AGEMA_signal_18326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( new_AGEMA_signal_17779 ), .Q ( new_AGEMA_signal_18328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( new_AGEMA_signal_17781 ), .Q ( new_AGEMA_signal_18330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_18332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_18334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_1087 ), .Q ( new_AGEMA_signal_18336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( new_AGEMA_signal_1088 ), .Q ( new_AGEMA_signal_18338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_1089 ), .Q ( new_AGEMA_signal_18340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( new_AGEMA_signal_17783 ), .Q ( new_AGEMA_signal_18342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( new_AGEMA_signal_17785 ), .Q ( new_AGEMA_signal_18344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( new_AGEMA_signal_17787 ), .Q ( new_AGEMA_signal_18346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_17789 ), .Q ( new_AGEMA_signal_18348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( new_AGEMA_signal_17791 ), .Q ( new_AGEMA_signal_18350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_18352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( new_AGEMA_signal_1022 ), .Q ( new_AGEMA_signal_18354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( new_AGEMA_signal_1023 ), .Q ( new_AGEMA_signal_18356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( new_AGEMA_signal_1024 ), .Q ( new_AGEMA_signal_18358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( new_AGEMA_signal_1025 ), .Q ( new_AGEMA_signal_18360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( new_AGEMA_signal_17843 ), .Q ( new_AGEMA_signal_18362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( new_AGEMA_signal_17845 ), .Q ( new_AGEMA_signal_18364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( new_AGEMA_signal_17847 ), .Q ( new_AGEMA_signal_18366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( new_AGEMA_signal_17849 ), .Q ( new_AGEMA_signal_18368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_17851 ), .Q ( new_AGEMA_signal_18370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_18372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( new_AGEMA_signal_1186 ), .Q ( new_AGEMA_signal_18374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_1187 ), .Q ( new_AGEMA_signal_18376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( new_AGEMA_signal_1188 ), .Q ( new_AGEMA_signal_18378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( new_AGEMA_signal_1189 ), .Q ( new_AGEMA_signal_18380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_18382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_18384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_18386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_1192 ), .Q ( new_AGEMA_signal_18388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_18390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_18392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_1162 ), .Q ( new_AGEMA_signal_18394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_1163 ), .Q ( new_AGEMA_signal_18396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( new_AGEMA_signal_1164 ), .Q ( new_AGEMA_signal_18398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_1165 ), .Q ( new_AGEMA_signal_18400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_18402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_1374 ), .Q ( new_AGEMA_signal_18404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( new_AGEMA_signal_1375 ), .Q ( new_AGEMA_signal_18406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_1376 ), .Q ( new_AGEMA_signal_18408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_1377 ), .Q ( new_AGEMA_signal_18410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_18412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( new_AGEMA_signal_1278 ), .Q ( new_AGEMA_signal_18414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( new_AGEMA_signal_1279 ), .Q ( new_AGEMA_signal_18416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( new_AGEMA_signal_1280 ), .Q ( new_AGEMA_signal_18418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_1281 ), .Q ( new_AGEMA_signal_18420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_18422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_18424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( new_AGEMA_signal_1059 ), .Q ( new_AGEMA_signal_18426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_18428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_18430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_18432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( new_AGEMA_signal_1054 ), .Q ( new_AGEMA_signal_18434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_1055 ), .Q ( new_AGEMA_signal_18436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( new_AGEMA_signal_1056 ), .Q ( new_AGEMA_signal_18438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( new_AGEMA_signal_1057 ), .Q ( new_AGEMA_signal_18440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_18442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_1290 ), .Q ( new_AGEMA_signal_18444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( new_AGEMA_signal_1291 ), .Q ( new_AGEMA_signal_18446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_1292 ), .Q ( new_AGEMA_signal_18448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( new_AGEMA_signal_1293 ), .Q ( new_AGEMA_signal_18450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_18452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( new_AGEMA_signal_1142 ), .Q ( new_AGEMA_signal_18454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_1143 ), .Q ( new_AGEMA_signal_18456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( new_AGEMA_signal_1144 ), .Q ( new_AGEMA_signal_18458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_1145 ), .Q ( new_AGEMA_signal_18460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_18462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( new_AGEMA_signal_1322 ), .Q ( new_AGEMA_signal_18464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1323 ), .Q ( new_AGEMA_signal_18466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_18468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( new_AGEMA_signal_1325 ), .Q ( new_AGEMA_signal_18470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_18472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_1302 ), .Q ( new_AGEMA_signal_18474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( new_AGEMA_signal_1303 ), .Q ( new_AGEMA_signal_18476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( new_AGEMA_signal_1304 ), .Q ( new_AGEMA_signal_18478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_1305 ), .Q ( new_AGEMA_signal_18480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_18482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_18484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( new_AGEMA_signal_1439 ), .Q ( new_AGEMA_signal_18486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( new_AGEMA_signal_1440 ), .Q ( new_AGEMA_signal_18488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_18490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_18492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( new_AGEMA_signal_1070 ), .Q ( new_AGEMA_signal_18494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_18496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_18498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_18500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_18502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_18504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( new_AGEMA_signal_1195 ), .Q ( new_AGEMA_signal_18506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( new_AGEMA_signal_1196 ), .Q ( new_AGEMA_signal_18508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_18510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_18512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_1154 ), .Q ( new_AGEMA_signal_18514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_1155 ), .Q ( new_AGEMA_signal_18516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( new_AGEMA_signal_1156 ), .Q ( new_AGEMA_signal_18518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_18520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_18522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( new_AGEMA_signal_1174 ), .Q ( new_AGEMA_signal_18524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( new_AGEMA_signal_1175 ), .Q ( new_AGEMA_signal_18526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_1176 ), .Q ( new_AGEMA_signal_18528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( new_AGEMA_signal_1177 ), .Q ( new_AGEMA_signal_18530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_18552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_18556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_18560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_1356 ), .Q ( new_AGEMA_signal_18564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_1357 ), .Q ( new_AGEMA_signal_18568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_18682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( new_AGEMA_signal_1042 ), .Q ( new_AGEMA_signal_18686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( new_AGEMA_signal_1043 ), .Q ( new_AGEMA_signal_18690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_18694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_18698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_18772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( new_AGEMA_signal_1218 ), .Q ( new_AGEMA_signal_18776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_1219 ), .Q ( new_AGEMA_signal_18780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_18784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_18788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_18842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( new_AGEMA_signal_1426 ), .Q ( new_AGEMA_signal_18846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( new_AGEMA_signal_1427 ), .Q ( new_AGEMA_signal_18850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( new_AGEMA_signal_1428 ), .Q ( new_AGEMA_signal_18854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( new_AGEMA_signal_1429 ), .Q ( new_AGEMA_signal_18858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_18892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( new_AGEMA_signal_1226 ), .Q ( new_AGEMA_signal_18896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_1227 ), .Q ( new_AGEMA_signal_18900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_1228 ), .Q ( new_AGEMA_signal_18904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( new_AGEMA_signal_1229 ), .Q ( new_AGEMA_signal_18908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_18942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( new_AGEMA_signal_1018 ), .Q ( new_AGEMA_signal_18946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( new_AGEMA_signal_1019 ), .Q ( new_AGEMA_signal_18950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( new_AGEMA_signal_1020 ), .Q ( new_AGEMA_signal_18954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( new_AGEMA_signal_1021 ), .Q ( new_AGEMA_signal_18958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( new_AGEMA_signal_19133 ), .Q ( new_AGEMA_signal_19134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_19139 ), .Q ( new_AGEMA_signal_19140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( new_AGEMA_signal_19145 ), .Q ( new_AGEMA_signal_19146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_19151 ), .Q ( new_AGEMA_signal_19152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( new_AGEMA_signal_19157 ), .Q ( new_AGEMA_signal_19158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_17723 ), .Q ( new_AGEMA_signal_19192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( new_AGEMA_signal_17725 ), .Q ( new_AGEMA_signal_19196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_17727 ), .Q ( new_AGEMA_signal_19200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_17729 ), .Q ( new_AGEMA_signal_19204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( new_AGEMA_signal_17731 ), .Q ( new_AGEMA_signal_19208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_19242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_1110 ), .Q ( new_AGEMA_signal_19246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( new_AGEMA_signal_1111 ), .Q ( new_AGEMA_signal_19250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( new_AGEMA_signal_1112 ), .Q ( new_AGEMA_signal_19254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_19258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_19332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_1062 ), .Q ( new_AGEMA_signal_19336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_19340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_19344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_19348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_17793 ), .Q ( new_AGEMA_signal_19372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( new_AGEMA_signal_17795 ), .Q ( new_AGEMA_signal_19376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_17797 ), .Q ( new_AGEMA_signal_19380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_17799 ), .Q ( new_AGEMA_signal_19384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C ( clk ), .D ( new_AGEMA_signal_17801 ), .Q ( new_AGEMA_signal_19388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_19742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C ( clk ), .D ( new_AGEMA_signal_1274 ), .Q ( new_AGEMA_signal_19748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_19754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C ( clk ), .D ( new_AGEMA_signal_1276 ), .Q ( new_AGEMA_signal_19760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C ( clk ), .D ( new_AGEMA_signal_1277 ), .Q ( new_AGEMA_signal_19766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_19872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C ( clk ), .D ( new_AGEMA_signal_1130 ), .Q ( new_AGEMA_signal_19878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C ( clk ), .D ( new_AGEMA_signal_1131 ), .Q ( new_AGEMA_signal_19884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_19890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_19896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_20452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_20460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_20468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_20476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_20484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_20502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C ( clk ), .D ( new_AGEMA_signal_1158 ), .Q ( new_AGEMA_signal_20510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C ( clk ), .D ( new_AGEMA_signal_1159 ), .Q ( new_AGEMA_signal_20518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C ( clk ), .D ( new_AGEMA_signal_1160 ), .Q ( new_AGEMA_signal_20526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C ( clk ), .D ( new_AGEMA_signal_1161 ), .Q ( new_AGEMA_signal_20534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_20882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C ( clk ), .D ( new_AGEMA_signal_1434 ), .Q ( new_AGEMA_signal_20890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C ( clk ), .D ( new_AGEMA_signal_1435 ), .Q ( new_AGEMA_signal_20898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C ( clk ), .D ( new_AGEMA_signal_1436 ), .Q ( new_AGEMA_signal_20906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C ( clk ), .D ( new_AGEMA_signal_1437 ), .Q ( new_AGEMA_signal_20914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_21312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C ( clk ), .D ( new_AGEMA_signal_1114 ), .Q ( new_AGEMA_signal_21320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C ( clk ), .D ( new_AGEMA_signal_1115 ), .Q ( new_AGEMA_signal_21328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C ( clk ), .D ( new_AGEMA_signal_1116 ), .Q ( new_AGEMA_signal_21336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C ( clk ), .D ( new_AGEMA_signal_1117 ), .Q ( new_AGEMA_signal_21344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_21462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C ( clk ), .D ( new_AGEMA_signal_1442 ), .Q ( new_AGEMA_signal_21470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C ( clk ), .D ( new_AGEMA_signal_1443 ), .Q ( new_AGEMA_signal_21478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C ( clk ), .D ( new_AGEMA_signal_1444 ), .Q ( new_AGEMA_signal_21486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C ( clk ), .D ( new_AGEMA_signal_1445 ), .Q ( new_AGEMA_signal_21494 ) ) ;

    /* cells in depth 4 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1954 ( .ina ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .inb ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2640}), .clk ( clk ), .rnd ({Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .outt ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, n2575}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1959 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}), .inb ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .clk ( clk ), .rnd ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795]}), .outt ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n1962}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1964 ( .ina ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2317}), .clk ( clk ), .rnd ({Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .outt ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, n1922}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1974 ( .ina ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .clk ( clk ), .rnd ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825]}), .outt ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, new_AGEMA_signal_1294, n2755}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1977 ( .ina ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2317}), .inb ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}), .clk ( clk ), .rnd ({Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .outt ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1694, n1926}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1980 ( .ina ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .inb ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2541}), .clk ( clk ), .rnd ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855]}), .outt ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n1925}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1986 ( .ina ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, n2086}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2317}), .clk ( clk ), .rnd ({Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .outt ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, n2151}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1988 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}), .inb ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2600}), .clk ( clk ), .rnd ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885]}), .outt ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2631}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2631}), .b ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2734}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1992 ( .ina ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .inb ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .clk ( clk ), .rnd ({Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .outt ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2763}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1997 ( .ina ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .clk ( clk ), .rnd ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915]}), .outt ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, new_AGEMA_signal_1318, n1930}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2005 ( .ina ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2400}), .inb ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .clk ( clk ), .rnd ({Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .outt ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2010 ( .ina ({new_AGEMA_signal_17711, new_AGEMA_signal_17709, new_AGEMA_signal_17707, new_AGEMA_signal_17705, new_AGEMA_signal_17703}), .inb ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .clk ( clk ), .rnd ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945]}), .outt ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1718, n1937}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2022 ( .ina ({new_AGEMA_signal_17721, new_AGEMA_signal_17719, new_AGEMA_signal_17717, new_AGEMA_signal_17715, new_AGEMA_signal_17713}), .inb ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n2493}), .clk ( clk ), .rnd ({Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .outt ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, new_AGEMA_signal_1343, new_AGEMA_signal_1342, n1942}) ) ;
    or_HPC1 #(.security_order(4), .pipeline(1)) U2026 ( .ina ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2587}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .clk ( clk ), .rnd ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975]}), .outt ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2676}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2030 ( .ina ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}), .clk ( clk ), .rnd ({Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .outt ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1730, n1944}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2037 ( .ina ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .inb ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}), .clk ( clk ), .rnd ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005]}), .outt ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n1950}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2039 ( .ina ({new_AGEMA_signal_17731, new_AGEMA_signal_17729, new_AGEMA_signal_17727, new_AGEMA_signal_17725, new_AGEMA_signal_17723}), .inb ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2739}), .clk ( clk ), .rnd ({Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .outt ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, n1949}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2042 ( .ina ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .inb ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2600}), .clk ( clk ), .rnd ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035]}), .outt ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2677}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2677}), .b ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2662}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2047 ( .ina ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}), .inb ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .clk ( clk ), .rnd ({Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .outt ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2053 ( .ina ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2452}), .clk ( clk ), .rnd ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065]}), .outt ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, new_AGEMA_signal_1370, n1957}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2056 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2600}), .clk ( clk ), .rnd ({Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .outt ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, n2088}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2062 ( .ina ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .inb ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .clk ( clk ), .rnd ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095]}), .outt ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n1964}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2063 ( .ina ({new_AGEMA_signal_17741, new_AGEMA_signal_17739, new_AGEMA_signal_17737, new_AGEMA_signal_17735, new_AGEMA_signal_17733}), .inb ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .clk ( clk ), .rnd ({Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .outt ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2736}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2069 ( .ina ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2772}), .inb ({new_AGEMA_signal_17751, new_AGEMA_signal_17749, new_AGEMA_signal_17747, new_AGEMA_signal_17745, new_AGEMA_signal_17743}), .clk ( clk ), .rnd ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125]}), .outt ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, n2673}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2072 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .clk ( clk ), .rnd ({Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .outt ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2720}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2075 ( .ina ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2313}), .inb ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .clk ( clk ), .rnd ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155]}), .outt ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, n2412}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, n2412}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2079 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}), .inb ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}), .clk ( clk ), .rnd ({Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .outt ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2571}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2571}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2505}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2081 ( .ina ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .inb ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}), .clk ( clk ), .rnd ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185]}), .outt ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2083 ( .ina ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .inb ({new_AGEMA_signal_17751, new_AGEMA_signal_17749, new_AGEMA_signal_17747, new_AGEMA_signal_17745, new_AGEMA_signal_17743}), .clk ( clk ), .rnd ({Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .outt ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, n2359}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2086 ( .ina ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .inb ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .clk ( clk ), .rnd ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215]}), .outt ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, new_AGEMA_signal_1402, n2101}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, new_AGEMA_signal_1402, n2101}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2625}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2091 ( .ina ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .inb ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2609}), .clk ( clk ), .rnd ({Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .outt ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2190}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2095 ( .ina ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2739}), .inb ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2779}), .clk ( clk ), .rnd ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245]}), .outt ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, new_AGEMA_signal_1415, new_AGEMA_signal_1414, n1976}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2098 ( .ina ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2242}), .clk ( clk ), .rnd ({Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .outt ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, n2535}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2101 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}), .inb ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2356}), .clk ( clk ), .rnd ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275]}), .outt ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, n1973}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2105 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .inb ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .clk ( clk ), .rnd ({Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .outt ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2690}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2111 ( .ina ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n2493}), .inb ({new_AGEMA_signal_17761, new_AGEMA_signal_17759, new_AGEMA_signal_17757, new_AGEMA_signal_17755, new_AGEMA_signal_17753}), .clk ( clk ), .rnd ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305]}), .outt ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2113 ( .ina ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .inb ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2779}), .clk ( clk ), .rnd ({Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .outt ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, n2741}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2118 ( .ina ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .inb ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .clk ( clk ), .rnd ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335]}), .outt ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, n1992}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2120 ( .ina ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2823}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .outt ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n1991}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2123 ( .ina ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .inb ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}), .clk ( clk ), .rnd ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365]}), .outt ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, n1993}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2125 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}), .inb ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .clk ( clk ), .rnd ({Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .outt ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, n1995}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2132 ( .ina ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .inb ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .clk ( clk ), .rnd ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395]}), .outt ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, n2241}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2135 ( .ina ({new_AGEMA_signal_17771, new_AGEMA_signal_17769, new_AGEMA_signal_17767, new_AGEMA_signal_17765, new_AGEMA_signal_17763}), .inb ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, n2679}), .clk ( clk ), .rnd ({Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .outt ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2003}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2140 ( .ina ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .inb ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2809}), .clk ( clk ), .rnd ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425]}), .outt ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, n2008}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2141 ( .ina ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, n2679}), .inb ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}), .clk ( clk ), .rnd ({Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .outt ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2572}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2143 ( .ina ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2809}), .inb ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2356}), .clk ( clk ), .rnd ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455]}), .outt ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2004}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2147 ( .ina ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .outt ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, n2009}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2151 ( .ina ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .inb ({new_AGEMA_signal_17761, new_AGEMA_signal_17759, new_AGEMA_signal_17757, new_AGEMA_signal_17755, new_AGEMA_signal_17753}), .clk ( clk ), .rnd ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485]}), .outt ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2157 ( .ina ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}), .clk ( clk ), .rnd ({Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .outt ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, n2026}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2158 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n2493}), .clk ( clk ), .rnd ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515]}), .outt ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2022}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2159 ( .ina ({new_AGEMA_signal_17781, new_AGEMA_signal_17779, new_AGEMA_signal_17777, new_AGEMA_signal_17775, new_AGEMA_signal_17773}), .inb ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .clk ( clk ), .rnd ({Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .outt ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, n2227}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2167 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .inb ({new_AGEMA_signal_17761, new_AGEMA_signal_17759, new_AGEMA_signal_17757, new_AGEMA_signal_17755, new_AGEMA_signal_17753}), .clk ( clk ), .rnd ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545]}), .outt ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, n2027}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2171 ( .ina ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .inb ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .clk ( clk ), .rnd ({Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .outt ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2214}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2173 ( .ina ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575]}), .outt ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, n2290}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2174 ( .ina ({new_AGEMA_signal_17741, new_AGEMA_signal_17739, new_AGEMA_signal_17737, new_AGEMA_signal_17735, new_AGEMA_signal_17733}), .inb ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .clk ( clk ), .rnd ({Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .outt ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2178 ( .ina ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .inb ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2400}), .clk ( clk ), .rnd ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605]}), .outt ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, new_AGEMA_signal_1462, n2034}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2182 ( .ina ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}), .inb ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .clk ( clk ), .rnd ({Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .outt ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, n2171}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2183 ( .ina ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2828}), .inb ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}), .clk ( clk ), .rnd ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635]}), .outt ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2039}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2188 ( .ina ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .outt ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1862, n2042}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2191 ( .ina ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .inb ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .clk ( clk ), .rnd ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665]}), .outt ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2754}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2192 ( .ina ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2313}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .clk ( clk ), .rnd ({Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .outt ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, n2044}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2198 ( .ina ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2313}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}), .clk ( clk ), .rnd ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695]}), .outt ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2654}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2202 ( .ina ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}), .inb ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2577}), .clk ( clk ), .rnd ({Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .outt ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2055}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2205 ( .ina ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2395}), .inb ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .clk ( clk ), .rnd ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725]}), .outt ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, n2057}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2208 ( .ina ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, n2679}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}), .clk ( clk ), .rnd ({Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .outt ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, n2407}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2212 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}), .inb ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, n2061}), .clk ( clk ), .rnd ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755]}), .outt ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2062}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2216 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}), .clk ( clk ), .rnd ({Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .outt ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2731}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2690}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, n2068}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2224 ( .ina ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}), .inb ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .clk ( clk ), .rnd ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785]}), .outt ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2642}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2225 ( .ina ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .inb ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .clk ( clk ), .rnd ({Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .outt ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2252}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2228 ( .ina ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2739}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .clk ( clk ), .rnd ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815]}), .outt ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, n2075}) ) ;
    or_HPC1 #(.security_order(4), .pipeline(1)) U2233 ( .ina ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}), .inb ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2723}), .clk ( clk ), .rnd ({Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .outt ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1478, n2081}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2234 ( .ina ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}), .clk ( clk ), .rnd ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845]}), .outt ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, n2080}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2237 ( .ina ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2600}), .inb ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2719}), .clk ( clk ), .rnd ({Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .outt ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, new_AGEMA_signal_1910, n2773}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2239 ( .ina ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .inb ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .clk ( clk ), .rnd ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875]}), .outt ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2083}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2244 ( .ina ({new_AGEMA_signal_17771, new_AGEMA_signal_17769, new_AGEMA_signal_17767, new_AGEMA_signal_17765, new_AGEMA_signal_17763}), .inb ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, n2086}), .clk ( clk ), .rnd ({Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .outt ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, n2562}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2247 ( .ina ({new_AGEMA_signal_17741, new_AGEMA_signal_17739, new_AGEMA_signal_17737, new_AGEMA_signal_17735, new_AGEMA_signal_17733}), .inb ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2661}), .clk ( clk ), .rnd ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905]}), .outt ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, n2087}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2251 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2563}), .inb ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2174}), .clk ( clk ), .rnd ({Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .outt ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, n2156}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2260 ( .ina ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}), .inb ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2401}), .clk ( clk ), .rnd ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935]}), .outt ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2100}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2277 ( .ina ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2739}), .inb ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2298}), .clk ( clk ), .rnd ({Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .outt ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, n2544}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2279 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2356}), .inb ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2118}), .clk ( clk ), .rnd ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965]}), .outt ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2121}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2284 ( .ina ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .inb ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2570}), .clk ( clk ), .rnd ({Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .outt ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1946, n2122}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2286 ( .ina ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .inb ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .clk ( clk ), .rnd ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995]}), .outt ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2811}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2294 ( .ina ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .clk ( clk ), .rnd ({Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .outt ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, n2647}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2297 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .inb ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .clk ( clk ), .rnd ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025]}), .outt ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, n2132}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2304 ( .ina ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2616}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .outt ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1970, n2220}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2305 ( .ina ({new_AGEMA_signal_17711, new_AGEMA_signal_17709, new_AGEMA_signal_17707, new_AGEMA_signal_17705, new_AGEMA_signal_17703}), .inb ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .clk ( clk ), .rnd ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055]}), .outt ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2138}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2312 ( .ina ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .inb ({new_AGEMA_signal_17791, new_AGEMA_signal_17789, new_AGEMA_signal_17787, new_AGEMA_signal_17785, new_AGEMA_signal_17783}), .clk ( clk ), .rnd ({Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .outt ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, n2555}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2322 ( .ina ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .inb ({new_AGEMA_signal_17801, new_AGEMA_signal_17799, new_AGEMA_signal_17797, new_AGEMA_signal_17795, new_AGEMA_signal_17793}), .clk ( clk ), .rnd ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085]}), .outt ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2429}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2328 ( .ina ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}), .inb ({new_AGEMA_signal_17761, new_AGEMA_signal_17759, new_AGEMA_signal_17757, new_AGEMA_signal_17755, new_AGEMA_signal_17753}), .clk ( clk ), .rnd ({Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .outt ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n2162}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2337 ( .ina ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2242}), .clk ( clk ), .rnd ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115]}), .outt ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2545}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2340 ( .ina ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}), .inb ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .clk ( clk ), .rnd ({Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .outt ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, n2178}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2342 ( .ina ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2430}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145]}), .outt ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, n2176}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2343 ( .ina ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2174}), .inb ({new_AGEMA_signal_17771, new_AGEMA_signal_17769, new_AGEMA_signal_17767, new_AGEMA_signal_17765, new_AGEMA_signal_17763}), .clk ( clk ), .rnd ({Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .outt ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, n2175}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2348 ( .ina ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}), .inb ({new_AGEMA_signal_17801, new_AGEMA_signal_17799, new_AGEMA_signal_17797, new_AGEMA_signal_17795, new_AGEMA_signal_17793}), .clk ( clk ), .rnd ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175]}), .outt ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, n2182}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2353 ( .ina ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .inb ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2430}), .clk ( clk ), .rnd ({Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .outt ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2188}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2355 ( .ina ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .inb ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .clk ( clk ), .rnd ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205]}), .outt ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, n2189}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2357 ( .ina ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}), .inb ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}), .clk ( clk ), .rnd ({Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .outt ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, n2446}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2362 ( .ina ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}), .clk ( clk ), .rnd ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235]}), .outt ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2576}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2363 ( .ina ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2609}), .inb ({new_AGEMA_signal_17811, new_AGEMA_signal_17809, new_AGEMA_signal_17807, new_AGEMA_signal_17805, new_AGEMA_signal_17803}), .clk ( clk ), .rnd ({Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .outt ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, n2748}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2654}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2674}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2378 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .inb ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .clk ( clk ), .rnd ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265]}), .outt ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n2213}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2380 ( .ina ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}), .inb ({new_AGEMA_signal_17741, new_AGEMA_signal_17739, new_AGEMA_signal_17737, new_AGEMA_signal_17735, new_AGEMA_signal_17733}), .clk ( clk ), .rnd ({Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .outt ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, n2215}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2384 ( .ina ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2712}), .inb ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2769}), .clk ( clk ), .rnd ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295]}), .outt ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, n2218}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2386 ( .ina ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2298}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .outt ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2219}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2405 ( .ina ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .clk ( clk ), .rnd ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325]}), .outt ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, n2240}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2407 ( .ina ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2709}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2242}), .clk ( clk ), .rnd ({Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .outt ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n2561}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2408 ( .ina ({new_AGEMA_signal_17771, new_AGEMA_signal_17769, new_AGEMA_signal_17767, new_AGEMA_signal_17765, new_AGEMA_signal_17763}), .inb ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .clk ( clk ), .rnd ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355]}), .outt ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, n2243}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2411 ( .ina ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}), .inb ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .clk ( clk ), .rnd ({Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .outt ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, n2245}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2422 ( .ina ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .inb ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2430}), .clk ( clk ), .rnd ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385]}), .outt ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n2540}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2423 ( .ina ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}), .inb ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2640}), .clk ( clk ), .rnd ({Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .outt ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, n2259}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2426 ( .ina ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2261}), .inb ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2661}), .clk ( clk ), .rnd ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415]}), .outt ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, n2262}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2431 ( .ina ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .inb ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n2777}), .clk ( clk ), .rnd ({Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .outt ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2266}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2432 ( .ina ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2772}), .inb ({new_AGEMA_signal_17801, new_AGEMA_signal_17799, new_AGEMA_signal_17797, new_AGEMA_signal_17795, new_AGEMA_signal_17793}), .clk ( clk ), .rnd ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445]}), .outt ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, n2645}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2436 ( .ina ({new_AGEMA_signal_17711, new_AGEMA_signal_17709, new_AGEMA_signal_17707, new_AGEMA_signal_17705, new_AGEMA_signal_17703}), .inb ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .clk ( clk ), .rnd ({Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .outt ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, n2268}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2443 ( .ina ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}), .inb ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .clk ( clk ), .rnd ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475]}), .outt ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, n2278}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2448 ( .ina ({new_AGEMA_signal_17821, new_AGEMA_signal_17819, new_AGEMA_signal_17817, new_AGEMA_signal_17815, new_AGEMA_signal_17813}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .clk ( clk ), .rnd ({Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .outt ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2383}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2455 ( .ina ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .inb ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2570}), .clk ( clk ), .rnd ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505]}), .outt ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2774}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2458 ( .ina ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2823}), .inb ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .clk ( clk ), .rnd ({Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .outt ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, n2287}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2470 ( .ina ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535]}), .outt ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2438}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2471 ( .ina ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2298}), .inb ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .clk ( clk ), .rnd ({Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .outt ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, n2299}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2481 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2313}), .clk ( clk ), .rnd ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565]}), .outt ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, n2371}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2484 ( .ina ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2315}), .inb ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .clk ( clk ), .rnd ({Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .outt ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, n2316}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2486 ( .ina ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, n2624}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2317}), .clk ( clk ), .rnd ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595]}), .outt ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2318}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2492 ( .ina ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .outt ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, n2325}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2494 ( .ina ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625]}), .outt ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2328}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2495 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .inb ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2723}), .clk ( clk ), .rnd ({Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .outt ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, n2327}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2505 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}), .inb ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}), .clk ( clk ), .rnd ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655]}), .outt ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, n2343}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2510 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2563}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .outt ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2344}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(1)) U2512 ( .ina ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2395}), .inb ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, new_AGEMA_signal_1226, n2346}), .clk ( clk ), .rnd ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685]}), .outt ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, n2348}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2513 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .inb ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .clk ( clk ), .rnd ({Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .outt ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n2347}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2520 ( .ina ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}), .inb ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2753}), .clk ( clk ), .rnd ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715]}), .outt ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, new_AGEMA_signal_1582, n2363}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2521 ( .ina ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2809}), .inb ({new_AGEMA_signal_17751, new_AGEMA_signal_17749, new_AGEMA_signal_17747, new_AGEMA_signal_17745, new_AGEMA_signal_17743}), .clk ( clk ), .rnd ({Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .outt ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, n2353}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2524 ( .ina ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .clk ( clk ), .rnd ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745]}), .outt ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, n2355}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2530 ( .ina ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2712}), .inb ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2672}), .clk ( clk ), .rnd ({Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .outt ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2364}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2543 ( .ina ({new_AGEMA_signal_17711, new_AGEMA_signal_17709, new_AGEMA_signal_17707, new_AGEMA_signal_17705, new_AGEMA_signal_17703}), .inb ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2401}), .clk ( clk ), .rnd ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775]}), .outt ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, n2415}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2558 ( .ina ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2395}), .inb ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .clk ( clk ), .rnd ({Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .outt ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2700}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2563 ( .ina ({new_AGEMA_signal_17831, new_AGEMA_signal_17829, new_AGEMA_signal_17827, new_AGEMA_signal_17825, new_AGEMA_signal_17823}), .inb ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2400}), .clk ( clk ), .rnd ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805]}), .outt ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, n2594}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2564 ( .ina ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2401}), .inb ({new_AGEMA_signal_17761, new_AGEMA_signal_17759, new_AGEMA_signal_17757, new_AGEMA_signal_17755, new_AGEMA_signal_17753}), .clk ( clk ), .rnd ({Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .outt ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, n2402}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2585 ( .ina ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2712}), .inb ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2823}), .clk ( clk ), .rnd ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835]}), .outt ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, n2428}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2588 ( .ina ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2430}), .inb ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2570}), .clk ( clk ), .rnd ({Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .outt ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, n2431}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2594 ( .ina ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2437}), .inb ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}), .clk ( clk ), .rnd ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865]}), .outt ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2483}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2599 ( .ina ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2442}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .clk ( clk ), .rnd ({Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .outt ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, n2443}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2606 ( .ina ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .inb ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2609}), .clk ( clk ), .rnd ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895]}), .outt ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, n2693}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2608 ( .ina ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2452}), .inb ({new_AGEMA_signal_17841, new_AGEMA_signal_17839, new_AGEMA_signal_17837, new_AGEMA_signal_17835, new_AGEMA_signal_17833}), .clk ( clk ), .rnd ({Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .outt ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, n2453}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2616 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, n2463}), .clk ( clk ), .rnd ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925]}), .outt ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, n2464}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2620 ( .ina ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2742}), .clk ( clk ), .rnd ({Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .outt ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2468}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2624 ( .ina ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .inb ({new_AGEMA_signal_17751, new_AGEMA_signal_17749, new_AGEMA_signal_17747, new_AGEMA_signal_17745, new_AGEMA_signal_17743}), .clk ( clk ), .rnd ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955]}), .outt ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, new_AGEMA_signal_1618, n2473}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2625 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .inb ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .clk ( clk ), .rnd ({Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .outt ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, n2472}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2628 ( .ina ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2661}), .inb ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n2474}), .clk ( clk ), .rnd ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985]}), .outt ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2475}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2632 ( .ina ({new_AGEMA_signal_17851, new_AGEMA_signal_17849, new_AGEMA_signal_17847, new_AGEMA_signal_17845, new_AGEMA_signal_17843}), .inb ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2828}), .clk ( clk ), .rnd ({Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .outt ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2480}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2638 ( .ina ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2577}), .inb ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}), .clk ( clk ), .rnd ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015]}), .outt ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, n2487}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2641 ( .ina ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2616}), .inb ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}), .clk ( clk ), .rnd ({Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .outt ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, n2488}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2665 ( .ina ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .inb ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2519}), .clk ( clk ), .rnd ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045]}), .outt ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, n2520}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2667 ( .ina ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .inb ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2587}), .clk ( clk ), .rnd ({Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .outt ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, n2521}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2674 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}), .inb ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2595}), .clk ( clk ), .rnd ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075]}), .outt ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, n2531}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2689 ( .ina ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}), .inb ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .clk ( clk ), .rnd ({Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .outt ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, n2553}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2691 ( .ina ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}), .inb ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .clk ( clk ), .rnd ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105]}), .outt ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, n2554}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(1)) U2695 ( .ina ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2559}), .inb ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .clk ( clk ), .rnd ({Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .outt ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2560}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2698 ( .ina ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, new_AGEMA_signal_1334, n2724}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2563}), .clk ( clk ), .rnd ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135]}), .outt ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2564}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2714 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2688}), .inb ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2694}), .clk ( clk ), .rnd ({Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .outt ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2586}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2720 ( .ina ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2595}), .inb ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, n2643}), .clk ( clk ), .rnd ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165]}), .outt ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, n2597}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2721 ( .ina ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2640}), .inb ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .clk ( clk ), .rnd ({Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .outt ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, n2596}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2723 ( .ina ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, new_AGEMA_signal_1334, n2724}), .inb ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .clk ( clk ), .rnd ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195]}), .outt ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2598}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2725 ( .ina ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2635}), .inb ({new_AGEMA_signal_17741, new_AGEMA_signal_17739, new_AGEMA_signal_17737, new_AGEMA_signal_17735, new_AGEMA_signal_17733}), .clk ( clk ), .rnd ({Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .outt ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, new_AGEMA_signal_1258, n2599}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2732 ( .ina ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .inb ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2818}), .clk ( clk ), .rnd ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225]}), .outt ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, n2610}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2734 ( .ina ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .inb ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2611}), .clk ( clk ), .rnd ({Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .outt ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2614}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2735 ( .ina ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2612}), .inb ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .clk ( clk ), .rnd ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255]}), .outt ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, n2613}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2737 ( .ina ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2616}), .inb ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2615}), .clk ( clk ), .rnd ({Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .outt ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2617}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2742 ( .ina ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, n2624}), .inb ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2750}), .clk ( clk ), .rnd ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285]}), .outt ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, new_AGEMA_signal_1654, n2629}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2751 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2641}), .inb ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2640}), .clk ( clk ), .rnd ({Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .outt ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2784}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2757 ( .ina ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, n2785}), .inb ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n2777}), .clk ( clk ), .rnd ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315]}), .outt ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, n2650}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2775 ( .ina ({new_AGEMA_signal_17791, new_AGEMA_signal_17789, new_AGEMA_signal_17787, new_AGEMA_signal_17785, new_AGEMA_signal_17783}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2682}), .clk ( clk ), .rnd ({Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .outt ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, new_AGEMA_signal_1262, n2683}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2789 ( .ina ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2723}), .inb ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2707}), .clk ( clk ), .rnd ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345]}), .outt ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, n2711}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2790 ( .ina ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2709}), .inb ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2708}), .clk ( clk ), .rnd ({Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .outt ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, n2710}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2792 ( .ina ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2713}), .inb ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2712}), .clk ( clk ), .rnd ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375]}), .outt ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2714}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2797 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .inb ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2721}), .clk ( clk ), .rnd ({Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .outt ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, n2722}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2799 ( .ina ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2725}), .inb ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, new_AGEMA_signal_1334, n2724}), .clk ( clk ), .rnd ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405]}), .outt ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, n2726}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2806 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2737}), .inb ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2753}), .clk ( clk ), .rnd ({Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .outt ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, n2738}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2822 ( .ina ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2767}), .inb ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2766}), .clk ( clk ), .rnd ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435]}), .outt ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, n2768}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2828 ( .ina ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2778}), .inb ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n2777}), .clk ( clk ), .rnd ({Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .outt ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, n2782}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2829 ( .ina ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2780}), .inb ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2779}), .clk ( clk ), .rnd ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465]}), .outt ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2781}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2832 ( .ina ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2786}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, n2785}), .clk ( clk ), .rnd ({Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .outt ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, n2787}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2834 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2790}), .inb ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2789}), .clk ( clk ), .rnd ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495]}), .outt ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, n2794}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2835 ( .ina ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, n2792}), .inb ({new_AGEMA_signal_17821, new_AGEMA_signal_17819, new_AGEMA_signal_17817, new_AGEMA_signal_17815, new_AGEMA_signal_17813}), .clk ( clk ), .rnd ({Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .outt ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2793}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2844 ( .ina ({new_AGEMA_signal_17851, new_AGEMA_signal_17849, new_AGEMA_signal_17847, new_AGEMA_signal_17845, new_AGEMA_signal_17843}), .inb ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2809}), .clk ( clk ), .rnd ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525]}), .outt ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, n2812}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2847 ( .ina ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2816}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2815}), .clk ( clk ), .rnd ({Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .outt ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, n2820}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2851 ( .ina ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n2824}), .inb ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2823}), .clk ( clk ), .rnd ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555]}), .outt ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_17852 ), .Q ( new_AGEMA_signal_17853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_17854 ), .Q ( new_AGEMA_signal_17855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_17856 ), .Q ( new_AGEMA_signal_17857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_17858 ), .Q ( new_AGEMA_signal_17859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_17860 ), .Q ( new_AGEMA_signal_17861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_17862 ), .Q ( new_AGEMA_signal_17863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_17864 ), .Q ( new_AGEMA_signal_17865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_17866 ), .Q ( new_AGEMA_signal_17867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_17868 ), .Q ( new_AGEMA_signal_17869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_17870 ), .Q ( new_AGEMA_signal_17871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_17872 ), .Q ( new_AGEMA_signal_17873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_17874 ), .Q ( new_AGEMA_signal_17875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_17876 ), .Q ( new_AGEMA_signal_17877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_17878 ), .Q ( new_AGEMA_signal_17879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_17880 ), .Q ( new_AGEMA_signal_17881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_17882 ), .Q ( new_AGEMA_signal_17883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_17884 ), .Q ( new_AGEMA_signal_17885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_17886 ), .Q ( new_AGEMA_signal_17887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_17888 ), .Q ( new_AGEMA_signal_17889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_17890 ), .Q ( new_AGEMA_signal_17891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_17892 ), .Q ( new_AGEMA_signal_17893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_17894 ), .Q ( new_AGEMA_signal_17895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_17896 ), .Q ( new_AGEMA_signal_17897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_17898 ), .Q ( new_AGEMA_signal_17899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_17900 ), .Q ( new_AGEMA_signal_17901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_17902 ), .Q ( new_AGEMA_signal_17903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_17904 ), .Q ( new_AGEMA_signal_17905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_17906 ), .Q ( new_AGEMA_signal_17907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_17908 ), .Q ( new_AGEMA_signal_17909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_17910 ), .Q ( new_AGEMA_signal_17911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_17912 ), .Q ( new_AGEMA_signal_17913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_17914 ), .Q ( new_AGEMA_signal_17915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_17916 ), .Q ( new_AGEMA_signal_17917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_17918 ), .Q ( new_AGEMA_signal_17919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_17920 ), .Q ( new_AGEMA_signal_17921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_17922 ), .Q ( new_AGEMA_signal_17923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_17924 ), .Q ( new_AGEMA_signal_17925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_17926 ), .Q ( new_AGEMA_signal_17927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_17928 ), .Q ( new_AGEMA_signal_17929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_17930 ), .Q ( new_AGEMA_signal_17931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_17932 ), .Q ( new_AGEMA_signal_17933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_17934 ), .Q ( new_AGEMA_signal_17935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_17936 ), .Q ( new_AGEMA_signal_17937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_17938 ), .Q ( new_AGEMA_signal_17939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_17940 ), .Q ( new_AGEMA_signal_17941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_17942 ), .Q ( new_AGEMA_signal_17943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_17944 ), .Q ( new_AGEMA_signal_17945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_17946 ), .Q ( new_AGEMA_signal_17947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_17948 ), .Q ( new_AGEMA_signal_17949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_17950 ), .Q ( new_AGEMA_signal_17951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_17952 ), .Q ( new_AGEMA_signal_17953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_17954 ), .Q ( new_AGEMA_signal_17955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_17956 ), .Q ( new_AGEMA_signal_17957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_17958 ), .Q ( new_AGEMA_signal_17959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_17960 ), .Q ( new_AGEMA_signal_17961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_17962 ), .Q ( new_AGEMA_signal_17963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_17964 ), .Q ( new_AGEMA_signal_17965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_17966 ), .Q ( new_AGEMA_signal_17967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_17968 ), .Q ( new_AGEMA_signal_17969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_17970 ), .Q ( new_AGEMA_signal_17971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_17972 ), .Q ( new_AGEMA_signal_17973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_17974 ), .Q ( new_AGEMA_signal_17975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_17976 ), .Q ( new_AGEMA_signal_17977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_17978 ), .Q ( new_AGEMA_signal_17979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_17980 ), .Q ( new_AGEMA_signal_17981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_17982 ), .Q ( new_AGEMA_signal_17983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_17984 ), .Q ( new_AGEMA_signal_17985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_17986 ), .Q ( new_AGEMA_signal_17987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_17988 ), .Q ( new_AGEMA_signal_17989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( new_AGEMA_signal_17990 ), .Q ( new_AGEMA_signal_17991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_17992 ), .Q ( new_AGEMA_signal_17993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_17994 ), .Q ( new_AGEMA_signal_17995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_17996 ), .Q ( new_AGEMA_signal_17997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_17998 ), .Q ( new_AGEMA_signal_17999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_18000 ), .Q ( new_AGEMA_signal_18001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_18002 ), .Q ( new_AGEMA_signal_18003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_18004 ), .Q ( new_AGEMA_signal_18005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_18006 ), .Q ( new_AGEMA_signal_18007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_18008 ), .Q ( new_AGEMA_signal_18009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_18010 ), .Q ( new_AGEMA_signal_18011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_18012 ), .Q ( new_AGEMA_signal_18013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_18014 ), .Q ( new_AGEMA_signal_18015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_18016 ), .Q ( new_AGEMA_signal_18017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_18018 ), .Q ( new_AGEMA_signal_18019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_18020 ), .Q ( new_AGEMA_signal_18021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_18022 ), .Q ( new_AGEMA_signal_18023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_18024 ), .Q ( new_AGEMA_signal_18025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_18026 ), .Q ( new_AGEMA_signal_18027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_18028 ), .Q ( new_AGEMA_signal_18029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_18030 ), .Q ( new_AGEMA_signal_18031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_18032 ), .Q ( new_AGEMA_signal_18033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_18034 ), .Q ( new_AGEMA_signal_18035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_18036 ), .Q ( new_AGEMA_signal_18037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_18038 ), .Q ( new_AGEMA_signal_18039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_18040 ), .Q ( new_AGEMA_signal_18041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_18042 ), .Q ( new_AGEMA_signal_18043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_18044 ), .Q ( new_AGEMA_signal_18045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_18046 ), .Q ( new_AGEMA_signal_18047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_18048 ), .Q ( new_AGEMA_signal_18049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_18050 ), .Q ( new_AGEMA_signal_18051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_18052 ), .Q ( new_AGEMA_signal_18053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_18054 ), .Q ( new_AGEMA_signal_18055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_18056 ), .Q ( new_AGEMA_signal_18057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_18058 ), .Q ( new_AGEMA_signal_18059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_18060 ), .Q ( new_AGEMA_signal_18061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_18062 ), .Q ( new_AGEMA_signal_18063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_18064 ), .Q ( new_AGEMA_signal_18065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_18066 ), .Q ( new_AGEMA_signal_18067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_18068 ), .Q ( new_AGEMA_signal_18069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_18070 ), .Q ( new_AGEMA_signal_18071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_18072 ), .Q ( new_AGEMA_signal_18073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_18074 ), .Q ( new_AGEMA_signal_18075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_18076 ), .Q ( new_AGEMA_signal_18077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_18078 ), .Q ( new_AGEMA_signal_18079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_18080 ), .Q ( new_AGEMA_signal_18081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_18082 ), .Q ( new_AGEMA_signal_18083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_18084 ), .Q ( new_AGEMA_signal_18085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_18086 ), .Q ( new_AGEMA_signal_18087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_18088 ), .Q ( new_AGEMA_signal_18089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_18090 ), .Q ( new_AGEMA_signal_18091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_18092 ), .Q ( new_AGEMA_signal_18093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_18094 ), .Q ( new_AGEMA_signal_18095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_18096 ), .Q ( new_AGEMA_signal_18097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_18098 ), .Q ( new_AGEMA_signal_18099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_18100 ), .Q ( new_AGEMA_signal_18101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_18102 ), .Q ( new_AGEMA_signal_18103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_18104 ), .Q ( new_AGEMA_signal_18105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_18106 ), .Q ( new_AGEMA_signal_18107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_18108 ), .Q ( new_AGEMA_signal_18109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_18110 ), .Q ( new_AGEMA_signal_18111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_18112 ), .Q ( new_AGEMA_signal_18113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_18114 ), .Q ( new_AGEMA_signal_18115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_18116 ), .Q ( new_AGEMA_signal_18117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_18118 ), .Q ( new_AGEMA_signal_18119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_18120 ), .Q ( new_AGEMA_signal_18121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_18122 ), .Q ( new_AGEMA_signal_18123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_18124 ), .Q ( new_AGEMA_signal_18125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_18126 ), .Q ( new_AGEMA_signal_18127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_18128 ), .Q ( new_AGEMA_signal_18129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_18130 ), .Q ( new_AGEMA_signal_18131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_18132 ), .Q ( new_AGEMA_signal_18133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_18134 ), .Q ( new_AGEMA_signal_18135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_18136 ), .Q ( new_AGEMA_signal_18137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_18138 ), .Q ( new_AGEMA_signal_18139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_18140 ), .Q ( new_AGEMA_signal_18141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_18142 ), .Q ( new_AGEMA_signal_18143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_18144 ), .Q ( new_AGEMA_signal_18145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_18146 ), .Q ( new_AGEMA_signal_18147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_18148 ), .Q ( new_AGEMA_signal_18149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_18150 ), .Q ( new_AGEMA_signal_18151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_18152 ), .Q ( new_AGEMA_signal_18153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_18154 ), .Q ( new_AGEMA_signal_18155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_18156 ), .Q ( new_AGEMA_signal_18157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_18158 ), .Q ( new_AGEMA_signal_18159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_18160 ), .Q ( new_AGEMA_signal_18161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_18162 ), .Q ( new_AGEMA_signal_18163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_18164 ), .Q ( new_AGEMA_signal_18165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_18166 ), .Q ( new_AGEMA_signal_18167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_18168 ), .Q ( new_AGEMA_signal_18169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_18170 ), .Q ( new_AGEMA_signal_18171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_18172 ), .Q ( new_AGEMA_signal_18173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_18174 ), .Q ( new_AGEMA_signal_18175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_18176 ), .Q ( new_AGEMA_signal_18177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_18178 ), .Q ( new_AGEMA_signal_18179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_18180 ), .Q ( new_AGEMA_signal_18181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_18182 ), .Q ( new_AGEMA_signal_18183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_18184 ), .Q ( new_AGEMA_signal_18185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_18186 ), .Q ( new_AGEMA_signal_18187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_18188 ), .Q ( new_AGEMA_signal_18189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_18190 ), .Q ( new_AGEMA_signal_18191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_18192 ), .Q ( new_AGEMA_signal_18193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_18194 ), .Q ( new_AGEMA_signal_18195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_18196 ), .Q ( new_AGEMA_signal_18197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_18198 ), .Q ( new_AGEMA_signal_18199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_18200 ), .Q ( new_AGEMA_signal_18201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_18202 ), .Q ( new_AGEMA_signal_18203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_18204 ), .Q ( new_AGEMA_signal_18205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_18206 ), .Q ( new_AGEMA_signal_18207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_18208 ), .Q ( new_AGEMA_signal_18209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_18210 ), .Q ( new_AGEMA_signal_18211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_18212 ), .Q ( new_AGEMA_signal_18213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_18214 ), .Q ( new_AGEMA_signal_18215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_18216 ), .Q ( new_AGEMA_signal_18217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_18218 ), .Q ( new_AGEMA_signal_18219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_18220 ), .Q ( new_AGEMA_signal_18221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_18222 ), .Q ( new_AGEMA_signal_18223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_18224 ), .Q ( new_AGEMA_signal_18225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_18226 ), .Q ( new_AGEMA_signal_18227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_18228 ), .Q ( new_AGEMA_signal_18229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_18230 ), .Q ( new_AGEMA_signal_18231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_18232 ), .Q ( new_AGEMA_signal_18233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_18234 ), .Q ( new_AGEMA_signal_18235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_18236 ), .Q ( new_AGEMA_signal_18237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_18238 ), .Q ( new_AGEMA_signal_18239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_18240 ), .Q ( new_AGEMA_signal_18241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_18242 ), .Q ( new_AGEMA_signal_18243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_18244 ), .Q ( new_AGEMA_signal_18245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_18246 ), .Q ( new_AGEMA_signal_18247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_18248 ), .Q ( new_AGEMA_signal_18249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_18250 ), .Q ( new_AGEMA_signal_18251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_18252 ), .Q ( new_AGEMA_signal_18253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_18254 ), .Q ( new_AGEMA_signal_18255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_18256 ), .Q ( new_AGEMA_signal_18257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_18258 ), .Q ( new_AGEMA_signal_18259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_18260 ), .Q ( new_AGEMA_signal_18261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_18262 ), .Q ( new_AGEMA_signal_18263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_18264 ), .Q ( new_AGEMA_signal_18265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_18266 ), .Q ( new_AGEMA_signal_18267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_18268 ), .Q ( new_AGEMA_signal_18269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_18270 ), .Q ( new_AGEMA_signal_18271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_18272 ), .Q ( new_AGEMA_signal_18273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_18274 ), .Q ( new_AGEMA_signal_18275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_18276 ), .Q ( new_AGEMA_signal_18277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_18278 ), .Q ( new_AGEMA_signal_18279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_18280 ), .Q ( new_AGEMA_signal_18281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_18282 ), .Q ( new_AGEMA_signal_18283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_18284 ), .Q ( new_AGEMA_signal_18285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_18286 ), .Q ( new_AGEMA_signal_18287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_18288 ), .Q ( new_AGEMA_signal_18289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_18290 ), .Q ( new_AGEMA_signal_18291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_18292 ), .Q ( new_AGEMA_signal_18293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_18294 ), .Q ( new_AGEMA_signal_18295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_18296 ), .Q ( new_AGEMA_signal_18297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_18298 ), .Q ( new_AGEMA_signal_18299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_18300 ), .Q ( new_AGEMA_signal_18301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_18302 ), .Q ( new_AGEMA_signal_18303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_18304 ), .Q ( new_AGEMA_signal_18305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_18306 ), .Q ( new_AGEMA_signal_18307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_18308 ), .Q ( new_AGEMA_signal_18309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_18310 ), .Q ( new_AGEMA_signal_18311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_18312 ), .Q ( new_AGEMA_signal_18313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_18314 ), .Q ( new_AGEMA_signal_18315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_18316 ), .Q ( new_AGEMA_signal_18317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_18318 ), .Q ( new_AGEMA_signal_18319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_18320 ), .Q ( new_AGEMA_signal_18321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_18322 ), .Q ( new_AGEMA_signal_18323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_18324 ), .Q ( new_AGEMA_signal_18325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_18326 ), .Q ( new_AGEMA_signal_18327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_18328 ), .Q ( new_AGEMA_signal_18329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_18330 ), .Q ( new_AGEMA_signal_18331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_18332 ), .Q ( new_AGEMA_signal_18333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_18334 ), .Q ( new_AGEMA_signal_18335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_18336 ), .Q ( new_AGEMA_signal_18337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_18338 ), .Q ( new_AGEMA_signal_18339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_18340 ), .Q ( new_AGEMA_signal_18341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_18342 ), .Q ( new_AGEMA_signal_18343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_18344 ), .Q ( new_AGEMA_signal_18345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_18346 ), .Q ( new_AGEMA_signal_18347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_18348 ), .Q ( new_AGEMA_signal_18349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_18350 ), .Q ( new_AGEMA_signal_18351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_18352 ), .Q ( new_AGEMA_signal_18353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_18354 ), .Q ( new_AGEMA_signal_18355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_18356 ), .Q ( new_AGEMA_signal_18357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_18358 ), .Q ( new_AGEMA_signal_18359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_18360 ), .Q ( new_AGEMA_signal_18361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_18362 ), .Q ( new_AGEMA_signal_18363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_18364 ), .Q ( new_AGEMA_signal_18365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_18366 ), .Q ( new_AGEMA_signal_18367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_18368 ), .Q ( new_AGEMA_signal_18369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_18370 ), .Q ( new_AGEMA_signal_18371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_18372 ), .Q ( new_AGEMA_signal_18373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_18374 ), .Q ( new_AGEMA_signal_18375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_18376 ), .Q ( new_AGEMA_signal_18377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_18378 ), .Q ( new_AGEMA_signal_18379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_18380 ), .Q ( new_AGEMA_signal_18381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_18382 ), .Q ( new_AGEMA_signal_18383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_18384 ), .Q ( new_AGEMA_signal_18385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_18386 ), .Q ( new_AGEMA_signal_18387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_18388 ), .Q ( new_AGEMA_signal_18389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_18390 ), .Q ( new_AGEMA_signal_18391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_18392 ), .Q ( new_AGEMA_signal_18393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_18394 ), .Q ( new_AGEMA_signal_18395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_18396 ), .Q ( new_AGEMA_signal_18397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_18398 ), .Q ( new_AGEMA_signal_18399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_18400 ), .Q ( new_AGEMA_signal_18401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_18402 ), .Q ( new_AGEMA_signal_18403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_18404 ), .Q ( new_AGEMA_signal_18405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_18406 ), .Q ( new_AGEMA_signal_18407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_18408 ), .Q ( new_AGEMA_signal_18409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_18410 ), .Q ( new_AGEMA_signal_18411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_18412 ), .Q ( new_AGEMA_signal_18413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_18414 ), .Q ( new_AGEMA_signal_18415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_18416 ), .Q ( new_AGEMA_signal_18417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_18418 ), .Q ( new_AGEMA_signal_18419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_18420 ), .Q ( new_AGEMA_signal_18421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_18422 ), .Q ( new_AGEMA_signal_18423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_18424 ), .Q ( new_AGEMA_signal_18425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_18426 ), .Q ( new_AGEMA_signal_18427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_18428 ), .Q ( new_AGEMA_signal_18429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_18430 ), .Q ( new_AGEMA_signal_18431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_18432 ), .Q ( new_AGEMA_signal_18433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_18434 ), .Q ( new_AGEMA_signal_18435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_18436 ), .Q ( new_AGEMA_signal_18437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_18438 ), .Q ( new_AGEMA_signal_18439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_18440 ), .Q ( new_AGEMA_signal_18441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_18442 ), .Q ( new_AGEMA_signal_18443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_18444 ), .Q ( new_AGEMA_signal_18445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_18446 ), .Q ( new_AGEMA_signal_18447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_18448 ), .Q ( new_AGEMA_signal_18449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_18450 ), .Q ( new_AGEMA_signal_18451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_18452 ), .Q ( new_AGEMA_signal_18453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_18454 ), .Q ( new_AGEMA_signal_18455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_18456 ), .Q ( new_AGEMA_signal_18457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_18458 ), .Q ( new_AGEMA_signal_18459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_18460 ), .Q ( new_AGEMA_signal_18461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_18462 ), .Q ( new_AGEMA_signal_18463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_18464 ), .Q ( new_AGEMA_signal_18465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_18466 ), .Q ( new_AGEMA_signal_18467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_18468 ), .Q ( new_AGEMA_signal_18469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_18470 ), .Q ( new_AGEMA_signal_18471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_18472 ), .Q ( new_AGEMA_signal_18473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_18474 ), .Q ( new_AGEMA_signal_18475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_18476 ), .Q ( new_AGEMA_signal_18477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_18478 ), .Q ( new_AGEMA_signal_18479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_18480 ), .Q ( new_AGEMA_signal_18481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_18482 ), .Q ( new_AGEMA_signal_18483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_18484 ), .Q ( new_AGEMA_signal_18485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_18486 ), .Q ( new_AGEMA_signal_18487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_18488 ), .Q ( new_AGEMA_signal_18489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_18490 ), .Q ( new_AGEMA_signal_18491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_18492 ), .Q ( new_AGEMA_signal_18493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_18494 ), .Q ( new_AGEMA_signal_18495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_18496 ), .Q ( new_AGEMA_signal_18497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_18498 ), .Q ( new_AGEMA_signal_18499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_18500 ), .Q ( new_AGEMA_signal_18501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_18502 ), .Q ( new_AGEMA_signal_18503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_18504 ), .Q ( new_AGEMA_signal_18505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_18506 ), .Q ( new_AGEMA_signal_18507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_18508 ), .Q ( new_AGEMA_signal_18509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_18510 ), .Q ( new_AGEMA_signal_18511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_18512 ), .Q ( new_AGEMA_signal_18513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_18514 ), .Q ( new_AGEMA_signal_18515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_18516 ), .Q ( new_AGEMA_signal_18517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_18518 ), .Q ( new_AGEMA_signal_18519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_18520 ), .Q ( new_AGEMA_signal_18521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_18522 ), .Q ( new_AGEMA_signal_18523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_18524 ), .Q ( new_AGEMA_signal_18525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_18526 ), .Q ( new_AGEMA_signal_18527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_18528 ), .Q ( new_AGEMA_signal_18529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_18530 ), .Q ( new_AGEMA_signal_18531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_18552 ), .Q ( new_AGEMA_signal_18553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_18556 ), .Q ( new_AGEMA_signal_18557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_18560 ), .Q ( new_AGEMA_signal_18561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_18564 ), .Q ( new_AGEMA_signal_18565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_18568 ), .Q ( new_AGEMA_signal_18569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_18682 ), .Q ( new_AGEMA_signal_18683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_18686 ), .Q ( new_AGEMA_signal_18687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_18690 ), .Q ( new_AGEMA_signal_18691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_18694 ), .Q ( new_AGEMA_signal_18695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_18698 ), .Q ( new_AGEMA_signal_18699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_18772 ), .Q ( new_AGEMA_signal_18773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_18776 ), .Q ( new_AGEMA_signal_18777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_18780 ), .Q ( new_AGEMA_signal_18781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_18784 ), .Q ( new_AGEMA_signal_18785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_18788 ), .Q ( new_AGEMA_signal_18789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_18842 ), .Q ( new_AGEMA_signal_18843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_18846 ), .Q ( new_AGEMA_signal_18847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_18850 ), .Q ( new_AGEMA_signal_18851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_18854 ), .Q ( new_AGEMA_signal_18855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_18858 ), .Q ( new_AGEMA_signal_18859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_18892 ), .Q ( new_AGEMA_signal_18893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_18896 ), .Q ( new_AGEMA_signal_18897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_18900 ), .Q ( new_AGEMA_signal_18901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_18904 ), .Q ( new_AGEMA_signal_18905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_18908 ), .Q ( new_AGEMA_signal_18909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_18942 ), .Q ( new_AGEMA_signal_18943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_18946 ), .Q ( new_AGEMA_signal_18947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_18950 ), .Q ( new_AGEMA_signal_18951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_18954 ), .Q ( new_AGEMA_signal_18955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_18958 ), .Q ( new_AGEMA_signal_18959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_19134 ), .Q ( new_AGEMA_signal_19135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_19140 ), .Q ( new_AGEMA_signal_19141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_19146 ), .Q ( new_AGEMA_signal_19147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_19152 ), .Q ( new_AGEMA_signal_19153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_19158 ), .Q ( new_AGEMA_signal_19159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_19192 ), .Q ( new_AGEMA_signal_19193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_19196 ), .Q ( new_AGEMA_signal_19197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_19200 ), .Q ( new_AGEMA_signal_19201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_19204 ), .Q ( new_AGEMA_signal_19205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_19208 ), .Q ( new_AGEMA_signal_19209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_19242 ), .Q ( new_AGEMA_signal_19243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_19246 ), .Q ( new_AGEMA_signal_19247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_19250 ), .Q ( new_AGEMA_signal_19251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_19254 ), .Q ( new_AGEMA_signal_19255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_19258 ), .Q ( new_AGEMA_signal_19259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_19332 ), .Q ( new_AGEMA_signal_19333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_19336 ), .Q ( new_AGEMA_signal_19337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_19340 ), .Q ( new_AGEMA_signal_19341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_19344 ), .Q ( new_AGEMA_signal_19345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_19348 ), .Q ( new_AGEMA_signal_19349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_19372 ), .Q ( new_AGEMA_signal_19373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_19376 ), .Q ( new_AGEMA_signal_19377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_19380 ), .Q ( new_AGEMA_signal_19381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_19384 ), .Q ( new_AGEMA_signal_19385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C ( clk ), .D ( new_AGEMA_signal_19388 ), .Q ( new_AGEMA_signal_19389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C ( clk ), .D ( new_AGEMA_signal_19742 ), .Q ( new_AGEMA_signal_19743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C ( clk ), .D ( new_AGEMA_signal_19748 ), .Q ( new_AGEMA_signal_19749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C ( clk ), .D ( new_AGEMA_signal_19754 ), .Q ( new_AGEMA_signal_19755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C ( clk ), .D ( new_AGEMA_signal_19760 ), .Q ( new_AGEMA_signal_19761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C ( clk ), .D ( new_AGEMA_signal_19766 ), .Q ( new_AGEMA_signal_19767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C ( clk ), .D ( new_AGEMA_signal_19872 ), .Q ( new_AGEMA_signal_19873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C ( clk ), .D ( new_AGEMA_signal_19878 ), .Q ( new_AGEMA_signal_19879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C ( clk ), .D ( new_AGEMA_signal_19884 ), .Q ( new_AGEMA_signal_19885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C ( clk ), .D ( new_AGEMA_signal_19890 ), .Q ( new_AGEMA_signal_19891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C ( clk ), .D ( new_AGEMA_signal_19896 ), .Q ( new_AGEMA_signal_19897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C ( clk ), .D ( new_AGEMA_signal_20452 ), .Q ( new_AGEMA_signal_20453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C ( clk ), .D ( new_AGEMA_signal_20460 ), .Q ( new_AGEMA_signal_20461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C ( clk ), .D ( new_AGEMA_signal_20468 ), .Q ( new_AGEMA_signal_20469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C ( clk ), .D ( new_AGEMA_signal_20476 ), .Q ( new_AGEMA_signal_20477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C ( clk ), .D ( new_AGEMA_signal_20484 ), .Q ( new_AGEMA_signal_20485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C ( clk ), .D ( new_AGEMA_signal_20502 ), .Q ( new_AGEMA_signal_20503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C ( clk ), .D ( new_AGEMA_signal_20510 ), .Q ( new_AGEMA_signal_20511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C ( clk ), .D ( new_AGEMA_signal_20518 ), .Q ( new_AGEMA_signal_20519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C ( clk ), .D ( new_AGEMA_signal_20526 ), .Q ( new_AGEMA_signal_20527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C ( clk ), .D ( new_AGEMA_signal_20534 ), .Q ( new_AGEMA_signal_20535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C ( clk ), .D ( new_AGEMA_signal_20882 ), .Q ( new_AGEMA_signal_20883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C ( clk ), .D ( new_AGEMA_signal_20890 ), .Q ( new_AGEMA_signal_20891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C ( clk ), .D ( new_AGEMA_signal_20898 ), .Q ( new_AGEMA_signal_20899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C ( clk ), .D ( new_AGEMA_signal_20906 ), .Q ( new_AGEMA_signal_20907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C ( clk ), .D ( new_AGEMA_signal_20914 ), .Q ( new_AGEMA_signal_20915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C ( clk ), .D ( new_AGEMA_signal_21312 ), .Q ( new_AGEMA_signal_21313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C ( clk ), .D ( new_AGEMA_signal_21320 ), .Q ( new_AGEMA_signal_21321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C ( clk ), .D ( new_AGEMA_signal_21328 ), .Q ( new_AGEMA_signal_21329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C ( clk ), .D ( new_AGEMA_signal_21336 ), .Q ( new_AGEMA_signal_21337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C ( clk ), .D ( new_AGEMA_signal_21344 ), .Q ( new_AGEMA_signal_21345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C ( clk ), .D ( new_AGEMA_signal_21462 ), .Q ( new_AGEMA_signal_21463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C ( clk ), .D ( new_AGEMA_signal_21470 ), .Q ( new_AGEMA_signal_21471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C ( clk ), .D ( new_AGEMA_signal_21478 ), .Q ( new_AGEMA_signal_21479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C ( clk ), .D ( new_AGEMA_signal_21486 ), .Q ( new_AGEMA_signal_21487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C ( clk ), .D ( new_AGEMA_signal_21494 ), .Q ( new_AGEMA_signal_21495 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_18532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_1294 ), .Q ( new_AGEMA_signal_18534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( new_AGEMA_signal_1295 ), .Q ( new_AGEMA_signal_18536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_1296 ), .Q ( new_AGEMA_signal_18538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_18540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_18542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_1702 ), .Q ( new_AGEMA_signal_18544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( new_AGEMA_signal_1703 ), .Q ( new_AGEMA_signal_18546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( new_AGEMA_signal_1704 ), .Q ( new_AGEMA_signal_18548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( new_AGEMA_signal_1705 ), .Q ( new_AGEMA_signal_18550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( new_AGEMA_signal_18553 ), .Q ( new_AGEMA_signal_18554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( new_AGEMA_signal_18557 ), .Q ( new_AGEMA_signal_18558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( new_AGEMA_signal_18561 ), .Q ( new_AGEMA_signal_18562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( new_AGEMA_signal_18565 ), .Q ( new_AGEMA_signal_18566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( new_AGEMA_signal_18569 ), .Q ( new_AGEMA_signal_18570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( new_AGEMA_signal_17933 ), .Q ( new_AGEMA_signal_18572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( new_AGEMA_signal_17935 ), .Q ( new_AGEMA_signal_18574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( new_AGEMA_signal_17937 ), .Q ( new_AGEMA_signal_18576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( new_AGEMA_signal_17939 ), .Q ( new_AGEMA_signal_18578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_17941 ), .Q ( new_AGEMA_signal_18580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( new_AGEMA_signal_17903 ), .Q ( new_AGEMA_signal_18582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( new_AGEMA_signal_17905 ), .Q ( new_AGEMA_signal_18584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( new_AGEMA_signal_17907 ), .Q ( new_AGEMA_signal_18586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_17909 ), .Q ( new_AGEMA_signal_18588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( new_AGEMA_signal_17911 ), .Q ( new_AGEMA_signal_18590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_18592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( new_AGEMA_signal_1170 ), .Q ( new_AGEMA_signal_18594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( new_AGEMA_signal_1171 ), .Q ( new_AGEMA_signal_18596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( new_AGEMA_signal_1172 ), .Q ( new_AGEMA_signal_18598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_1173 ), .Q ( new_AGEMA_signal_18600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_18602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_1382 ), .Q ( new_AGEMA_signal_18604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( new_AGEMA_signal_1383 ), .Q ( new_AGEMA_signal_18606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_1384 ), .Q ( new_AGEMA_signal_18608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( new_AGEMA_signal_1385 ), .Q ( new_AGEMA_signal_18610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_18612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( new_AGEMA_signal_1762 ), .Q ( new_AGEMA_signal_18614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_18616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_1764 ), .Q ( new_AGEMA_signal_18618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( new_AGEMA_signal_1765 ), .Q ( new_AGEMA_signal_18620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_18622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( new_AGEMA_signal_1778 ), .Q ( new_AGEMA_signal_18624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( new_AGEMA_signal_1779 ), .Q ( new_AGEMA_signal_18626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_1780 ), .Q ( new_AGEMA_signal_18628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_18630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_18632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_1418 ), .Q ( new_AGEMA_signal_18634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_1419 ), .Q ( new_AGEMA_signal_18636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( new_AGEMA_signal_1420 ), .Q ( new_AGEMA_signal_18638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_1421 ), .Q ( new_AGEMA_signal_18640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_18642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( new_AGEMA_signal_1786 ), .Q ( new_AGEMA_signal_18644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( new_AGEMA_signal_1787 ), .Q ( new_AGEMA_signal_18646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_1788 ), .Q ( new_AGEMA_signal_18648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( new_AGEMA_signal_1789 ), .Q ( new_AGEMA_signal_18650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_18652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( new_AGEMA_signal_1430 ), .Q ( new_AGEMA_signal_18654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( new_AGEMA_signal_1431 ), .Q ( new_AGEMA_signal_18656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( new_AGEMA_signal_1432 ), .Q ( new_AGEMA_signal_18658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( new_AGEMA_signal_1433 ), .Q ( new_AGEMA_signal_18660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_18662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( new_AGEMA_signal_1802 ), .Q ( new_AGEMA_signal_18664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( new_AGEMA_signal_1803 ), .Q ( new_AGEMA_signal_18666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( new_AGEMA_signal_1804 ), .Q ( new_AGEMA_signal_18668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( new_AGEMA_signal_1805 ), .Q ( new_AGEMA_signal_18670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( new_AGEMA_signal_18203 ), .Q ( new_AGEMA_signal_18672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( new_AGEMA_signal_18205 ), .Q ( new_AGEMA_signal_18674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_18207 ), .Q ( new_AGEMA_signal_18676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( new_AGEMA_signal_18209 ), .Q ( new_AGEMA_signal_18678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( new_AGEMA_signal_18211 ), .Q ( new_AGEMA_signal_18680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_18683 ), .Q ( new_AGEMA_signal_18684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( new_AGEMA_signal_18687 ), .Q ( new_AGEMA_signal_18688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( new_AGEMA_signal_18691 ), .Q ( new_AGEMA_signal_18692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( new_AGEMA_signal_18695 ), .Q ( new_AGEMA_signal_18696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_18699 ), .Q ( new_AGEMA_signal_18700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_18702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_1846 ), .Q ( new_AGEMA_signal_18704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( new_AGEMA_signal_1847 ), .Q ( new_AGEMA_signal_18706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_1848 ), .Q ( new_AGEMA_signal_18708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( new_AGEMA_signal_1849 ), .Q ( new_AGEMA_signal_18710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_18712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( new_AGEMA_signal_1466 ), .Q ( new_AGEMA_signal_18714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( new_AGEMA_signal_1467 ), .Q ( new_AGEMA_signal_18716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( new_AGEMA_signal_1468 ), .Q ( new_AGEMA_signal_18718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( new_AGEMA_signal_1469 ), .Q ( new_AGEMA_signal_18720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_18722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_1862 ), .Q ( new_AGEMA_signal_18724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( new_AGEMA_signal_1863 ), .Q ( new_AGEMA_signal_18726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( new_AGEMA_signal_1864 ), .Q ( new_AGEMA_signal_18728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_18730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_18732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( new_AGEMA_signal_1866 ), .Q ( new_AGEMA_signal_18734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_1867 ), .Q ( new_AGEMA_signal_18736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( new_AGEMA_signal_1868 ), .Q ( new_AGEMA_signal_18738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_1869 ), .Q ( new_AGEMA_signal_18740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( new_AGEMA_signal_17853 ), .Q ( new_AGEMA_signal_18742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_17855 ), .Q ( new_AGEMA_signal_18744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( new_AGEMA_signal_17857 ), .Q ( new_AGEMA_signal_18746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_17859 ), .Q ( new_AGEMA_signal_18748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( new_AGEMA_signal_17861 ), .Q ( new_AGEMA_signal_18750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_18752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( new_AGEMA_signal_1774 ), .Q ( new_AGEMA_signal_18754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_1775 ), .Q ( new_AGEMA_signal_18756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( new_AGEMA_signal_1776 ), .Q ( new_AGEMA_signal_18758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_1777 ), .Q ( new_AGEMA_signal_18760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_18762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_1470 ), .Q ( new_AGEMA_signal_18764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_1471 ), .Q ( new_AGEMA_signal_18766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_1472 ), .Q ( new_AGEMA_signal_18768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( new_AGEMA_signal_1473 ), .Q ( new_AGEMA_signal_18770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( new_AGEMA_signal_18773 ), .Q ( new_AGEMA_signal_18774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( new_AGEMA_signal_18777 ), .Q ( new_AGEMA_signal_18778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( new_AGEMA_signal_18781 ), .Q ( new_AGEMA_signal_18782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_18785 ), .Q ( new_AGEMA_signal_18786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( new_AGEMA_signal_18789 ), .Q ( new_AGEMA_signal_18790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_18792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( new_AGEMA_signal_1910 ), .Q ( new_AGEMA_signal_18794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_1911 ), .Q ( new_AGEMA_signal_18796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( new_AGEMA_signal_1912 ), .Q ( new_AGEMA_signal_18798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_1913 ), .Q ( new_AGEMA_signal_18800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_18802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_1366 ), .Q ( new_AGEMA_signal_18804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( new_AGEMA_signal_1367 ), .Q ( new_AGEMA_signal_18806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_18808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( new_AGEMA_signal_1369 ), .Q ( new_AGEMA_signal_18810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( new_AGEMA_signal_18053 ), .Q ( new_AGEMA_signal_18812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_18055 ), .Q ( new_AGEMA_signal_18814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_18057 ), .Q ( new_AGEMA_signal_18816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( new_AGEMA_signal_18059 ), .Q ( new_AGEMA_signal_18818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_18061 ), .Q ( new_AGEMA_signal_18820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_18822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( new_AGEMA_signal_1310 ), .Q ( new_AGEMA_signal_18824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_1311 ), .Q ( new_AGEMA_signal_18826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_1312 ), .Q ( new_AGEMA_signal_18828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( new_AGEMA_signal_1313 ), .Q ( new_AGEMA_signal_18830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_18832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_1850 ), .Q ( new_AGEMA_signal_18834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_1851 ), .Q ( new_AGEMA_signal_18836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( new_AGEMA_signal_1852 ), .Q ( new_AGEMA_signal_18838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_18840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_18843 ), .Q ( new_AGEMA_signal_18844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( new_AGEMA_signal_18847 ), .Q ( new_AGEMA_signal_18848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( new_AGEMA_signal_18851 ), .Q ( new_AGEMA_signal_18852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_18855 ), .Q ( new_AGEMA_signal_18856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_18859 ), .Q ( new_AGEMA_signal_18860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_18283 ), .Q ( new_AGEMA_signal_18862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( new_AGEMA_signal_18285 ), .Q ( new_AGEMA_signal_18864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( new_AGEMA_signal_18287 ), .Q ( new_AGEMA_signal_18866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( new_AGEMA_signal_18289 ), .Q ( new_AGEMA_signal_18868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( new_AGEMA_signal_18291 ), .Q ( new_AGEMA_signal_18870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_18103 ), .Q ( new_AGEMA_signal_18872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_18105 ), .Q ( new_AGEMA_signal_18874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_18107 ), .Q ( new_AGEMA_signal_18876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( new_AGEMA_signal_18109 ), .Q ( new_AGEMA_signal_18878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_18111 ), .Q ( new_AGEMA_signal_18880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_18143 ), .Q ( new_AGEMA_signal_18882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( new_AGEMA_signal_18145 ), .Q ( new_AGEMA_signal_18884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( new_AGEMA_signal_18147 ), .Q ( new_AGEMA_signal_18886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_18149 ), .Q ( new_AGEMA_signal_18888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( new_AGEMA_signal_18151 ), .Q ( new_AGEMA_signal_18890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_18893 ), .Q ( new_AGEMA_signal_18894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( new_AGEMA_signal_18897 ), .Q ( new_AGEMA_signal_18898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( new_AGEMA_signal_18901 ), .Q ( new_AGEMA_signal_18902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_18905 ), .Q ( new_AGEMA_signal_18906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( new_AGEMA_signal_18909 ), .Q ( new_AGEMA_signal_18910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_18483 ), .Q ( new_AGEMA_signal_18912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_18485 ), .Q ( new_AGEMA_signal_18914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( new_AGEMA_signal_18487 ), .Q ( new_AGEMA_signal_18916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( new_AGEMA_signal_18489 ), .Q ( new_AGEMA_signal_18918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_18491 ), .Q ( new_AGEMA_signal_18920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_18922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_18924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( new_AGEMA_signal_1483 ), .Q ( new_AGEMA_signal_18926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_1484 ), .Q ( new_AGEMA_signal_18928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( new_AGEMA_signal_1485 ), .Q ( new_AGEMA_signal_18930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_18932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( new_AGEMA_signal_1514 ), .Q ( new_AGEMA_signal_18934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( new_AGEMA_signal_1515 ), .Q ( new_AGEMA_signal_18936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_18938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_1517 ), .Q ( new_AGEMA_signal_18940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_18943 ), .Q ( new_AGEMA_signal_18944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_18947 ), .Q ( new_AGEMA_signal_18948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( new_AGEMA_signal_18951 ), .Q ( new_AGEMA_signal_18952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( new_AGEMA_signal_18955 ), .Q ( new_AGEMA_signal_18956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_18959 ), .Q ( new_AGEMA_signal_18960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_18962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_18964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( new_AGEMA_signal_1759 ), .Q ( new_AGEMA_signal_18966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_18968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_1761 ), .Q ( new_AGEMA_signal_18970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_18972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( new_AGEMA_signal_2058 ), .Q ( new_AGEMA_signal_18974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_2059 ), .Q ( new_AGEMA_signal_18976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( new_AGEMA_signal_2060 ), .Q ( new_AGEMA_signal_18978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( new_AGEMA_signal_2061 ), .Q ( new_AGEMA_signal_18980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_18982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( new_AGEMA_signal_1542 ), .Q ( new_AGEMA_signal_18984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( new_AGEMA_signal_1543 ), .Q ( new_AGEMA_signal_18986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( new_AGEMA_signal_1544 ), .Q ( new_AGEMA_signal_18988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( new_AGEMA_signal_1545 ), .Q ( new_AGEMA_signal_18990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_18992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_2074 ), .Q ( new_AGEMA_signal_18994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_2075 ), .Q ( new_AGEMA_signal_18996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( new_AGEMA_signal_2076 ), .Q ( new_AGEMA_signal_18998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( new_AGEMA_signal_2077 ), .Q ( new_AGEMA_signal_19000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( new_AGEMA_signal_18263 ), .Q ( new_AGEMA_signal_19002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( new_AGEMA_signal_18265 ), .Q ( new_AGEMA_signal_19004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( new_AGEMA_signal_18267 ), .Q ( new_AGEMA_signal_19006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_18269 ), .Q ( new_AGEMA_signal_19008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( new_AGEMA_signal_18271 ), .Q ( new_AGEMA_signal_19010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_18373 ), .Q ( new_AGEMA_signal_19012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( new_AGEMA_signal_18375 ), .Q ( new_AGEMA_signal_19014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_18377 ), .Q ( new_AGEMA_signal_19016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( new_AGEMA_signal_18379 ), .Q ( new_AGEMA_signal_19018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_18381 ), .Q ( new_AGEMA_signal_19020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( new_AGEMA_signal_18033 ), .Q ( new_AGEMA_signal_19022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( new_AGEMA_signal_18035 ), .Q ( new_AGEMA_signal_19024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( new_AGEMA_signal_18037 ), .Q ( new_AGEMA_signal_19026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( new_AGEMA_signal_18039 ), .Q ( new_AGEMA_signal_19028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( new_AGEMA_signal_18041 ), .Q ( new_AGEMA_signal_19030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( new_AGEMA_signal_18013 ), .Q ( new_AGEMA_signal_19032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( new_AGEMA_signal_18015 ), .Q ( new_AGEMA_signal_19034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_18017 ), .Q ( new_AGEMA_signal_19036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_18019 ), .Q ( new_AGEMA_signal_19038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( new_AGEMA_signal_18021 ), .Q ( new_AGEMA_signal_19040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_19042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( new_AGEMA_signal_1566 ), .Q ( new_AGEMA_signal_19044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( new_AGEMA_signal_1567 ), .Q ( new_AGEMA_signal_19046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_1568 ), .Q ( new_AGEMA_signal_19048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_1569 ), .Q ( new_AGEMA_signal_19050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_19052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( new_AGEMA_signal_2114 ), .Q ( new_AGEMA_signal_19054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_2115 ), .Q ( new_AGEMA_signal_19056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( new_AGEMA_signal_2116 ), .Q ( new_AGEMA_signal_19058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_2117 ), .Q ( new_AGEMA_signal_19060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_19062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( new_AGEMA_signal_1362 ), .Q ( new_AGEMA_signal_19064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_1363 ), .Q ( new_AGEMA_signal_19066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_1364 ), .Q ( new_AGEMA_signal_19068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( new_AGEMA_signal_1365 ), .Q ( new_AGEMA_signal_19070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_18463 ), .Q ( new_AGEMA_signal_19072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_18465 ), .Q ( new_AGEMA_signal_19074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_18467 ), .Q ( new_AGEMA_signal_19076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( new_AGEMA_signal_18469 ), .Q ( new_AGEMA_signal_19078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_18471 ), .Q ( new_AGEMA_signal_19080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_18503 ), .Q ( new_AGEMA_signal_19082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_18505 ), .Q ( new_AGEMA_signal_19084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( new_AGEMA_signal_18507 ), .Q ( new_AGEMA_signal_19086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_18509 ), .Q ( new_AGEMA_signal_19088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_18511 ), .Q ( new_AGEMA_signal_19090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_18123 ), .Q ( new_AGEMA_signal_19092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( new_AGEMA_signal_18125 ), .Q ( new_AGEMA_signal_19094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_18127 ), .Q ( new_AGEMA_signal_19096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_18129 ), .Q ( new_AGEMA_signal_19098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( new_AGEMA_signal_18131 ), .Q ( new_AGEMA_signal_19100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( new_AGEMA_signal_17873 ), .Q ( new_AGEMA_signal_19102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_17875 ), .Q ( new_AGEMA_signal_19104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_17877 ), .Q ( new_AGEMA_signal_19106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( new_AGEMA_signal_17879 ), .Q ( new_AGEMA_signal_19108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( new_AGEMA_signal_17881 ), .Q ( new_AGEMA_signal_19110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_19112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_19114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( new_AGEMA_signal_1767 ), .Q ( new_AGEMA_signal_19116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_1768 ), .Q ( new_AGEMA_signal_19118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( new_AGEMA_signal_1769 ), .Q ( new_AGEMA_signal_19120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_19122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( new_AGEMA_signal_2198 ), .Q ( new_AGEMA_signal_19124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_2199 ), .Q ( new_AGEMA_signal_19126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_2200 ), .Q ( new_AGEMA_signal_19128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_2201 ), .Q ( new_AGEMA_signal_19130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( new_AGEMA_signal_19135 ), .Q ( new_AGEMA_signal_19136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( new_AGEMA_signal_19141 ), .Q ( new_AGEMA_signal_19142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( new_AGEMA_signal_19147 ), .Q ( new_AGEMA_signal_19148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( new_AGEMA_signal_19153 ), .Q ( new_AGEMA_signal_19154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( new_AGEMA_signal_19159 ), .Q ( new_AGEMA_signal_19160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_19162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_1606 ), .Q ( new_AGEMA_signal_19164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( new_AGEMA_signal_1607 ), .Q ( new_AGEMA_signal_19166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_19168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( new_AGEMA_signal_1609 ), .Q ( new_AGEMA_signal_19170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_19172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( new_AGEMA_signal_1626 ), .Q ( new_AGEMA_signal_19174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_1627 ), .Q ( new_AGEMA_signal_19176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_1628 ), .Q ( new_AGEMA_signal_19178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_1629 ), .Q ( new_AGEMA_signal_19180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_19182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( new_AGEMA_signal_2230 ), .Q ( new_AGEMA_signal_19184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_2231 ), .Q ( new_AGEMA_signal_19186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( new_AGEMA_signal_2232 ), .Q ( new_AGEMA_signal_19188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( new_AGEMA_signal_2233 ), .Q ( new_AGEMA_signal_19190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( new_AGEMA_signal_19193 ), .Q ( new_AGEMA_signal_19194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( new_AGEMA_signal_19197 ), .Q ( new_AGEMA_signal_19198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( new_AGEMA_signal_19201 ), .Q ( new_AGEMA_signal_19202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( new_AGEMA_signal_19205 ), .Q ( new_AGEMA_signal_19206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( new_AGEMA_signal_19209 ), .Q ( new_AGEMA_signal_19210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_18223 ), .Q ( new_AGEMA_signal_19212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( new_AGEMA_signal_18225 ), .Q ( new_AGEMA_signal_19214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_18227 ), .Q ( new_AGEMA_signal_19216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_18229 ), .Q ( new_AGEMA_signal_19218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( new_AGEMA_signal_18231 ), .Q ( new_AGEMA_signal_19220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( new_AGEMA_signal_18243 ), .Q ( new_AGEMA_signal_19222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_18245 ), .Q ( new_AGEMA_signal_19224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( new_AGEMA_signal_18247 ), .Q ( new_AGEMA_signal_19226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_18249 ), .Q ( new_AGEMA_signal_19228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_18251 ), .Q ( new_AGEMA_signal_19230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_19232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( new_AGEMA_signal_2274 ), .Q ( new_AGEMA_signal_19234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_2275 ), .Q ( new_AGEMA_signal_19236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( new_AGEMA_signal_2276 ), .Q ( new_AGEMA_signal_19238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_2277 ), .Q ( new_AGEMA_signal_19240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_19243 ), .Q ( new_AGEMA_signal_19244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_19247 ), .Q ( new_AGEMA_signal_19248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_19251 ), .Q ( new_AGEMA_signal_19252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( new_AGEMA_signal_19255 ), .Q ( new_AGEMA_signal_19256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_19259 ), .Q ( new_AGEMA_signal_19260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_19262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_1650 ), .Q ( new_AGEMA_signal_19264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_1651 ), .Q ( new_AGEMA_signal_19266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( new_AGEMA_signal_1652 ), .Q ( new_AGEMA_signal_19268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_19270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_19272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( new_AGEMA_signal_1498 ), .Q ( new_AGEMA_signal_19274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_1499 ), .Q ( new_AGEMA_signal_19276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( new_AGEMA_signal_1500 ), .Q ( new_AGEMA_signal_19278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( new_AGEMA_signal_1501 ), .Q ( new_AGEMA_signal_19280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_19282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_2674 ), .Q ( new_AGEMA_signal_19284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( new_AGEMA_signal_2675 ), .Q ( new_AGEMA_signal_19286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_2676 ), .Q ( new_AGEMA_signal_19288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( new_AGEMA_signal_2677 ), .Q ( new_AGEMA_signal_19290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_19292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( new_AGEMA_signal_1262 ), .Q ( new_AGEMA_signal_19294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_1263 ), .Q ( new_AGEMA_signal_19296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( new_AGEMA_signal_1264 ), .Q ( new_AGEMA_signal_19298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_1265 ), .Q ( new_AGEMA_signal_19300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_19302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_1662 ), .Q ( new_AGEMA_signal_19304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_1663 ), .Q ( new_AGEMA_signal_19306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_1664 ), .Q ( new_AGEMA_signal_19308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( new_AGEMA_signal_1665 ), .Q ( new_AGEMA_signal_19310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_19312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( new_AGEMA_signal_2362 ), .Q ( new_AGEMA_signal_19314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( new_AGEMA_signal_2363 ), .Q ( new_AGEMA_signal_19316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_2364 ), .Q ( new_AGEMA_signal_19318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_2365 ), .Q ( new_AGEMA_signal_19320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_19322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( new_AGEMA_signal_1706 ), .Q ( new_AGEMA_signal_19324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_1707 ), .Q ( new_AGEMA_signal_19326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_1708 ), .Q ( new_AGEMA_signal_19328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_1709 ), .Q ( new_AGEMA_signal_19330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( new_AGEMA_signal_19333 ), .Q ( new_AGEMA_signal_19334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( new_AGEMA_signal_19337 ), .Q ( new_AGEMA_signal_19338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_19341 ), .Q ( new_AGEMA_signal_19342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( new_AGEMA_signal_19345 ), .Q ( new_AGEMA_signal_19346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( new_AGEMA_signal_19349 ), .Q ( new_AGEMA_signal_19350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_19352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( new_AGEMA_signal_1710 ), .Q ( new_AGEMA_signal_19354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_1711 ), .Q ( new_AGEMA_signal_19356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( new_AGEMA_signal_1712 ), .Q ( new_AGEMA_signal_19358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_1713 ), .Q ( new_AGEMA_signal_19360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_19362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_2322 ), .Q ( new_AGEMA_signal_19364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_2323 ), .Q ( new_AGEMA_signal_19366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_2324 ), .Q ( new_AGEMA_signal_19368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( new_AGEMA_signal_2325 ), .Q ( new_AGEMA_signal_19370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_19373 ), .Q ( new_AGEMA_signal_19374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( new_AGEMA_signal_19377 ), .Q ( new_AGEMA_signal_19378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( new_AGEMA_signal_19381 ), .Q ( new_AGEMA_signal_19382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C ( clk ), .D ( new_AGEMA_signal_19385 ), .Q ( new_AGEMA_signal_19386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C ( clk ), .D ( new_AGEMA_signal_19389 ), .Q ( new_AGEMA_signal_19390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_19392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C ( clk ), .D ( new_AGEMA_signal_1678 ), .Q ( new_AGEMA_signal_19394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C ( clk ), .D ( new_AGEMA_signal_1679 ), .Q ( new_AGEMA_signal_19396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C ( clk ), .D ( new_AGEMA_signal_1680 ), .Q ( new_AGEMA_signal_19398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C ( clk ), .D ( new_AGEMA_signal_1681 ), .Q ( new_AGEMA_signal_19400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C ( clk ), .D ( new_AGEMA_signal_18443 ), .Q ( new_AGEMA_signal_19402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C ( clk ), .D ( new_AGEMA_signal_18445 ), .Q ( new_AGEMA_signal_19406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C ( clk ), .D ( new_AGEMA_signal_18447 ), .Q ( new_AGEMA_signal_19410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C ( clk ), .D ( new_AGEMA_signal_18449 ), .Q ( new_AGEMA_signal_19414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C ( clk ), .D ( new_AGEMA_signal_18451 ), .Q ( new_AGEMA_signal_19418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_19422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C ( clk ), .D ( new_AGEMA_signal_1318 ), .Q ( new_AGEMA_signal_19426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C ( clk ), .D ( new_AGEMA_signal_1319 ), .Q ( new_AGEMA_signal_19430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C ( clk ), .D ( new_AGEMA_signal_1320 ), .Q ( new_AGEMA_signal_19434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C ( clk ), .D ( new_AGEMA_signal_1321 ), .Q ( new_AGEMA_signal_19438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_19462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C ( clk ), .D ( new_AGEMA_signal_1414 ), .Q ( new_AGEMA_signal_19466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C ( clk ), .D ( new_AGEMA_signal_1415 ), .Q ( new_AGEMA_signal_19470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C ( clk ), .D ( new_AGEMA_signal_1416 ), .Q ( new_AGEMA_signal_19474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C ( clk ), .D ( new_AGEMA_signal_1417 ), .Q ( new_AGEMA_signal_19478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C ( clk ), .D ( new_AGEMA_signal_18023 ), .Q ( new_AGEMA_signal_19492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C ( clk ), .D ( new_AGEMA_signal_18025 ), .Q ( new_AGEMA_signal_19496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C ( clk ), .D ( new_AGEMA_signal_18027 ), .Q ( new_AGEMA_signal_19500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C ( clk ), .D ( new_AGEMA_signal_18029 ), .Q ( new_AGEMA_signal_19504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C ( clk ), .D ( new_AGEMA_signal_18031 ), .Q ( new_AGEMA_signal_19508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_19522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C ( clk ), .D ( new_AGEMA_signal_1810 ), .Q ( new_AGEMA_signal_19526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C ( clk ), .D ( new_AGEMA_signal_1811 ), .Q ( new_AGEMA_signal_19530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C ( clk ), .D ( new_AGEMA_signal_1812 ), .Q ( new_AGEMA_signal_19534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C ( clk ), .D ( new_AGEMA_signal_1813 ), .Q ( new_AGEMA_signal_19538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_19542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C ( clk ), .D ( new_AGEMA_signal_1830 ), .Q ( new_AGEMA_signal_19546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C ( clk ), .D ( new_AGEMA_signal_1831 ), .Q ( new_AGEMA_signal_19550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C ( clk ), .D ( new_AGEMA_signal_1832 ), .Q ( new_AGEMA_signal_19554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C ( clk ), .D ( new_AGEMA_signal_1833 ), .Q ( new_AGEMA_signal_19558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_19602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C ( clk ), .D ( new_AGEMA_signal_1882 ), .Q ( new_AGEMA_signal_19606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C ( clk ), .D ( new_AGEMA_signal_1883 ), .Q ( new_AGEMA_signal_19610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C ( clk ), .D ( new_AGEMA_signal_1884 ), .Q ( new_AGEMA_signal_19614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C ( clk ), .D ( new_AGEMA_signal_1885 ), .Q ( new_AGEMA_signal_19618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_19622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C ( clk ), .D ( new_AGEMA_signal_1890 ), .Q ( new_AGEMA_signal_19626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C ( clk ), .D ( new_AGEMA_signal_1891 ), .Q ( new_AGEMA_signal_19630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C ( clk ), .D ( new_AGEMA_signal_1892 ), .Q ( new_AGEMA_signal_19634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C ( clk ), .D ( new_AGEMA_signal_1893 ), .Q ( new_AGEMA_signal_19638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_19642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C ( clk ), .D ( new_AGEMA_signal_1474 ), .Q ( new_AGEMA_signal_19646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C ( clk ), .D ( new_AGEMA_signal_1475 ), .Q ( new_AGEMA_signal_19650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C ( clk ), .D ( new_AGEMA_signal_1476 ), .Q ( new_AGEMA_signal_19654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C ( clk ), .D ( new_AGEMA_signal_1477 ), .Q ( new_AGEMA_signal_19658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_19692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C ( clk ), .D ( new_AGEMA_signal_1938 ), .Q ( new_AGEMA_signal_19696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C ( clk ), .D ( new_AGEMA_signal_1939 ), .Q ( new_AGEMA_signal_19700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C ( clk ), .D ( new_AGEMA_signal_1940 ), .Q ( new_AGEMA_signal_19704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C ( clk ), .D ( new_AGEMA_signal_1941 ), .Q ( new_AGEMA_signal_19708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C ( clk ), .D ( new_AGEMA_signal_17973 ), .Q ( new_AGEMA_signal_19722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C ( clk ), .D ( new_AGEMA_signal_17975 ), .Q ( new_AGEMA_signal_19726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C ( clk ), .D ( new_AGEMA_signal_17977 ), .Q ( new_AGEMA_signal_19730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C ( clk ), .D ( new_AGEMA_signal_17979 ), .Q ( new_AGEMA_signal_19734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C ( clk ), .D ( new_AGEMA_signal_17981 ), .Q ( new_AGEMA_signal_19738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C ( clk ), .D ( new_AGEMA_signal_19743 ), .Q ( new_AGEMA_signal_19744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C ( clk ), .D ( new_AGEMA_signal_19749 ), .Q ( new_AGEMA_signal_19750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C ( clk ), .D ( new_AGEMA_signal_19755 ), .Q ( new_AGEMA_signal_19756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C ( clk ), .D ( new_AGEMA_signal_19761 ), .Q ( new_AGEMA_signal_19762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C ( clk ), .D ( new_AGEMA_signal_19767 ), .Q ( new_AGEMA_signal_19768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C ( clk ), .D ( new_AGEMA_signal_18333 ), .Q ( new_AGEMA_signal_19772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C ( clk ), .D ( new_AGEMA_signal_18335 ), .Q ( new_AGEMA_signal_19776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C ( clk ), .D ( new_AGEMA_signal_18337 ), .Q ( new_AGEMA_signal_19780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C ( clk ), .D ( new_AGEMA_signal_18339 ), .Q ( new_AGEMA_signal_19784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C ( clk ), .D ( new_AGEMA_signal_18341 ), .Q ( new_AGEMA_signal_19788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C ( clk ), .D ( new_AGEMA_signal_18403 ), .Q ( new_AGEMA_signal_19792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C ( clk ), .D ( new_AGEMA_signal_18405 ), .Q ( new_AGEMA_signal_19796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C ( clk ), .D ( new_AGEMA_signal_18407 ), .Q ( new_AGEMA_signal_19800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C ( clk ), .D ( new_AGEMA_signal_18409 ), .Q ( new_AGEMA_signal_19804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C ( clk ), .D ( new_AGEMA_signal_18411 ), .Q ( new_AGEMA_signal_19808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_19852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C ( clk ), .D ( new_AGEMA_signal_2054 ), .Q ( new_AGEMA_signal_19856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C ( clk ), .D ( new_AGEMA_signal_2055 ), .Q ( new_AGEMA_signal_19860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C ( clk ), .D ( new_AGEMA_signal_2056 ), .Q ( new_AGEMA_signal_19864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C ( clk ), .D ( new_AGEMA_signal_2057 ), .Q ( new_AGEMA_signal_19868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C ( clk ), .D ( new_AGEMA_signal_19873 ), .Q ( new_AGEMA_signal_19874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C ( clk ), .D ( new_AGEMA_signal_19879 ), .Q ( new_AGEMA_signal_19880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C ( clk ), .D ( new_AGEMA_signal_19885 ), .Q ( new_AGEMA_signal_19886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C ( clk ), .D ( new_AGEMA_signal_19891 ), .Q ( new_AGEMA_signal_19892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C ( clk ), .D ( new_AGEMA_signal_19897 ), .Q ( new_AGEMA_signal_19898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_19902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C ( clk ), .D ( new_AGEMA_signal_1538 ), .Q ( new_AGEMA_signal_19906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C ( clk ), .D ( new_AGEMA_signal_1539 ), .Q ( new_AGEMA_signal_19910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C ( clk ), .D ( new_AGEMA_signal_1540 ), .Q ( new_AGEMA_signal_19914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C ( clk ), .D ( new_AGEMA_signal_1541 ), .Q ( new_AGEMA_signal_19918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_19952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C ( clk ), .D ( new_AGEMA_signal_2122 ), .Q ( new_AGEMA_signal_19956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C ( clk ), .D ( new_AGEMA_signal_2123 ), .Q ( new_AGEMA_signal_19960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C ( clk ), .D ( new_AGEMA_signal_2124 ), .Q ( new_AGEMA_signal_19964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C ( clk ), .D ( new_AGEMA_signal_2125 ), .Q ( new_AGEMA_signal_19968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C ( clk ), .D ( new_AGEMA_signal_18343 ), .Q ( new_AGEMA_signal_19992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C ( clk ), .D ( new_AGEMA_signal_18345 ), .Q ( new_AGEMA_signal_19996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C ( clk ), .D ( new_AGEMA_signal_18347 ), .Q ( new_AGEMA_signal_20000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C ( clk ), .D ( new_AGEMA_signal_18349 ), .Q ( new_AGEMA_signal_20004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C ( clk ), .D ( new_AGEMA_signal_18351 ), .Q ( new_AGEMA_signal_20008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C ( clk ), .D ( new_AGEMA_signal_18303 ), .Q ( new_AGEMA_signal_20012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C ( clk ), .D ( new_AGEMA_signal_18305 ), .Q ( new_AGEMA_signal_20016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C ( clk ), .D ( new_AGEMA_signal_18307 ), .Q ( new_AGEMA_signal_20020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C ( clk ), .D ( new_AGEMA_signal_18309 ), .Q ( new_AGEMA_signal_20024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C ( clk ), .D ( new_AGEMA_signal_18311 ), .Q ( new_AGEMA_signal_20028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C ( clk ), .D ( new_AGEMA_signal_17953 ), .Q ( new_AGEMA_signal_20032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C ( clk ), .D ( new_AGEMA_signal_17955 ), .Q ( new_AGEMA_signal_20036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C ( clk ), .D ( new_AGEMA_signal_17957 ), .Q ( new_AGEMA_signal_20040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C ( clk ), .D ( new_AGEMA_signal_17959 ), .Q ( new_AGEMA_signal_20044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C ( clk ), .D ( new_AGEMA_signal_17961 ), .Q ( new_AGEMA_signal_20048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C ( clk ), .D ( new_AGEMA_signal_18083 ), .Q ( new_AGEMA_signal_20052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C ( clk ), .D ( new_AGEMA_signal_18085 ), .Q ( new_AGEMA_signal_20056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C ( clk ), .D ( new_AGEMA_signal_18087 ), .Q ( new_AGEMA_signal_20060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C ( clk ), .D ( new_AGEMA_signal_18089 ), .Q ( new_AGEMA_signal_20064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C ( clk ), .D ( new_AGEMA_signal_18091 ), .Q ( new_AGEMA_signal_20068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_20072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C ( clk ), .D ( new_AGEMA_signal_2470 ), .Q ( new_AGEMA_signal_20076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C ( clk ), .D ( new_AGEMA_signal_2471 ), .Q ( new_AGEMA_signal_20080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C ( clk ), .D ( new_AGEMA_signal_2472 ), .Q ( new_AGEMA_signal_20084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C ( clk ), .D ( new_AGEMA_signal_2473 ), .Q ( new_AGEMA_signal_20088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C ( clk ), .D ( new_AGEMA_signal_18433 ), .Q ( new_AGEMA_signal_20132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C ( clk ), .D ( new_AGEMA_signal_18435 ), .Q ( new_AGEMA_signal_20136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C ( clk ), .D ( new_AGEMA_signal_18437 ), .Q ( new_AGEMA_signal_20140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C ( clk ), .D ( new_AGEMA_signal_18439 ), .Q ( new_AGEMA_signal_20144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C ( clk ), .D ( new_AGEMA_signal_18441 ), .Q ( new_AGEMA_signal_20148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_20152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C ( clk ), .D ( new_AGEMA_signal_1602 ), .Q ( new_AGEMA_signal_20156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C ( clk ), .D ( new_AGEMA_signal_1603 ), .Q ( new_AGEMA_signal_20160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C ( clk ), .D ( new_AGEMA_signal_1604 ), .Q ( new_AGEMA_signal_20164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C ( clk ), .D ( new_AGEMA_signal_1605 ), .Q ( new_AGEMA_signal_20168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_20262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C ( clk ), .D ( new_AGEMA_signal_1654 ), .Q ( new_AGEMA_signal_20266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_20270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C ( clk ), .D ( new_AGEMA_signal_1656 ), .Q ( new_AGEMA_signal_20274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C ( clk ), .D ( new_AGEMA_signal_1657 ), .Q ( new_AGEMA_signal_20278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_20332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C ( clk ), .D ( new_AGEMA_signal_1378 ), .Q ( new_AGEMA_signal_20336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C ( clk ), .D ( new_AGEMA_signal_1379 ), .Q ( new_AGEMA_signal_20340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C ( clk ), .D ( new_AGEMA_signal_1380 ), .Q ( new_AGEMA_signal_20344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C ( clk ), .D ( new_AGEMA_signal_1381 ), .Q ( new_AGEMA_signal_20348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C ( clk ), .D ( new_AGEMA_signal_18213 ), .Q ( new_AGEMA_signal_20352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C ( clk ), .D ( new_AGEMA_signal_18215 ), .Q ( new_AGEMA_signal_20356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C ( clk ), .D ( new_AGEMA_signal_18217 ), .Q ( new_AGEMA_signal_20360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C ( clk ), .D ( new_AGEMA_signal_18219 ), .Q ( new_AGEMA_signal_20364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C ( clk ), .D ( new_AGEMA_signal_18221 ), .Q ( new_AGEMA_signal_20368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C ( clk ), .D ( new_AGEMA_signal_18073 ), .Q ( new_AGEMA_signal_20372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C ( clk ), .D ( new_AGEMA_signal_18075 ), .Q ( new_AGEMA_signal_20376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C ( clk ), .D ( new_AGEMA_signal_18077 ), .Q ( new_AGEMA_signal_20380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C ( clk ), .D ( new_AGEMA_signal_18079 ), .Q ( new_AGEMA_signal_20384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C ( clk ), .D ( new_AGEMA_signal_18081 ), .Q ( new_AGEMA_signal_20388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_20392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C ( clk ), .D ( new_AGEMA_signal_2386 ), .Q ( new_AGEMA_signal_20396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C ( clk ), .D ( new_AGEMA_signal_2387 ), .Q ( new_AGEMA_signal_20400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C ( clk ), .D ( new_AGEMA_signal_2388 ), .Q ( new_AGEMA_signal_20404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C ( clk ), .D ( new_AGEMA_signal_2389 ), .Q ( new_AGEMA_signal_20408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C ( clk ), .D ( new_AGEMA_signal_20453 ), .Q ( new_AGEMA_signal_20454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C ( clk ), .D ( new_AGEMA_signal_20461 ), .Q ( new_AGEMA_signal_20462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C ( clk ), .D ( new_AGEMA_signal_20469 ), .Q ( new_AGEMA_signal_20470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C ( clk ), .D ( new_AGEMA_signal_20477 ), .Q ( new_AGEMA_signal_20478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C ( clk ), .D ( new_AGEMA_signal_20485 ), .Q ( new_AGEMA_signal_20486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C ( clk ), .D ( new_AGEMA_signal_20503 ), .Q ( new_AGEMA_signal_20504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C ( clk ), .D ( new_AGEMA_signal_20511 ), .Q ( new_AGEMA_signal_20512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C ( clk ), .D ( new_AGEMA_signal_20519 ), .Q ( new_AGEMA_signal_20520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C ( clk ), .D ( new_AGEMA_signal_20527 ), .Q ( new_AGEMA_signal_20528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C ( clk ), .D ( new_AGEMA_signal_20535 ), .Q ( new_AGEMA_signal_20536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_20542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_20548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C ( clk ), .D ( new_AGEMA_signal_1823 ), .Q ( new_AGEMA_signal_20554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C ( clk ), .D ( new_AGEMA_signal_1824 ), .Q ( new_AGEMA_signal_20560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C ( clk ), .D ( new_AGEMA_signal_1825 ), .Q ( new_AGEMA_signal_20566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_20592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C ( clk ), .D ( new_AGEMA_signal_1462 ), .Q ( new_AGEMA_signal_20598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C ( clk ), .D ( new_AGEMA_signal_1463 ), .Q ( new_AGEMA_signal_20604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C ( clk ), .D ( new_AGEMA_signal_1464 ), .Q ( new_AGEMA_signal_20610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C ( clk ), .D ( new_AGEMA_signal_1465 ), .Q ( new_AGEMA_signal_20616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C ( clk ), .D ( new_AGEMA_signal_18423 ), .Q ( new_AGEMA_signal_20632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C ( clk ), .D ( new_AGEMA_signal_18425 ), .Q ( new_AGEMA_signal_20638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C ( clk ), .D ( new_AGEMA_signal_18427 ), .Q ( new_AGEMA_signal_20644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C ( clk ), .D ( new_AGEMA_signal_18429 ), .Q ( new_AGEMA_signal_20650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C ( clk ), .D ( new_AGEMA_signal_18431 ), .Q ( new_AGEMA_signal_20656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C ( clk ), .D ( new_AGEMA_signal_18493 ), .Q ( new_AGEMA_signal_20662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C ( clk ), .D ( new_AGEMA_signal_18495 ), .Q ( new_AGEMA_signal_20668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C ( clk ), .D ( new_AGEMA_signal_18497 ), .Q ( new_AGEMA_signal_20674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C ( clk ), .D ( new_AGEMA_signal_18499 ), .Q ( new_AGEMA_signal_20680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C ( clk ), .D ( new_AGEMA_signal_18501 ), .Q ( new_AGEMA_signal_20686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C ( clk ), .D ( new_AGEMA_signal_17863 ), .Q ( new_AGEMA_signal_20722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C ( clk ), .D ( new_AGEMA_signal_17865 ), .Q ( new_AGEMA_signal_20728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C ( clk ), .D ( new_AGEMA_signal_17867 ), .Q ( new_AGEMA_signal_20734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C ( clk ), .D ( new_AGEMA_signal_17869 ), .Q ( new_AGEMA_signal_20740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C ( clk ), .D ( new_AGEMA_signal_17871 ), .Q ( new_AGEMA_signal_20746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_20752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C ( clk ), .D ( new_AGEMA_signal_1946 ), .Q ( new_AGEMA_signal_20758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C ( clk ), .D ( new_AGEMA_signal_1947 ), .Q ( new_AGEMA_signal_20764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C ( clk ), .D ( new_AGEMA_signal_1948 ), .Q ( new_AGEMA_signal_20770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C ( clk ), .D ( new_AGEMA_signal_1949 ), .Q ( new_AGEMA_signal_20776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_20792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C ( clk ), .D ( new_AGEMA_signal_1970 ), .Q ( new_AGEMA_signal_20798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C ( clk ), .D ( new_AGEMA_signal_1971 ), .Q ( new_AGEMA_signal_20804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C ( clk ), .D ( new_AGEMA_signal_1972 ), .Q ( new_AGEMA_signal_20810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C ( clk ), .D ( new_AGEMA_signal_1973 ), .Q ( new_AGEMA_signal_20816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C ( clk ), .D ( new_AGEMA_signal_20883 ), .Q ( new_AGEMA_signal_20884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C ( clk ), .D ( new_AGEMA_signal_20891 ), .Q ( new_AGEMA_signal_20892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C ( clk ), .D ( new_AGEMA_signal_20899 ), .Q ( new_AGEMA_signal_20900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C ( clk ), .D ( new_AGEMA_signal_20907 ), .Q ( new_AGEMA_signal_20908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C ( clk ), .D ( new_AGEMA_signal_20915 ), .Q ( new_AGEMA_signal_20916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C ( clk ), .D ( new_AGEMA_signal_18113 ), .Q ( new_AGEMA_signal_20922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C ( clk ), .D ( new_AGEMA_signal_18115 ), .Q ( new_AGEMA_signal_20928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C ( clk ), .D ( new_AGEMA_signal_18117 ), .Q ( new_AGEMA_signal_20934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C ( clk ), .D ( new_AGEMA_signal_18119 ), .Q ( new_AGEMA_signal_20940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C ( clk ), .D ( new_AGEMA_signal_18121 ), .Q ( new_AGEMA_signal_20946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_21062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C ( clk ), .D ( new_AGEMA_signal_2130 ), .Q ( new_AGEMA_signal_21068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C ( clk ), .D ( new_AGEMA_signal_2131 ), .Q ( new_AGEMA_signal_21074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C ( clk ), .D ( new_AGEMA_signal_2132 ), .Q ( new_AGEMA_signal_21080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C ( clk ), .D ( new_AGEMA_signal_2133 ), .Q ( new_AGEMA_signal_21086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_21222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C ( clk ), .D ( new_AGEMA_signal_1614 ), .Q ( new_AGEMA_signal_21228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C ( clk ), .D ( new_AGEMA_signal_1615 ), .Q ( new_AGEMA_signal_21234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C ( clk ), .D ( new_AGEMA_signal_1616 ), .Q ( new_AGEMA_signal_21240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C ( clk ), .D ( new_AGEMA_signal_1617 ), .Q ( new_AGEMA_signal_21246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_21252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C ( clk ), .D ( new_AGEMA_signal_1750 ), .Q ( new_AGEMA_signal_21258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C ( clk ), .D ( new_AGEMA_signal_1751 ), .Q ( new_AGEMA_signal_21264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C ( clk ), .D ( new_AGEMA_signal_1752 ), .Q ( new_AGEMA_signal_21270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C ( clk ), .D ( new_AGEMA_signal_1753 ), .Q ( new_AGEMA_signal_21276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C ( clk ), .D ( new_AGEMA_signal_21313 ), .Q ( new_AGEMA_signal_21314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C ( clk ), .D ( new_AGEMA_signal_21321 ), .Q ( new_AGEMA_signal_21322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C ( clk ), .D ( new_AGEMA_signal_21329 ), .Q ( new_AGEMA_signal_21330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C ( clk ), .D ( new_AGEMA_signal_21337 ), .Q ( new_AGEMA_signal_21338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C ( clk ), .D ( new_AGEMA_signal_21345 ), .Q ( new_AGEMA_signal_21346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C ( clk ), .D ( new_AGEMA_signal_21463 ), .Q ( new_AGEMA_signal_21464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C ( clk ), .D ( new_AGEMA_signal_21471 ), .Q ( new_AGEMA_signal_21472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C ( clk ), .D ( new_AGEMA_signal_21479 ), .Q ( new_AGEMA_signal_21480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C ( clk ), .D ( new_AGEMA_signal_21487 ), .Q ( new_AGEMA_signal_21488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C ( clk ), .D ( new_AGEMA_signal_21495 ), .Q ( new_AGEMA_signal_21496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_21542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C ( clk ), .D ( new_AGEMA_signal_2406 ), .Q ( new_AGEMA_signal_21548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C ( clk ), .D ( new_AGEMA_signal_2407 ), .Q ( new_AGEMA_signal_21554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C ( clk ), .D ( new_AGEMA_signal_2408 ), .Q ( new_AGEMA_signal_21560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C ( clk ), .D ( new_AGEMA_signal_2409 ), .Q ( new_AGEMA_signal_21566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_21582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C ( clk ), .D ( new_AGEMA_signal_1370 ), .Q ( new_AGEMA_signal_21590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C ( clk ), .D ( new_AGEMA_signal_1371 ), .Q ( new_AGEMA_signal_21598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_21606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C ( clk ), .D ( new_AGEMA_signal_1373 ), .Q ( new_AGEMA_signal_21614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_21652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C ( clk ), .D ( new_AGEMA_signal_1450 ), .Q ( new_AGEMA_signal_21660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C ( clk ), .D ( new_AGEMA_signal_1451 ), .Q ( new_AGEMA_signal_21668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C ( clk ), .D ( new_AGEMA_signal_1452 ), .Q ( new_AGEMA_signal_21676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C ( clk ), .D ( new_AGEMA_signal_1453 ), .Q ( new_AGEMA_signal_21684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_21752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C ( clk ), .D ( new_AGEMA_signal_1950 ), .Q ( new_AGEMA_signal_21760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C ( clk ), .D ( new_AGEMA_signal_1951 ), .Q ( new_AGEMA_signal_21768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C ( clk ), .D ( new_AGEMA_signal_1952 ), .Q ( new_AGEMA_signal_21776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C ( clk ), .D ( new_AGEMA_signal_1953 ), .Q ( new_AGEMA_signal_21784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C ( clk ), .D ( new_AGEMA_signal_18523 ), .Q ( new_AGEMA_signal_21982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C ( clk ), .D ( new_AGEMA_signal_18525 ), .Q ( new_AGEMA_signal_21990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C ( clk ), .D ( new_AGEMA_signal_18527 ), .Q ( new_AGEMA_signal_21998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C ( clk ), .D ( new_AGEMA_signal_18529 ), .Q ( new_AGEMA_signal_22006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C ( clk ), .D ( new_AGEMA_signal_18531 ), .Q ( new_AGEMA_signal_22014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_22072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C ( clk ), .D ( new_AGEMA_signal_1582 ), .Q ( new_AGEMA_signal_22080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C ( clk ), .D ( new_AGEMA_signal_1583 ), .Q ( new_AGEMA_signal_22088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C ( clk ), .D ( new_AGEMA_signal_1584 ), .Q ( new_AGEMA_signal_22096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C ( clk ), .D ( new_AGEMA_signal_1585 ), .Q ( new_AGEMA_signal_22104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C ( clk ), .D ( new_AGEMA_signal_18413 ), .Q ( new_AGEMA_signal_22232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C ( clk ), .D ( new_AGEMA_signal_18415 ), .Q ( new_AGEMA_signal_22240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C ( clk ), .D ( new_AGEMA_signal_18417 ), .Q ( new_AGEMA_signal_22248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C ( clk ), .D ( new_AGEMA_signal_18419 ), .Q ( new_AGEMA_signal_22256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C ( clk ), .D ( new_AGEMA_signal_18421 ), .Q ( new_AGEMA_signal_22264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C ( clk ), .D ( new_AGEMA_signal_17913 ), .Q ( new_AGEMA_signal_22272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C ( clk ), .D ( new_AGEMA_signal_17915 ), .Q ( new_AGEMA_signal_22280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C ( clk ), .D ( new_AGEMA_signal_17917 ), .Q ( new_AGEMA_signal_22288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C ( clk ), .D ( new_AGEMA_signal_17919 ), .Q ( new_AGEMA_signal_22296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C ( clk ), .D ( new_AGEMA_signal_17921 ), .Q ( new_AGEMA_signal_22304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_22702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C ( clk ), .D ( new_AGEMA_signal_1490 ), .Q ( new_AGEMA_signal_22712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C ( clk ), .D ( new_AGEMA_signal_1491 ), .Q ( new_AGEMA_signal_22722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C ( clk ), .D ( new_AGEMA_signal_1492 ), .Q ( new_AGEMA_signal_22732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C ( clk ), .D ( new_AGEMA_signal_1493 ), .Q ( new_AGEMA_signal_22742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_22952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C ( clk ), .D ( new_AGEMA_signal_2154 ), .Q ( new_AGEMA_signal_22962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C ( clk ), .D ( new_AGEMA_signal_2155 ), .Q ( new_AGEMA_signal_22972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C ( clk ), .D ( new_AGEMA_signal_2156 ), .Q ( new_AGEMA_signal_22982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C ( clk ), .D ( new_AGEMA_signal_2157 ), .Q ( new_AGEMA_signal_22992 ) ) ;

    /* cells in depth 6 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1960 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, n2575}), .inb ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n1962}), .clk ( clk ), .rnd ({Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .outt ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, n1924}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1967 ( .ina ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, n1922}), .inb ({new_AGEMA_signal_17861, new_AGEMA_signal_17859, new_AGEMA_signal_17857, new_AGEMA_signal_17855, new_AGEMA_signal_17853}), .clk ( clk ), .rnd ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585]}), .outt ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, n1923}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1981 ( .ina ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1694, n1926}), .inb ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n1925}), .clk ( clk ), .rnd ({Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .outt ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n1927}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1993 ( .ina ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2734}), .inb ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2763}), .clk ( clk ), .rnd ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615]}), .outt ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, n1929}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2007 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .clk ( clk ), .rnd ({Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .outt ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, n2665}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2011 ( .ina ({new_AGEMA_signal_17881, new_AGEMA_signal_17879, new_AGEMA_signal_17877, new_AGEMA_signal_17875, new_AGEMA_signal_17873}), .inb ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1718, n1937}), .clk ( clk ), .rnd ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645]}), .outt ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n1938}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2019 ( .ina ({new_AGEMA_signal_17891, new_AGEMA_signal_17889, new_AGEMA_signal_17887, new_AGEMA_signal_17885, new_AGEMA_signal_17883}), .inb ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .clk ( clk ), .rnd ({Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .outt ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, n2235}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2023 ( .ina ({new_AGEMA_signal_17901, new_AGEMA_signal_17899, new_AGEMA_signal_17897, new_AGEMA_signal_17895, new_AGEMA_signal_17893}), .inb ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, new_AGEMA_signal_1343, new_AGEMA_signal_1342, n1942}), .clk ( clk ), .rnd ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675]}), .outt ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n1943}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2027 ( .ina ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2676}), .inb ({new_AGEMA_signal_17911, new_AGEMA_signal_17909, new_AGEMA_signal_17907, new_AGEMA_signal_17905, new_AGEMA_signal_17903}), .clk ( clk ), .rnd ({Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .outt ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, n1946}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2031 ( .ina ({new_AGEMA_signal_17921, new_AGEMA_signal_17919, new_AGEMA_signal_17917, new_AGEMA_signal_17915, new_AGEMA_signal_17913}), .inb ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1730, n1944}), .clk ( clk ), .rnd ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705]}), .outt ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, n1945}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2034 ( .ina ({new_AGEMA_signal_17931, new_AGEMA_signal_17929, new_AGEMA_signal_17927, new_AGEMA_signal_17925, new_AGEMA_signal_17923}), .inb ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2734}), .clk ( clk ), .rnd ({Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .outt ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n1956}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2040 ( .ina ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n1950}), .inb ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, n1949}), .clk ( clk ), .rnd ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735]}), .outt ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, n1951}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2048 ( .ina ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2662}), .inb ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}), .clk ( clk ), .rnd ({Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .outt ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, n1952}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2057 ( .ina ({new_AGEMA_signal_17941, new_AGEMA_signal_17939, new_AGEMA_signal_17937, new_AGEMA_signal_17935, new_AGEMA_signal_17933}), .inb ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, n2088}), .clk ( clk ), .rnd ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765]}), .outt ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2687}) ) ;
    or_HPC1 #(.security_order(4), .pipeline(1)) U2061 ( .ina ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n1962}), .inb ({new_AGEMA_signal_17951, new_AGEMA_signal_17949, new_AGEMA_signal_17947, new_AGEMA_signal_17945, new_AGEMA_signal_17943}), .clk ( clk ), .rnd ({Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .outt ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, n1966}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2064 ( .ina ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2736}), .inb ({new_AGEMA_signal_17961, new_AGEMA_signal_17959, new_AGEMA_signal_17957, new_AGEMA_signal_17955, new_AGEMA_signal_17953}), .clk ( clk ), .rnd ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795]}), .outt ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n1963}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2077 ( .ina ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2720}), .inb ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .clk ( clk ), .rnd ({Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .outt ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, n1968}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2082 ( .ina ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2505}), .inb ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825]}), .outt ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, n2684}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2088 ( .ina ({new_AGEMA_signal_17971, new_AGEMA_signal_17969, new_AGEMA_signal_17967, new_AGEMA_signal_17965, new_AGEMA_signal_17963}), .inb ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2625}), .clk ( clk ), .rnd ({Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .outt ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n1972}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2092 ( .ina ({new_AGEMA_signal_17981, new_AGEMA_signal_17979, new_AGEMA_signal_17977, new_AGEMA_signal_17975, new_AGEMA_signal_17973}), .inb ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2190}), .clk ( clk ), .rnd ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855]}), .outt ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n1971}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2099 ( .ina ({new_AGEMA_signal_17991, new_AGEMA_signal_17989, new_AGEMA_signal_17987, new_AGEMA_signal_17985, new_AGEMA_signal_17983}), .inb ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, n2535}), .clk ( clk ), .rnd ({Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .outt ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, n1974}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2106 ( .ina ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .inb ({new_AGEMA_signal_17941, new_AGEMA_signal_17939, new_AGEMA_signal_17937, new_AGEMA_signal_17935, new_AGEMA_signal_17933}), .clk ( clk ), .rnd ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885]}), .outt ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, n1979}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2112 ( .ina ({new_AGEMA_signal_18001, new_AGEMA_signal_17999, new_AGEMA_signal_17997, new_AGEMA_signal_17995, new_AGEMA_signal_17993}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .outt ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n1985}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2121 ( .ina ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, n1992}), .inb ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n1991}), .clk ( clk ), .rnd ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915]}), .outt ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, n1994}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2126 ( .ina ({new_AGEMA_signal_18011, new_AGEMA_signal_18009, new_AGEMA_signal_18007, new_AGEMA_signal_18005, new_AGEMA_signal_18003}), .inb ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, n1995}), .clk ( clk ), .rnd ({Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .outt ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, n1996}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2136 ( .ina ({new_AGEMA_signal_18021, new_AGEMA_signal_18019, new_AGEMA_signal_18017, new_AGEMA_signal_18015, new_AGEMA_signal_18013}), .inb ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2003}), .clk ( clk ), .rnd ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945]}), .outt ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2137}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2142 ( .ina ({new_AGEMA_signal_18031, new_AGEMA_signal_18029, new_AGEMA_signal_18027, new_AGEMA_signal_18025, new_AGEMA_signal_18023}), .inb ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2572}), .clk ( clk ), .rnd ({Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .outt ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, n2006}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2144 ( .ina ({new_AGEMA_signal_18041, new_AGEMA_signal_18039, new_AGEMA_signal_18037, new_AGEMA_signal_18035, new_AGEMA_signal_18033}), .inb ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2004}), .clk ( clk ), .rnd ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975]}), .outt ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, n2005}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2152 ( .ina ({new_AGEMA_signal_18051, new_AGEMA_signal_18049, new_AGEMA_signal_18047, new_AGEMA_signal_18045, new_AGEMA_signal_18043}), .inb ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .clk ( clk ), .rnd ({Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .outt ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2013}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2160 ( .ina ({new_AGEMA_signal_18061, new_AGEMA_signal_18059, new_AGEMA_signal_18057, new_AGEMA_signal_18055, new_AGEMA_signal_18053}), .inb ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, n2227}), .clk ( clk ), .rnd ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005]}), .outt ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, new_AGEMA_signal_1834, n2020}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2164 ( .ina ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .inb ({new_AGEMA_signal_18071, new_AGEMA_signal_18069, new_AGEMA_signal_18067, new_AGEMA_signal_18065, new_AGEMA_signal_18063}), .clk ( clk ), .rnd ({Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .outt ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, n2023}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2168 ( .ina ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, n2027}), .inb ({new_AGEMA_signal_18081, new_AGEMA_signal_18079, new_AGEMA_signal_18077, new_AGEMA_signal_18075, new_AGEMA_signal_18073}), .clk ( clk ), .rnd ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035]}), .outt ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2028}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2172 ( .ina ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2214}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .outt ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, new_AGEMA_signal_2522, n2033}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2175 ( .ina ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}), .inb ({new_AGEMA_signal_18101, new_AGEMA_signal_18099, new_AGEMA_signal_18097, new_AGEMA_signal_18095, new_AGEMA_signal_18093}), .clk ( clk ), .rnd ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065]}), .outt ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n2031}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2184 ( .ina ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}), .inb ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2039}), .clk ( clk ), .rnd ({Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .outt ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, n2040}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2187 ( .ina ({new_AGEMA_signal_18111, new_AGEMA_signal_18109, new_AGEMA_signal_18107, new_AGEMA_signal_18105, new_AGEMA_signal_18103}), .inb ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095]}), .outt ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, n2050}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2193 ( .ina ({new_AGEMA_signal_18121, new_AGEMA_signal_18119, new_AGEMA_signal_18117, new_AGEMA_signal_18115, new_AGEMA_signal_18113}), .inb ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, n2044}), .clk ( clk ), .rnd ({Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .outt ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, n2045}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2199 ( .ina ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2654}), .inb ({new_AGEMA_signal_17941, new_AGEMA_signal_17939, new_AGEMA_signal_17937, new_AGEMA_signal_17935, new_AGEMA_signal_17933}), .clk ( clk ), .rnd ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125]}), .outt ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n2051}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2203 ( .ina ({new_AGEMA_signal_18131, new_AGEMA_signal_18129, new_AGEMA_signal_18127, new_AGEMA_signal_18125, new_AGEMA_signal_18123}), .inb ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2055}), .clk ( clk ), .rnd ({Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .outt ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, n2056}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2209 ( .ina ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, n2407}), .inb ({new_AGEMA_signal_18141, new_AGEMA_signal_18139, new_AGEMA_signal_18137, new_AGEMA_signal_18135, new_AGEMA_signal_18133}), .clk ( clk ), .rnd ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155]}), .outt ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, n2060}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2215 ( .ina ({new_AGEMA_signal_18151, new_AGEMA_signal_18149, new_AGEMA_signal_18147, new_AGEMA_signal_18145, new_AGEMA_signal_18143}), .inb ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2654}), .clk ( clk ), .rnd ({Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .outt ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2066}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2217 ( .ina ({new_AGEMA_signal_18081, new_AGEMA_signal_18079, new_AGEMA_signal_18077, new_AGEMA_signal_18075, new_AGEMA_signal_18073}), .inb ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2731}), .clk ( clk ), .rnd ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185]}), .outt ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, n2065}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2221 ( .ina ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, n2068}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .outt ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, n2069}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2226 ( .ina ({new_AGEMA_signal_18161, new_AGEMA_signal_18159, new_AGEMA_signal_18157, new_AGEMA_signal_18155, new_AGEMA_signal_18153}), .inb ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2252}), .clk ( clk ), .rnd ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215]}), .outt ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n2074}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2235 ( .ina ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1478, n2081}), .inb ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, n2080}), .clk ( clk ), .rnd ({Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .outt ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, n2082}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2240 ( .ina ({new_AGEMA_signal_18041, new_AGEMA_signal_18039, new_AGEMA_signal_18037, new_AGEMA_signal_18035, new_AGEMA_signal_18033}), .inb ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2083}), .clk ( clk ), .rnd ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245]}), .outt ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, n2084}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2242 ( .ina ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .inb ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .clk ( clk ), .rnd ({Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .outt ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n2085}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2245 ( .ina ({new_AGEMA_signal_18171, new_AGEMA_signal_18169, new_AGEMA_signal_18167, new_AGEMA_signal_18165, new_AGEMA_signal_18163}), .inb ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, n2562}), .clk ( clk ), .rnd ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275]}), .outt ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, n2131}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2248 ( .ina ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, n2088}), .inb ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, n2087}), .clk ( clk ), .rnd ({Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .outt ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, new_AGEMA_signal_2582, n2089}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2252 ( .ina ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .inb ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, n2156}), .clk ( clk ), .rnd ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305]}), .outt ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2330}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2254 ( .ina ({new_AGEMA_signal_18181, new_AGEMA_signal_18179, new_AGEMA_signal_18177, new_AGEMA_signal_18175, new_AGEMA_signal_18173}), .inb ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, n2151}), .clk ( clk ), .rnd ({Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .outt ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, n2092}) ) ;
    or_HPC1 #(.security_order(4), .pipeline(1)) U2256 ( .ina ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}), .inb ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, n2359}), .clk ( clk ), .rnd ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335]}), .outt ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, n2094}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2261 ( .ina ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, new_AGEMA_signal_1402, n2101}), .inb ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2100}), .clk ( clk ), .rnd ({Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .outt ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2160}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2265 ( .ina ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365]}), .outt ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, n2504}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2271 ( .ina ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .inb ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .outt ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, n2114}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2273 ( .ina ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2677}), .inb ({new_AGEMA_signal_18041, new_AGEMA_signal_18039, new_AGEMA_signal_18037, new_AGEMA_signal_18035, new_AGEMA_signal_18033}), .clk ( clk ), .rnd ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395]}), .outt ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1934, n2115}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2280 ( .ina ({new_AGEMA_signal_18191, new_AGEMA_signal_18189, new_AGEMA_signal_18187, new_AGEMA_signal_18185, new_AGEMA_signal_18183}), .inb ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2731}), .clk ( clk ), .rnd ({Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .outt ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, n2291}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2281 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .clk ( clk ), .rnd ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425]}), .outt ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, new_AGEMA_signal_1942, n2119}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2291 ( .ina ({new_AGEMA_signal_18201, new_AGEMA_signal_18199, new_AGEMA_signal_18197, new_AGEMA_signal_18195, new_AGEMA_signal_18193}), .inb ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .clk ( clk ), .rnd ({Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .outt ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, n2130}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2292 ( .ina ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .inb ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2631}), .clk ( clk ), .rnd ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455]}), .outt ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, n2129}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2295 ( .ina ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, n2647}), .inb ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .clk ( clk ), .rnd ({Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .outt ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2150}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2298 ( .ina ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}), .inb ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, n2132}), .clk ( clk ), .rnd ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485]}), .outt ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, n2133}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2302 ( .ina ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .inb ({new_AGEMA_signal_18221, new_AGEMA_signal_18219, new_AGEMA_signal_18217, new_AGEMA_signal_18215, new_AGEMA_signal_18213}), .clk ( clk ), .rnd ({Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .outt ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, n2136}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2306 ( .ina ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2572}), .inb ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2138}), .clk ( clk ), .rnd ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515]}), .outt ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2139}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2313 ( .ina ({new_AGEMA_signal_18231, new_AGEMA_signal_18229, new_AGEMA_signal_18227, new_AGEMA_signal_18225, new_AGEMA_signal_18223}), .inb ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, n2555}), .clk ( clk ), .rnd ({Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .outt ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, n2144}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2318 ( .ina ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, n2151}), .inb ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .clk ( clk ), .rnd ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545]}), .outt ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, n2152}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2321 ( .ina ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}), .inb ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, n2156}), .clk ( clk ), .rnd ({Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .outt ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2170}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2323 ( .ina ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2429}), .inb ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .clk ( clk ), .rnd ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575]}), .outt ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, n2157}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2329 ( .ina ({new_AGEMA_signal_18241, new_AGEMA_signal_18239, new_AGEMA_signal_18237, new_AGEMA_signal_18235, new_AGEMA_signal_18233}), .inb ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n2162}), .clk ( clk ), .rnd ({Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .outt ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2163}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2335 ( .ina ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, n2171}), .inb ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}), .clk ( clk ), .rnd ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605]}), .outt ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2172}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2338 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2545}), .clk ( clk ), .rnd ({Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .outt ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, n2186}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2339 ( .ina ({new_AGEMA_signal_17991, new_AGEMA_signal_17989, new_AGEMA_signal_17987, new_AGEMA_signal_17985, new_AGEMA_signal_17983}), .inb ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, n2290}), .clk ( clk ), .rnd ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635]}), .outt ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, n2181}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2344 ( .ina ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, n2176}), .inb ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, n2175}), .clk ( clk ), .rnd ({Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .outt ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, n2177}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2349 ( .ina ({new_AGEMA_signal_17941, new_AGEMA_signal_17939, new_AGEMA_signal_17937, new_AGEMA_signal_17935, new_AGEMA_signal_17933}), .inb ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, n2182}), .clk ( clk ), .rnd ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665]}), .outt ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2183}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2354 ( .ina ({new_AGEMA_signal_18251, new_AGEMA_signal_18249, new_AGEMA_signal_18247, new_AGEMA_signal_18245, new_AGEMA_signal_18243}), .inb ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2188}), .clk ( clk ), .rnd ({Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .outt ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2195}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2356 ( .ina ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2190}), .inb ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, n2189}), .clk ( clk ), .rnd ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695]}), .outt ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, n2193}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2358 ( .ina ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .inb ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, n2446}), .clk ( clk ), .rnd ({Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .outt ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, n2191}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2364 ( .ina ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2576}), .inb ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, n2748}), .clk ( clk ), .rnd ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725]}), .outt ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2196}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2367 ( .ina ({new_AGEMA_signal_17911, new_AGEMA_signal_17909, new_AGEMA_signal_17907, new_AGEMA_signal_17905, new_AGEMA_signal_17903}), .inb ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2505}), .clk ( clk ), .rnd ({Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .outt ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2201}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2369 ( .ina ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2674}), .inb ({new_AGEMA_signal_18271, new_AGEMA_signal_18269, new_AGEMA_signal_18267, new_AGEMA_signal_18265, new_AGEMA_signal_18263}), .clk ( clk ), .rnd ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755]}), .outt ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2200}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2371 ( .ins ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2734}), .ina ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .clk ( clk ), .rnd ({Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .outt ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, n2202}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2379 ( .ina ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2214}), .inb ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n2213}), .clk ( clk ), .rnd ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785]}), .outt ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, n2217}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2381 ( .ina ({new_AGEMA_signal_18281, new_AGEMA_signal_18279, new_AGEMA_signal_18277, new_AGEMA_signal_18275, new_AGEMA_signal_18273}), .inb ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, n2215}), .clk ( clk ), .rnd ({Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .outt ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, new_AGEMA_signal_2014, n2216}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2385 ( .ina ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, n2218}), .inb ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .clk ( clk ), .rnd ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815]}), .outt ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2222}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2387 ( .ina ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1970, n2220}), .inb ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2219}), .clk ( clk ), .rnd ({Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .outt ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, n2221}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2391 ( .ina ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}), .inb ({new_AGEMA_signal_18291, new_AGEMA_signal_18289, new_AGEMA_signal_18287, new_AGEMA_signal_18285, new_AGEMA_signal_18283}), .clk ( clk ), .rnd ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845]}), .outt ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, n2226}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2393 ( .ins ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .ina ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, n2227}), .clk ( clk ), .rnd ({Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .outt ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, new_AGEMA_signal_2030, n2228}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2397 ( .ina ({new_AGEMA_signal_18061, new_AGEMA_signal_18059, new_AGEMA_signal_18057, new_AGEMA_signal_18055, new_AGEMA_signal_18053}), .inb ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875]}), .outt ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2237}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2398 ( .ina ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .inb ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .clk ( clk ), .rnd ({Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .outt ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, new_AGEMA_signal_3254, n2233}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2403 ( .ina ({new_AGEMA_signal_18301, new_AGEMA_signal_18299, new_AGEMA_signal_18297, new_AGEMA_signal_18295, new_AGEMA_signal_18293}), .inb ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2631}), .clk ( clk ), .rnd ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905]}), .outt ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, n2238}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2406 ( .ina ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, n2241}), .inb ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, n2240}), .clk ( clk ), .rnd ({Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .outt ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2248}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2409 ( .ina ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n2561}), .inb ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, n2243}), .clk ( clk ), .rnd ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935]}), .outt ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, n2244}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2414 ( .ina ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}), .inb ({new_AGEMA_signal_17861, new_AGEMA_signal_17859, new_AGEMA_signal_17857, new_AGEMA_signal_17855, new_AGEMA_signal_17853}), .clk ( clk ), .rnd ({Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .outt ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, n2249}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2417 ( .ins ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2252}), .ina ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965]}), .outt ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2253}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2424 ( .ina ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .inb ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, n2259}), .clk ( clk ), .rnd ({Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .outt ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, n2260}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2429 ( .ina ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .inb ({new_AGEMA_signal_18311, new_AGEMA_signal_18309, new_AGEMA_signal_18307, new_AGEMA_signal_18305, new_AGEMA_signal_18303}), .clk ( clk ), .rnd ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995]}), .outt ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2273}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2430 ( .ina ({new_AGEMA_signal_18321, new_AGEMA_signal_18319, new_AGEMA_signal_18317, new_AGEMA_signal_18315, new_AGEMA_signal_18313}), .inb ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2720}), .clk ( clk ), .rnd ({Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .outt ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, n2752}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2433 ( .ina ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, n2645}), .inb ({new_AGEMA_signal_18191, new_AGEMA_signal_18189, new_AGEMA_signal_18187, new_AGEMA_signal_18185, new_AGEMA_signal_18183}), .clk ( clk ), .rnd ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025]}), .outt ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, n2265}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2437 ( .ina ({new_AGEMA_signal_18331, new_AGEMA_signal_18329, new_AGEMA_signal_18327, new_AGEMA_signal_18325, new_AGEMA_signal_18323}), .inb ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, n2268}), .clk ( clk ), .rnd ({Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .outt ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n2269}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2444 ( .ina ({new_AGEMA_signal_17961, new_AGEMA_signal_17959, new_AGEMA_signal_17957, new_AGEMA_signal_17955, new_AGEMA_signal_17953}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055]}), .outt ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, n2277}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2449 ( .ina ({new_AGEMA_signal_18341, new_AGEMA_signal_18339, new_AGEMA_signal_18337, new_AGEMA_signal_18335, new_AGEMA_signal_18333}), .inb ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2383}), .clk ( clk ), .rnd ({Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .outt ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n2282}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2452 ( .ina ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2736}), .inb ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .clk ( clk ), .rnd ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085]}), .outt ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2284}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2456 ( .ina ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2774}), .inb ({new_AGEMA_signal_18351, new_AGEMA_signal_18349, new_AGEMA_signal_18347, new_AGEMA_signal_18345, new_AGEMA_signal_18343}), .clk ( clk ), .rnd ({Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .outt ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, n2459}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2459 ( .ina ({new_AGEMA_signal_17881, new_AGEMA_signal_17879, new_AGEMA_signal_17877, new_AGEMA_signal_17875, new_AGEMA_signal_17873}), .inb ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, n2287}), .clk ( clk ), .rnd ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115]}), .outt ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, n2288}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2462 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}), .clk ( clk ), .rnd ({Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .outt ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2458}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2464 ( .ina ({new_AGEMA_signal_18241, new_AGEMA_signal_18239, new_AGEMA_signal_18237, new_AGEMA_signal_18235, new_AGEMA_signal_18233}), .inb ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, n2290}), .clk ( clk ), .rnd ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145]}), .outt ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, n2293}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2467 ( .ina ({new_AGEMA_signal_18181, new_AGEMA_signal_18179, new_AGEMA_signal_18177, new_AGEMA_signal_18175, new_AGEMA_signal_18173}), .inb ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2642}), .clk ( clk ), .rnd ({Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .outt ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n2294}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2472 ( .ina ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2438}), .inb ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, n2299}), .clk ( clk ), .rnd ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175]}), .outt ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, n2300}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2480 ( .ina ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2734}), .inb ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .clk ( clk ), .rnd ({Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .outt ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2323}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(1)) U2482 ( .ina ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2571}), .inb ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, n2371}), .clk ( clk ), .rnd ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205]}), .outt ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, n2314}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2485 ( .ina ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, n2316}), .inb ({new_AGEMA_signal_18361, new_AGEMA_signal_18359, new_AGEMA_signal_18357, new_AGEMA_signal_18355, new_AGEMA_signal_18353}), .clk ( clk ), .rnd ({Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .outt ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, n2319}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2491 ( .ina ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2642}), .inb ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .clk ( clk ), .rnd ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235]}), .outt ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, n2326}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2496 ( .ina ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2328}), .inb ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, n2327}), .clk ( clk ), .rnd ({Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .outt ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2329}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2501 ( .ina ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2417}), .inb ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2674}), .clk ( clk ), .rnd ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265]}), .outt ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, n2335}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2506 ( .ina ({new_AGEMA_signal_18051, new_AGEMA_signal_18049, new_AGEMA_signal_18047, new_AGEMA_signal_18045, new_AGEMA_signal_18043}), .inb ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}), .clk ( clk ), .rnd ({Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290], Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .outt ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, n2341}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2507 ( .ina ({new_AGEMA_signal_18371, new_AGEMA_signal_18369, new_AGEMA_signal_18367, new_AGEMA_signal_18365, new_AGEMA_signal_18363}), .inb ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2736}), .clk ( clk ), .rnd ({Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300], Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295]}), .outt ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, n2340}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2514 ( .ina ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, n2348}), .inb ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n2347}), .clk ( clk ), .rnd ({Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320], Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310]}), .outt ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, n2349}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2517 ( .ina ({new_AGEMA_signal_18381, new_AGEMA_signal_18379, new_AGEMA_signal_18377, new_AGEMA_signal_18375, new_AGEMA_signal_18373}), .inb ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2690}), .clk ( clk ), .rnd ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330], Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325]}), .outt ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, n2375}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2518 ( .ina ({new_AGEMA_signal_18231, new_AGEMA_signal_18229, new_AGEMA_signal_18227, new_AGEMA_signal_18225, new_AGEMA_signal_18223}), .inb ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2736}), .clk ( clk ), .rnd ({Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350], Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .outt ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2352}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2522 ( .ina ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, n2353}), .inb ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .clk ( clk ), .rnd ({Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360], Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355]}), .outt ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2354}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2525 ( .ina ({new_AGEMA_signal_18391, new_AGEMA_signal_18389, new_AGEMA_signal_18387, new_AGEMA_signal_18385, new_AGEMA_signal_18383}), .inb ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, n2355}), .clk ( clk ), .rnd ({Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380], Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370]}), .outt ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, n2357}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2527 ( .ina ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, n2359}), .inb ({new_AGEMA_signal_18401, new_AGEMA_signal_18399, new_AGEMA_signal_18397, new_AGEMA_signal_18395, new_AGEMA_signal_18393}), .clk ( clk ), .rnd ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390], Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385]}), .outt ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, n2360}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2534 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2674}), .clk ( clk ), .rnd ({Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410], Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .outt ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, n2369}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2536 ( .ina ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, n2371}), .inb ({new_AGEMA_signal_18291, new_AGEMA_signal_18289, new_AGEMA_signal_18287, new_AGEMA_signal_18285, new_AGEMA_signal_18283}), .clk ( clk ), .rnd ({Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420], Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415]}), .outt ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2372}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2539 ( .ina ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2576}), .inb ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2376}), .clk ( clk ), .rnd ({Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440], Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430]}), .outt ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, n2377}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2544 ( .ina ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .inb ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, n2415}), .clk ( clk ), .rnd ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450], Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445]}), .outt ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, n2467}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2545 ( .ina ({new_AGEMA_signal_18411, new_AGEMA_signal_18409, new_AGEMA_signal_18407, new_AGEMA_signal_18405, new_AGEMA_signal_18403}), .inb ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2383}), .clk ( clk ), .rnd ({Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470], Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .outt ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, n2385}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2546 ( .ina ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480], Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475]}), .outt ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2384}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2548 ( .ina ({new_AGEMA_signal_18041, new_AGEMA_signal_18039, new_AGEMA_signal_18037, new_AGEMA_signal_18035, new_AGEMA_signal_18033}), .inb ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2429}), .clk ( clk ), .rnd ({Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500], Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490]}), .outt ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2386}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2552 ( .ina ({new_AGEMA_signal_18251, new_AGEMA_signal_18249, new_AGEMA_signal_18247, new_AGEMA_signal_18245, new_AGEMA_signal_18243}), .inb ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, n2647}), .clk ( clk ), .rnd ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510], Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505]}), .outt ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, n2394}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2553 ( .ina ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .inb ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .clk ( clk ), .rnd ({Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530], Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .outt ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, n2391}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2554 ( .ina ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2505}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540], Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535]}), .outt ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, n2390}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2559 ( .ina ({new_AGEMA_signal_18181, new_AGEMA_signal_18179, new_AGEMA_signal_18177, new_AGEMA_signal_18175, new_AGEMA_signal_18173}), .inb ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2700}), .clk ( clk ), .rnd ({Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560], Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550]}), .outt ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2396}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2562 ( .ina ({new_AGEMA_signal_18421, new_AGEMA_signal_18419, new_AGEMA_signal_18417, new_AGEMA_signal_18415, new_AGEMA_signal_18413}), .inb ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2438}), .clk ( clk ), .rnd ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570], Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565]}), .outt ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, n2406}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2565 ( .ina ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, n2594}), .inb ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, n2402}), .clk ( clk ), .rnd ({Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590], Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .outt ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, n2403}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2569 ( .ina ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, n2407}), .inb ({new_AGEMA_signal_18221, new_AGEMA_signal_18219, new_AGEMA_signal_18217, new_AGEMA_signal_18215, new_AGEMA_signal_18213}), .clk ( clk ), .rnd ({Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600], Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595]}), .outt ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, n2408}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2573 ( .ina ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, n2412}), .inb ({new_AGEMA_signal_18301, new_AGEMA_signal_18299, new_AGEMA_signal_18297, new_AGEMA_signal_18295, new_AGEMA_signal_18293}), .clk ( clk ), .rnd ({Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620], Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610]}), .outt ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, n2574}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2574 ( .ina ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .inb ({new_AGEMA_signal_18121, new_AGEMA_signal_18119, new_AGEMA_signal_18117, new_AGEMA_signal_18115, new_AGEMA_signal_18113}), .clk ( clk ), .rnd ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630], Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625]}), .outt ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, n2413}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2577 ( .ina ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, n2415}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650], Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .outt ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2416}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2586 ( .ina ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, n2428}), .inb ({new_AGEMA_signal_18431, new_AGEMA_signal_18429, new_AGEMA_signal_18427, new_AGEMA_signal_18425, new_AGEMA_signal_18423}), .clk ( clk ), .rnd ({Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660], Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655]}), .outt ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, n2433}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2587 ( .ina ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .inb ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2429}), .clk ( clk ), .rnd ({Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680], Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670]}), .outt ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, n2689}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2591 ( .ina ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, n2647}), .inb ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}), .clk ( clk ), .rnd ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690], Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685]}), .outt ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2434}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2595 ( .ina ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2438}), .inb ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2483}), .clk ( clk ), .rnd ({Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710], Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .outt ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, n2439}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2598 ( .ina ({new_AGEMA_signal_18411, new_AGEMA_signal_18409, new_AGEMA_signal_18407, new_AGEMA_signal_18405, new_AGEMA_signal_18403}), .inb ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n2540}), .clk ( clk ), .rnd ({Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720], Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715]}), .outt ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, n2445}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2600 ( .ina ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2690}), .inb ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, n2443}), .clk ( clk ), .rnd ({Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740], Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730]}), .outt ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2444}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2602 ( .ina ({new_AGEMA_signal_17991, new_AGEMA_signal_17989, new_AGEMA_signal_17987, new_AGEMA_signal_17985, new_AGEMA_signal_17983}), .inb ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, n2446}), .clk ( clk ), .rnd ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750], Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745]}), .outt ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, n2447}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2607 ( .ina ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}), .inb ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, n2693}), .clk ( clk ), .rnd ({Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770], Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .outt ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, n2454}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2617 ( .ina ({new_AGEMA_signal_18191, new_AGEMA_signal_18189, new_AGEMA_signal_18187, new_AGEMA_signal_18185, new_AGEMA_signal_18183}), .inb ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, n2464}), .clk ( clk ), .rnd ({Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780], Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775]}), .outt ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2465}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2622 ( .ina ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2576}), .clk ( clk ), .rnd ({Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800], Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790]}), .outt ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, n2470}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2626 ( .ina ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, new_AGEMA_signal_1618, n2473}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, n2472}), .clk ( clk ), .rnd ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810], Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805]}), .outt ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, n2476}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2633 ( .ina ({new_AGEMA_signal_18441, new_AGEMA_signal_18439, new_AGEMA_signal_18437, new_AGEMA_signal_18435, new_AGEMA_signal_18433}), .inb ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2480}), .clk ( clk ), .rnd ({Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830], Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .outt ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, n2481}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2639 ( .ina ({new_AGEMA_signal_18451, new_AGEMA_signal_18449, new_AGEMA_signal_18447, new_AGEMA_signal_18445, new_AGEMA_signal_18443}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840], Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835]}), .outt ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, n2486}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2642 ( .ina ({new_AGEMA_signal_18321, new_AGEMA_signal_18319, new_AGEMA_signal_18317, new_AGEMA_signal_18315, new_AGEMA_signal_18313}), .inb ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, n2488}), .clk ( clk ), .rnd ({Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860], Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850]}), .outt ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2489}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2645 ( .ina ({new_AGEMA_signal_18461, new_AGEMA_signal_18459, new_AGEMA_signal_18457, new_AGEMA_signal_18455, new_AGEMA_signal_18453}), .inb ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2492}), .clk ( clk ), .rnd ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870], Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865]}), .outt ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, n2497}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2646 ( .ina ({new_AGEMA_signal_18471, new_AGEMA_signal_18469, new_AGEMA_signal_18467, new_AGEMA_signal_18465, new_AGEMA_signal_18463}), .inb ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2700}), .clk ( clk ), .rnd ({Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890], Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .outt ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, n2495}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2647 ( .ina ({new_AGEMA_signal_18201, new_AGEMA_signal_18199, new_AGEMA_signal_18197, new_AGEMA_signal_18195, new_AGEMA_signal_18193}), .inb ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2625}), .clk ( clk ), .rnd ({Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900], Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895]}), .outt ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, n2494}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2650 ( .ina ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2498}), .inb ({new_AGEMA_signal_17911, new_AGEMA_signal_17909, new_AGEMA_signal_17907, new_AGEMA_signal_17905, new_AGEMA_signal_17903}), .clk ( clk ), .rnd ({Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920], Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910]}), .outt ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2499}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2653 ( .ina ({new_AGEMA_signal_17911, new_AGEMA_signal_17909, new_AGEMA_signal_17907, new_AGEMA_signal_17905, new_AGEMA_signal_17903}), .inb ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2674}), .clk ( clk ), .rnd ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930], Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925]}), .outt ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2503}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2655 ( .ins ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2505}), .ina ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .clk ( clk ), .rnd ({Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950], Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .outt ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, n2506}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2662 ( .ina ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2662}), .inb ({new_AGEMA_signal_18021, new_AGEMA_signal_18019, new_AGEMA_signal_18017, new_AGEMA_signal_18015, new_AGEMA_signal_18013}), .clk ( clk ), .rnd ({Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960], Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955]}), .outt ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n2518}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2663 ( .ina ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2720}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980], Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970]}), .outt ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, n2517}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2666 ( .ina ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, n2520}), .inb ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .clk ( clk ), .rnd ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990], Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985]}), .outt ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, n2523}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2668 ( .ina ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2774}), .inb ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, n2521}), .clk ( clk ), .rnd ({Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010], Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .outt ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, n2522}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2675 ( .ina ({new_AGEMA_signal_18021, new_AGEMA_signal_18019, new_AGEMA_signal_18017, new_AGEMA_signal_18015, new_AGEMA_signal_18013}), .inb ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, n2531}), .clk ( clk ), .rnd ({Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020], Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015]}), .outt ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n2532}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2677 ( .ina ({new_AGEMA_signal_17861, new_AGEMA_signal_17859, new_AGEMA_signal_17857, new_AGEMA_signal_17855, new_AGEMA_signal_17853}), .inb ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2533}), .clk ( clk ), .rnd ({Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040], Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030]}), .outt ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, n2534}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2681 ( .ina ({new_AGEMA_signal_18481, new_AGEMA_signal_18479, new_AGEMA_signal_18477, new_AGEMA_signal_18475, new_AGEMA_signal_18473}), .inb ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n2540}), .clk ( clk ), .rnd ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050], Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045]}), .outt ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, n2542}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2683 ( .ina ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2545}), .inb ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, n2544}), .clk ( clk ), .rnd ({Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070], Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .outt ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2546}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2687 ( .ina ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, n2673}), .inb ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .clk ( clk ), .rnd ({Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080], Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075]}), .outt ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, n2551}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2690 ( .ina ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, n2553}), .inb ({new_AGEMA_signal_18491, new_AGEMA_signal_18489, new_AGEMA_signal_18487, new_AGEMA_signal_18485, new_AGEMA_signal_18483}), .clk ( clk ), .rnd ({Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100], Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090]}), .outt ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, n2558}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2692 ( .ina ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, n2555}), .inb ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, n2554}), .clk ( clk ), .rnd ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110], Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105]}), .outt ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2556}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2696 ( .ina ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n2561}), .inb ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2560}), .clk ( clk ), .rnd ({Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130], Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .outt ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, n2566}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2697 ( .ina ({new_AGEMA_signal_18501, new_AGEMA_signal_18499, new_AGEMA_signal_18497, new_AGEMA_signal_18495, new_AGEMA_signal_18493}), .inb ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, n2562}), .clk ( clk ), .rnd ({Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140], Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135]}), .outt ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, n2715}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2703 ( .ina ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2572}), .inb ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2571}), .clk ( clk ), .rnd ({Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160], Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150]}), .outt ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2573}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2705 ( .ina ({new_AGEMA_signal_18421, new_AGEMA_signal_18419, new_AGEMA_signal_18417, new_AGEMA_signal_18415, new_AGEMA_signal_18413}), .inb ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2754}), .clk ( clk ), .rnd ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170], Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165]}), .outt ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, n2585}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2706 ( .ina ({new_AGEMA_signal_18311, new_AGEMA_signal_18309, new_AGEMA_signal_18307, new_AGEMA_signal_18305, new_AGEMA_signal_18303}), .inb ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, n2627}), .clk ( clk ), .rnd ({Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190], Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .outt ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, n2581}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2707 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, n2575}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200], Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195]}), .outt ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, n2579}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2708 ( .ina ({new_AGEMA_signal_18471, new_AGEMA_signal_18469, new_AGEMA_signal_18467, new_AGEMA_signal_18465, new_AGEMA_signal_18463}), .inb ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2576}), .clk ( clk ), .rnd ({Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220], Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210]}), .outt ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, n2578}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2711 ( .ina ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2625}), .inb ({new_AGEMA_signal_18271, new_AGEMA_signal_18269, new_AGEMA_signal_18267, new_AGEMA_signal_18265, new_AGEMA_signal_18263}), .clk ( clk ), .rnd ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230], Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225]}), .outt ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2582}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2715 ( .ina ({new_AGEMA_signal_17951, new_AGEMA_signal_17949, new_AGEMA_signal_17947, new_AGEMA_signal_17945, new_AGEMA_signal_17943}), .inb ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2586}), .clk ( clk ), .rnd ({Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250], Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .outt ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, n2588}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2719 ( .ina ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, n2594}), .inb ({new_AGEMA_signal_18421, new_AGEMA_signal_18419, new_AGEMA_signal_18417, new_AGEMA_signal_18415, new_AGEMA_signal_18413}), .clk ( clk ), .rnd ({Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260], Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255]}), .outt ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, n2607}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2722 ( .ina ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, n2597}), .inb ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, n2596}), .clk ( clk ), .rnd ({Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280], Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270]}), .outt ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, n2605}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2724 ( .ina ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2598}), .inb ({new_AGEMA_signal_18511, new_AGEMA_signal_18509, new_AGEMA_signal_18507, new_AGEMA_signal_18505, new_AGEMA_signal_18503}), .clk ( clk ), .rnd ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290], Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285]}), .outt ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2603}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2726 ( .ina ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, new_AGEMA_signal_1258, n2599}), .inb ({new_AGEMA_signal_18301, new_AGEMA_signal_18299, new_AGEMA_signal_18297, new_AGEMA_signal_18295, new_AGEMA_signal_18293}), .clk ( clk ), .rnd ({Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310], Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .outt ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, n2601}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2733 ( .ina ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, n2610}), .inb ({new_AGEMA_signal_18261, new_AGEMA_signal_18259, new_AGEMA_signal_18257, new_AGEMA_signal_18255, new_AGEMA_signal_18253}), .clk ( clk ), .rnd ({Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320], Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315]}), .outt ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, n2620}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2736 ( .ina ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2614}), .inb ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, n2613}), .clk ( clk ), .rnd ({Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340], Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330]}), .outt ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, n2618}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2743 ( .ina ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .inb ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2625}), .clk ( clk ), .rnd ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350], Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345]}), .outt ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2626}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2746 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2631}), .inb ({new_AGEMA_signal_18091, new_AGEMA_signal_18089, new_AGEMA_signal_18087, new_AGEMA_signal_18085, new_AGEMA_signal_18083}), .clk ( clk ), .rnd ({Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370], Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .outt ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, n2632}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2752 ( .ina ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2784}), .inb ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2642}), .clk ( clk ), .rnd ({Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380], Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375]}), .outt ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, n2644}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2754 ( .ina ({new_AGEMA_signal_17901, new_AGEMA_signal_17899, new_AGEMA_signal_17897, new_AGEMA_signal_17895, new_AGEMA_signal_17893}), .inb ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, n2645}), .clk ( clk ), .rnd ({Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400], Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390]}), .outt ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, n2646}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2758 ( .ina ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2651}), .inb ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, n2650}), .clk ( clk ), .rnd ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410], Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405]}), .outt ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, n2653}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2760 ( .ina ({new_AGEMA_signal_18301, new_AGEMA_signal_18299, new_AGEMA_signal_18297, new_AGEMA_signal_18295, new_AGEMA_signal_18293}), .inb ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2654}), .clk ( clk ), .rnd ({Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430], Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .outt ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, n2655}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2764 ( .ina ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2662}), .inb ({new_AGEMA_signal_18321, new_AGEMA_signal_18319, new_AGEMA_signal_18317, new_AGEMA_signal_18315, new_AGEMA_signal_18313}), .clk ( clk ), .rnd ({Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440], Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435]}), .outt ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, n2663}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2770 ( .ina ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, n2673}), .inb ({new_AGEMA_signal_18271, new_AGEMA_signal_18269, new_AGEMA_signal_18267, new_AGEMA_signal_18265, new_AGEMA_signal_18263}), .clk ( clk ), .rnd ({Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460], Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450]}), .outt ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2675}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2772 ( .ina ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2677}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2676}), .clk ( clk ), .rnd ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470], Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465]}), .outt ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, n2678}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2780 ( .ina ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2690}), .inb ({new_AGEMA_signal_18311, new_AGEMA_signal_18309, new_AGEMA_signal_18307, new_AGEMA_signal_18305, new_AGEMA_signal_18303}), .clk ( clk ), .rnd ({Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490], Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .outt ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, new_AGEMA_signal_2342, n2691}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2782 ( .ina ({new_AGEMA_signal_18341, new_AGEMA_signal_18339, new_AGEMA_signal_18337, new_AGEMA_signal_18335, new_AGEMA_signal_18333}), .inb ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, n2693}), .clk ( clk ), .rnd ({Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500], Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495]}), .outt ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, n2695}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2785 ( .ina ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2700}), .inb ({new_AGEMA_signal_18501, new_AGEMA_signal_18499, new_AGEMA_signal_18497, new_AGEMA_signal_18495, new_AGEMA_signal_18493}), .clk ( clk ), .rnd ({Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520], Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510]}), .outt ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2701}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2791 ( .ina ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, n2711}), .inb ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, n2710}), .clk ( clk ), .rnd ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530], Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525]}), .outt ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, n2717}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2796 ( .ina ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2720}), .inb ({new_AGEMA_signal_18211, new_AGEMA_signal_18209, new_AGEMA_signal_18207, new_AGEMA_signal_18205, new_AGEMA_signal_18203}), .clk ( clk ), .rnd ({Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550], Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .outt ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, n2729}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2798 ( .ina ({new_AGEMA_signal_18041, new_AGEMA_signal_18039, new_AGEMA_signal_18037, new_AGEMA_signal_18035, new_AGEMA_signal_18033}), .inb ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, n2722}), .clk ( clk ), .rnd ({Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560], Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555]}), .outt ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2727}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2803 ( .ina ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, n2732}), .inb ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2731}), .clk ( clk ), .rnd ({Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580], Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570]}), .outt ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2733}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2807 ( .ina ({new_AGEMA_signal_18521, new_AGEMA_signal_18519, new_AGEMA_signal_18517, new_AGEMA_signal_18515, new_AGEMA_signal_18513}), .inb ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, n2738}), .clk ( clk ), .rnd ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590], Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585]}), .outt ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, n2740}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2812 ( .ina ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, n2748}), .inb ({new_AGEMA_signal_17861, new_AGEMA_signal_17859, new_AGEMA_signal_17857, new_AGEMA_signal_17855, new_AGEMA_signal_17853}), .clk ( clk ), .rnd ({Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610], Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .outt ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2749}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2815 ( .ina ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2754}), .inb ({new_AGEMA_signal_18061, new_AGEMA_signal_18059, new_AGEMA_signal_18057, new_AGEMA_signal_18055, new_AGEMA_signal_18053}), .clk ( clk ), .rnd ({Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620], Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615]}), .outt ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2757}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2816 ( .ina ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, new_AGEMA_signal_1294, n2755}), .inb ({new_AGEMA_signal_18531, new_AGEMA_signal_18529, new_AGEMA_signal_18527, new_AGEMA_signal_18525, new_AGEMA_signal_18523}), .clk ( clk ), .rnd ({Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640], Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630]}), .outt ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, n2756}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2819 ( .ina ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2761}), .inb ({new_AGEMA_signal_18351, new_AGEMA_signal_18349, new_AGEMA_signal_18347, new_AGEMA_signal_18345, new_AGEMA_signal_18343}), .clk ( clk ), .rnd ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650], Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645]}), .outt ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, n2762}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2823 ( .ina ({new_AGEMA_signal_17861, new_AGEMA_signal_17859, new_AGEMA_signal_17857, new_AGEMA_signal_17855, new_AGEMA_signal_17853}), .inb ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, n2768}), .clk ( clk ), .rnd ({Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670], Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .outt ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, n2770}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2825 ( .ina ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, new_AGEMA_signal_1910, n2773}), .inb ({new_AGEMA_signal_18531, new_AGEMA_signal_18529, new_AGEMA_signal_18527, new_AGEMA_signal_18525, new_AGEMA_signal_18523}), .clk ( clk ), .rnd ({Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680], Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675]}), .outt ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2776}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2826 ( .ina ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2774}), .inb ({new_AGEMA_signal_17871, new_AGEMA_signal_17869, new_AGEMA_signal_17867, new_AGEMA_signal_17865, new_AGEMA_signal_17863}), .clk ( clk ), .rnd ({Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700], Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690]}), .outt ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, n2775}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2830 ( .ina ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, n2782}), .inb ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2781}), .clk ( clk ), .rnd ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710], Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705]}), .outt ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2783}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2836 ( .ina ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, n2794}), .inb ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2793}), .clk ( clk ), .rnd ({Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730], Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720]}), .outt ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2795}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2845 ( .ina ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, n2812}), .inb ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2811}), .clk ( clk ), .rnd ({Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740], Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735]}), .outt ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, n2814}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2848 ( .ina ({new_AGEMA_signal_17981, new_AGEMA_signal_17979, new_AGEMA_signal_17977, new_AGEMA_signal_17975, new_AGEMA_signal_17973}), .inb ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2817}), .clk ( clk ), .rnd ({Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760], Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750]}), .outt ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_18532 ), .Q ( new_AGEMA_signal_18533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_18534 ), .Q ( new_AGEMA_signal_18535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_18536 ), .Q ( new_AGEMA_signal_18537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_18538 ), .Q ( new_AGEMA_signal_18539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_18540 ), .Q ( new_AGEMA_signal_18541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_18542 ), .Q ( new_AGEMA_signal_18543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_18544 ), .Q ( new_AGEMA_signal_18545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_18546 ), .Q ( new_AGEMA_signal_18547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_18548 ), .Q ( new_AGEMA_signal_18549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_18550 ), .Q ( new_AGEMA_signal_18551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_18554 ), .Q ( new_AGEMA_signal_18555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_18558 ), .Q ( new_AGEMA_signal_18559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_18562 ), .Q ( new_AGEMA_signal_18563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_18566 ), .Q ( new_AGEMA_signal_18567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_18570 ), .Q ( new_AGEMA_signal_18571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_18572 ), .Q ( new_AGEMA_signal_18573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_18574 ), .Q ( new_AGEMA_signal_18575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_18576 ), .Q ( new_AGEMA_signal_18577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_18578 ), .Q ( new_AGEMA_signal_18579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_18580 ), .Q ( new_AGEMA_signal_18581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_18582 ), .Q ( new_AGEMA_signal_18583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_18584 ), .Q ( new_AGEMA_signal_18585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_18586 ), .Q ( new_AGEMA_signal_18587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_18588 ), .Q ( new_AGEMA_signal_18589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_18590 ), .Q ( new_AGEMA_signal_18591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_18592 ), .Q ( new_AGEMA_signal_18593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_18594 ), .Q ( new_AGEMA_signal_18595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_18596 ), .Q ( new_AGEMA_signal_18597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_18598 ), .Q ( new_AGEMA_signal_18599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_18600 ), .Q ( new_AGEMA_signal_18601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_18602 ), .Q ( new_AGEMA_signal_18603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_18604 ), .Q ( new_AGEMA_signal_18605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_18606 ), .Q ( new_AGEMA_signal_18607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_18608 ), .Q ( new_AGEMA_signal_18609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_18610 ), .Q ( new_AGEMA_signal_18611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_18612 ), .Q ( new_AGEMA_signal_18613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_18614 ), .Q ( new_AGEMA_signal_18615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_18616 ), .Q ( new_AGEMA_signal_18617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_18618 ), .Q ( new_AGEMA_signal_18619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_18620 ), .Q ( new_AGEMA_signal_18621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_18622 ), .Q ( new_AGEMA_signal_18623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_18624 ), .Q ( new_AGEMA_signal_18625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_18626 ), .Q ( new_AGEMA_signal_18627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_18628 ), .Q ( new_AGEMA_signal_18629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_18630 ), .Q ( new_AGEMA_signal_18631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_18632 ), .Q ( new_AGEMA_signal_18633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_18634 ), .Q ( new_AGEMA_signal_18635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_18636 ), .Q ( new_AGEMA_signal_18637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_18638 ), .Q ( new_AGEMA_signal_18639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_18640 ), .Q ( new_AGEMA_signal_18641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_18642 ), .Q ( new_AGEMA_signal_18643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_18644 ), .Q ( new_AGEMA_signal_18645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_18646 ), .Q ( new_AGEMA_signal_18647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_18648 ), .Q ( new_AGEMA_signal_18649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_18650 ), .Q ( new_AGEMA_signal_18651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_18652 ), .Q ( new_AGEMA_signal_18653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_18654 ), .Q ( new_AGEMA_signal_18655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_18656 ), .Q ( new_AGEMA_signal_18657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_18658 ), .Q ( new_AGEMA_signal_18659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_18660 ), .Q ( new_AGEMA_signal_18661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_18662 ), .Q ( new_AGEMA_signal_18663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_18664 ), .Q ( new_AGEMA_signal_18665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_18666 ), .Q ( new_AGEMA_signal_18667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_18668 ), .Q ( new_AGEMA_signal_18669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_18670 ), .Q ( new_AGEMA_signal_18671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_18672 ), .Q ( new_AGEMA_signal_18673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_18674 ), .Q ( new_AGEMA_signal_18675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_18676 ), .Q ( new_AGEMA_signal_18677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_18678 ), .Q ( new_AGEMA_signal_18679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_18680 ), .Q ( new_AGEMA_signal_18681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_18684 ), .Q ( new_AGEMA_signal_18685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_18688 ), .Q ( new_AGEMA_signal_18689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_18692 ), .Q ( new_AGEMA_signal_18693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_18696 ), .Q ( new_AGEMA_signal_18697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_18700 ), .Q ( new_AGEMA_signal_18701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_18702 ), .Q ( new_AGEMA_signal_18703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_18704 ), .Q ( new_AGEMA_signal_18705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_18706 ), .Q ( new_AGEMA_signal_18707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_18708 ), .Q ( new_AGEMA_signal_18709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_18710 ), .Q ( new_AGEMA_signal_18711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_18712 ), .Q ( new_AGEMA_signal_18713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_18714 ), .Q ( new_AGEMA_signal_18715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_18716 ), .Q ( new_AGEMA_signal_18717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_18718 ), .Q ( new_AGEMA_signal_18719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_18720 ), .Q ( new_AGEMA_signal_18721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_18722 ), .Q ( new_AGEMA_signal_18723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_18724 ), .Q ( new_AGEMA_signal_18725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_18726 ), .Q ( new_AGEMA_signal_18727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_18728 ), .Q ( new_AGEMA_signal_18729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_18730 ), .Q ( new_AGEMA_signal_18731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_18732 ), .Q ( new_AGEMA_signal_18733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_18734 ), .Q ( new_AGEMA_signal_18735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_18736 ), .Q ( new_AGEMA_signal_18737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_18738 ), .Q ( new_AGEMA_signal_18739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_18740 ), .Q ( new_AGEMA_signal_18741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_18742 ), .Q ( new_AGEMA_signal_18743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_18744 ), .Q ( new_AGEMA_signal_18745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_18746 ), .Q ( new_AGEMA_signal_18747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_18748 ), .Q ( new_AGEMA_signal_18749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_18750 ), .Q ( new_AGEMA_signal_18751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_18752 ), .Q ( new_AGEMA_signal_18753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_18754 ), .Q ( new_AGEMA_signal_18755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_18756 ), .Q ( new_AGEMA_signal_18757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_18758 ), .Q ( new_AGEMA_signal_18759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_18760 ), .Q ( new_AGEMA_signal_18761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_18762 ), .Q ( new_AGEMA_signal_18763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_18764 ), .Q ( new_AGEMA_signal_18765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_18766 ), .Q ( new_AGEMA_signal_18767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_18768 ), .Q ( new_AGEMA_signal_18769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_18770 ), .Q ( new_AGEMA_signal_18771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_18774 ), .Q ( new_AGEMA_signal_18775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_18778 ), .Q ( new_AGEMA_signal_18779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_18782 ), .Q ( new_AGEMA_signal_18783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_18786 ), .Q ( new_AGEMA_signal_18787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_18790 ), .Q ( new_AGEMA_signal_18791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_18792 ), .Q ( new_AGEMA_signal_18793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_18794 ), .Q ( new_AGEMA_signal_18795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_18796 ), .Q ( new_AGEMA_signal_18797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_18798 ), .Q ( new_AGEMA_signal_18799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_18800 ), .Q ( new_AGEMA_signal_18801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_18802 ), .Q ( new_AGEMA_signal_18803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_18804 ), .Q ( new_AGEMA_signal_18805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_18806 ), .Q ( new_AGEMA_signal_18807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_18808 ), .Q ( new_AGEMA_signal_18809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_18810 ), .Q ( new_AGEMA_signal_18811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_18812 ), .Q ( new_AGEMA_signal_18813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_18814 ), .Q ( new_AGEMA_signal_18815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_18816 ), .Q ( new_AGEMA_signal_18817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_18818 ), .Q ( new_AGEMA_signal_18819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_18820 ), .Q ( new_AGEMA_signal_18821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_18822 ), .Q ( new_AGEMA_signal_18823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_18824 ), .Q ( new_AGEMA_signal_18825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_18826 ), .Q ( new_AGEMA_signal_18827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_18828 ), .Q ( new_AGEMA_signal_18829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_18830 ), .Q ( new_AGEMA_signal_18831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_18832 ), .Q ( new_AGEMA_signal_18833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_18834 ), .Q ( new_AGEMA_signal_18835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_18836 ), .Q ( new_AGEMA_signal_18837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_18838 ), .Q ( new_AGEMA_signal_18839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_18840 ), .Q ( new_AGEMA_signal_18841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_18844 ), .Q ( new_AGEMA_signal_18845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_18848 ), .Q ( new_AGEMA_signal_18849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_18852 ), .Q ( new_AGEMA_signal_18853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_18856 ), .Q ( new_AGEMA_signal_18857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_18860 ), .Q ( new_AGEMA_signal_18861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_18862 ), .Q ( new_AGEMA_signal_18863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_18864 ), .Q ( new_AGEMA_signal_18865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_18866 ), .Q ( new_AGEMA_signal_18867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_18868 ), .Q ( new_AGEMA_signal_18869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_18870 ), .Q ( new_AGEMA_signal_18871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_18872 ), .Q ( new_AGEMA_signal_18873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_18874 ), .Q ( new_AGEMA_signal_18875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_18876 ), .Q ( new_AGEMA_signal_18877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_18878 ), .Q ( new_AGEMA_signal_18879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_18880 ), .Q ( new_AGEMA_signal_18881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_18882 ), .Q ( new_AGEMA_signal_18883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_18884 ), .Q ( new_AGEMA_signal_18885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_18886 ), .Q ( new_AGEMA_signal_18887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_18888 ), .Q ( new_AGEMA_signal_18889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_18890 ), .Q ( new_AGEMA_signal_18891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_18894 ), .Q ( new_AGEMA_signal_18895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_18898 ), .Q ( new_AGEMA_signal_18899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_18902 ), .Q ( new_AGEMA_signal_18903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_18906 ), .Q ( new_AGEMA_signal_18907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_18910 ), .Q ( new_AGEMA_signal_18911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_18912 ), .Q ( new_AGEMA_signal_18913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_18914 ), .Q ( new_AGEMA_signal_18915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_18916 ), .Q ( new_AGEMA_signal_18917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_18918 ), .Q ( new_AGEMA_signal_18919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_18920 ), .Q ( new_AGEMA_signal_18921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_18922 ), .Q ( new_AGEMA_signal_18923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_18924 ), .Q ( new_AGEMA_signal_18925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_18926 ), .Q ( new_AGEMA_signal_18927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_18928 ), .Q ( new_AGEMA_signal_18929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_18930 ), .Q ( new_AGEMA_signal_18931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_18932 ), .Q ( new_AGEMA_signal_18933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_18934 ), .Q ( new_AGEMA_signal_18935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_18936 ), .Q ( new_AGEMA_signal_18937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_18938 ), .Q ( new_AGEMA_signal_18939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_18940 ), .Q ( new_AGEMA_signal_18941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_18944 ), .Q ( new_AGEMA_signal_18945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_18948 ), .Q ( new_AGEMA_signal_18949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_18952 ), .Q ( new_AGEMA_signal_18953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_18956 ), .Q ( new_AGEMA_signal_18957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_18960 ), .Q ( new_AGEMA_signal_18961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_18962 ), .Q ( new_AGEMA_signal_18963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_18964 ), .Q ( new_AGEMA_signal_18965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_18966 ), .Q ( new_AGEMA_signal_18967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_18968 ), .Q ( new_AGEMA_signal_18969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_18970 ), .Q ( new_AGEMA_signal_18971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_18972 ), .Q ( new_AGEMA_signal_18973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_18974 ), .Q ( new_AGEMA_signal_18975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_18976 ), .Q ( new_AGEMA_signal_18977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_18978 ), .Q ( new_AGEMA_signal_18979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_18980 ), .Q ( new_AGEMA_signal_18981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_18982 ), .Q ( new_AGEMA_signal_18983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_18984 ), .Q ( new_AGEMA_signal_18985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_18986 ), .Q ( new_AGEMA_signal_18987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_18988 ), .Q ( new_AGEMA_signal_18989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_18990 ), .Q ( new_AGEMA_signal_18991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_18992 ), .Q ( new_AGEMA_signal_18993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_18994 ), .Q ( new_AGEMA_signal_18995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_18996 ), .Q ( new_AGEMA_signal_18997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_18998 ), .Q ( new_AGEMA_signal_18999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_19000 ), .Q ( new_AGEMA_signal_19001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_19002 ), .Q ( new_AGEMA_signal_19003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_19004 ), .Q ( new_AGEMA_signal_19005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_19006 ), .Q ( new_AGEMA_signal_19007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_19008 ), .Q ( new_AGEMA_signal_19009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_19010 ), .Q ( new_AGEMA_signal_19011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_19012 ), .Q ( new_AGEMA_signal_19013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_19014 ), .Q ( new_AGEMA_signal_19015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_19016 ), .Q ( new_AGEMA_signal_19017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_19018 ), .Q ( new_AGEMA_signal_19019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_19020 ), .Q ( new_AGEMA_signal_19021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_19022 ), .Q ( new_AGEMA_signal_19023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_19024 ), .Q ( new_AGEMA_signal_19025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_19026 ), .Q ( new_AGEMA_signal_19027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_19028 ), .Q ( new_AGEMA_signal_19029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_19030 ), .Q ( new_AGEMA_signal_19031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_19032 ), .Q ( new_AGEMA_signal_19033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_19034 ), .Q ( new_AGEMA_signal_19035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_19036 ), .Q ( new_AGEMA_signal_19037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_19038 ), .Q ( new_AGEMA_signal_19039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_19040 ), .Q ( new_AGEMA_signal_19041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_19042 ), .Q ( new_AGEMA_signal_19043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_19044 ), .Q ( new_AGEMA_signal_19045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_19046 ), .Q ( new_AGEMA_signal_19047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_19048 ), .Q ( new_AGEMA_signal_19049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_19050 ), .Q ( new_AGEMA_signal_19051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_19052 ), .Q ( new_AGEMA_signal_19053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_19054 ), .Q ( new_AGEMA_signal_19055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_19056 ), .Q ( new_AGEMA_signal_19057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_19058 ), .Q ( new_AGEMA_signal_19059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_19060 ), .Q ( new_AGEMA_signal_19061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_19062 ), .Q ( new_AGEMA_signal_19063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_19064 ), .Q ( new_AGEMA_signal_19065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_19066 ), .Q ( new_AGEMA_signal_19067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_19068 ), .Q ( new_AGEMA_signal_19069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_19070 ), .Q ( new_AGEMA_signal_19071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_19072 ), .Q ( new_AGEMA_signal_19073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_19074 ), .Q ( new_AGEMA_signal_19075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_19076 ), .Q ( new_AGEMA_signal_19077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_19078 ), .Q ( new_AGEMA_signal_19079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_19080 ), .Q ( new_AGEMA_signal_19081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_19082 ), .Q ( new_AGEMA_signal_19083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_19084 ), .Q ( new_AGEMA_signal_19085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_19086 ), .Q ( new_AGEMA_signal_19087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_19088 ), .Q ( new_AGEMA_signal_19089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_19090 ), .Q ( new_AGEMA_signal_19091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_19092 ), .Q ( new_AGEMA_signal_19093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_19094 ), .Q ( new_AGEMA_signal_19095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_19096 ), .Q ( new_AGEMA_signal_19097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_19098 ), .Q ( new_AGEMA_signal_19099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_19100 ), .Q ( new_AGEMA_signal_19101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_19102 ), .Q ( new_AGEMA_signal_19103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_19104 ), .Q ( new_AGEMA_signal_19105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_19106 ), .Q ( new_AGEMA_signal_19107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_19108 ), .Q ( new_AGEMA_signal_19109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_19110 ), .Q ( new_AGEMA_signal_19111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_19112 ), .Q ( new_AGEMA_signal_19113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_19114 ), .Q ( new_AGEMA_signal_19115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_19116 ), .Q ( new_AGEMA_signal_19117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_19118 ), .Q ( new_AGEMA_signal_19119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_19120 ), .Q ( new_AGEMA_signal_19121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_19122 ), .Q ( new_AGEMA_signal_19123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_19124 ), .Q ( new_AGEMA_signal_19125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_19126 ), .Q ( new_AGEMA_signal_19127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_19128 ), .Q ( new_AGEMA_signal_19129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_19130 ), .Q ( new_AGEMA_signal_19131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_19136 ), .Q ( new_AGEMA_signal_19137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_19142 ), .Q ( new_AGEMA_signal_19143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_19148 ), .Q ( new_AGEMA_signal_19149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_19154 ), .Q ( new_AGEMA_signal_19155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_19160 ), .Q ( new_AGEMA_signal_19161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_19162 ), .Q ( new_AGEMA_signal_19163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_19164 ), .Q ( new_AGEMA_signal_19165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_19166 ), .Q ( new_AGEMA_signal_19167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_19168 ), .Q ( new_AGEMA_signal_19169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_19170 ), .Q ( new_AGEMA_signal_19171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_19172 ), .Q ( new_AGEMA_signal_19173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_19174 ), .Q ( new_AGEMA_signal_19175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_19176 ), .Q ( new_AGEMA_signal_19177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_19178 ), .Q ( new_AGEMA_signal_19179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_19180 ), .Q ( new_AGEMA_signal_19181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_19182 ), .Q ( new_AGEMA_signal_19183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_19184 ), .Q ( new_AGEMA_signal_19185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_19186 ), .Q ( new_AGEMA_signal_19187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_19188 ), .Q ( new_AGEMA_signal_19189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_19190 ), .Q ( new_AGEMA_signal_19191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_19194 ), .Q ( new_AGEMA_signal_19195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_19198 ), .Q ( new_AGEMA_signal_19199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_19202 ), .Q ( new_AGEMA_signal_19203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_19206 ), .Q ( new_AGEMA_signal_19207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_19210 ), .Q ( new_AGEMA_signal_19211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_19212 ), .Q ( new_AGEMA_signal_19213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_19214 ), .Q ( new_AGEMA_signal_19215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_19216 ), .Q ( new_AGEMA_signal_19217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_19218 ), .Q ( new_AGEMA_signal_19219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_19220 ), .Q ( new_AGEMA_signal_19221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_19222 ), .Q ( new_AGEMA_signal_19223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_19224 ), .Q ( new_AGEMA_signal_19225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_19226 ), .Q ( new_AGEMA_signal_19227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_19228 ), .Q ( new_AGEMA_signal_19229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_19230 ), .Q ( new_AGEMA_signal_19231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_19232 ), .Q ( new_AGEMA_signal_19233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_19234 ), .Q ( new_AGEMA_signal_19235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_19236 ), .Q ( new_AGEMA_signal_19237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_19238 ), .Q ( new_AGEMA_signal_19239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_19240 ), .Q ( new_AGEMA_signal_19241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_19244 ), .Q ( new_AGEMA_signal_19245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_19248 ), .Q ( new_AGEMA_signal_19249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_19252 ), .Q ( new_AGEMA_signal_19253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_19256 ), .Q ( new_AGEMA_signal_19257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_19260 ), .Q ( new_AGEMA_signal_19261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_19262 ), .Q ( new_AGEMA_signal_19263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_19264 ), .Q ( new_AGEMA_signal_19265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_19266 ), .Q ( new_AGEMA_signal_19267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_19268 ), .Q ( new_AGEMA_signal_19269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_19270 ), .Q ( new_AGEMA_signal_19271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_19272 ), .Q ( new_AGEMA_signal_19273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_19274 ), .Q ( new_AGEMA_signal_19275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_19276 ), .Q ( new_AGEMA_signal_19277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_19278 ), .Q ( new_AGEMA_signal_19279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_19280 ), .Q ( new_AGEMA_signal_19281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_19282 ), .Q ( new_AGEMA_signal_19283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_19284 ), .Q ( new_AGEMA_signal_19285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_19286 ), .Q ( new_AGEMA_signal_19287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_19288 ), .Q ( new_AGEMA_signal_19289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_19290 ), .Q ( new_AGEMA_signal_19291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_19292 ), .Q ( new_AGEMA_signal_19293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_19294 ), .Q ( new_AGEMA_signal_19295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_19296 ), .Q ( new_AGEMA_signal_19297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_19298 ), .Q ( new_AGEMA_signal_19299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_19300 ), .Q ( new_AGEMA_signal_19301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_19302 ), .Q ( new_AGEMA_signal_19303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_19304 ), .Q ( new_AGEMA_signal_19305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_19306 ), .Q ( new_AGEMA_signal_19307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_19308 ), .Q ( new_AGEMA_signal_19309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_19310 ), .Q ( new_AGEMA_signal_19311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_19312 ), .Q ( new_AGEMA_signal_19313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_19314 ), .Q ( new_AGEMA_signal_19315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_19316 ), .Q ( new_AGEMA_signal_19317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_19318 ), .Q ( new_AGEMA_signal_19319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_19320 ), .Q ( new_AGEMA_signal_19321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_19322 ), .Q ( new_AGEMA_signal_19323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_19324 ), .Q ( new_AGEMA_signal_19325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_19326 ), .Q ( new_AGEMA_signal_19327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_19328 ), .Q ( new_AGEMA_signal_19329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_19330 ), .Q ( new_AGEMA_signal_19331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_19334 ), .Q ( new_AGEMA_signal_19335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_19338 ), .Q ( new_AGEMA_signal_19339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_19342 ), .Q ( new_AGEMA_signal_19343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_19346 ), .Q ( new_AGEMA_signal_19347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_19350 ), .Q ( new_AGEMA_signal_19351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_19352 ), .Q ( new_AGEMA_signal_19353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_19354 ), .Q ( new_AGEMA_signal_19355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_19356 ), .Q ( new_AGEMA_signal_19357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_19358 ), .Q ( new_AGEMA_signal_19359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_19360 ), .Q ( new_AGEMA_signal_19361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_19362 ), .Q ( new_AGEMA_signal_19363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_19364 ), .Q ( new_AGEMA_signal_19365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_19366 ), .Q ( new_AGEMA_signal_19367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_19368 ), .Q ( new_AGEMA_signal_19369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_19370 ), .Q ( new_AGEMA_signal_19371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_19374 ), .Q ( new_AGEMA_signal_19375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_19378 ), .Q ( new_AGEMA_signal_19379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_19382 ), .Q ( new_AGEMA_signal_19383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C ( clk ), .D ( new_AGEMA_signal_19386 ), .Q ( new_AGEMA_signal_19387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C ( clk ), .D ( new_AGEMA_signal_19390 ), .Q ( new_AGEMA_signal_19391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C ( clk ), .D ( new_AGEMA_signal_19392 ), .Q ( new_AGEMA_signal_19393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C ( clk ), .D ( new_AGEMA_signal_19394 ), .Q ( new_AGEMA_signal_19395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C ( clk ), .D ( new_AGEMA_signal_19396 ), .Q ( new_AGEMA_signal_19397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C ( clk ), .D ( new_AGEMA_signal_19398 ), .Q ( new_AGEMA_signal_19399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C ( clk ), .D ( new_AGEMA_signal_19400 ), .Q ( new_AGEMA_signal_19401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C ( clk ), .D ( new_AGEMA_signal_19402 ), .Q ( new_AGEMA_signal_19403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C ( clk ), .D ( new_AGEMA_signal_19406 ), .Q ( new_AGEMA_signal_19407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C ( clk ), .D ( new_AGEMA_signal_19410 ), .Q ( new_AGEMA_signal_19411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C ( clk ), .D ( new_AGEMA_signal_19414 ), .Q ( new_AGEMA_signal_19415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C ( clk ), .D ( new_AGEMA_signal_19418 ), .Q ( new_AGEMA_signal_19419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C ( clk ), .D ( new_AGEMA_signal_19422 ), .Q ( new_AGEMA_signal_19423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C ( clk ), .D ( new_AGEMA_signal_19426 ), .Q ( new_AGEMA_signal_19427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C ( clk ), .D ( new_AGEMA_signal_19430 ), .Q ( new_AGEMA_signal_19431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C ( clk ), .D ( new_AGEMA_signal_19434 ), .Q ( new_AGEMA_signal_19435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C ( clk ), .D ( new_AGEMA_signal_19438 ), .Q ( new_AGEMA_signal_19439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C ( clk ), .D ( new_AGEMA_signal_19462 ), .Q ( new_AGEMA_signal_19463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C ( clk ), .D ( new_AGEMA_signal_19466 ), .Q ( new_AGEMA_signal_19467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C ( clk ), .D ( new_AGEMA_signal_19470 ), .Q ( new_AGEMA_signal_19471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C ( clk ), .D ( new_AGEMA_signal_19474 ), .Q ( new_AGEMA_signal_19475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C ( clk ), .D ( new_AGEMA_signal_19478 ), .Q ( new_AGEMA_signal_19479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C ( clk ), .D ( new_AGEMA_signal_19492 ), .Q ( new_AGEMA_signal_19493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C ( clk ), .D ( new_AGEMA_signal_19496 ), .Q ( new_AGEMA_signal_19497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C ( clk ), .D ( new_AGEMA_signal_19500 ), .Q ( new_AGEMA_signal_19501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C ( clk ), .D ( new_AGEMA_signal_19504 ), .Q ( new_AGEMA_signal_19505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C ( clk ), .D ( new_AGEMA_signal_19508 ), .Q ( new_AGEMA_signal_19509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C ( clk ), .D ( new_AGEMA_signal_19522 ), .Q ( new_AGEMA_signal_19523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C ( clk ), .D ( new_AGEMA_signal_19526 ), .Q ( new_AGEMA_signal_19527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C ( clk ), .D ( new_AGEMA_signal_19530 ), .Q ( new_AGEMA_signal_19531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C ( clk ), .D ( new_AGEMA_signal_19534 ), .Q ( new_AGEMA_signal_19535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C ( clk ), .D ( new_AGEMA_signal_19538 ), .Q ( new_AGEMA_signal_19539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C ( clk ), .D ( new_AGEMA_signal_19542 ), .Q ( new_AGEMA_signal_19543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C ( clk ), .D ( new_AGEMA_signal_19546 ), .Q ( new_AGEMA_signal_19547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C ( clk ), .D ( new_AGEMA_signal_19550 ), .Q ( new_AGEMA_signal_19551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C ( clk ), .D ( new_AGEMA_signal_19554 ), .Q ( new_AGEMA_signal_19555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C ( clk ), .D ( new_AGEMA_signal_19558 ), .Q ( new_AGEMA_signal_19559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C ( clk ), .D ( new_AGEMA_signal_19602 ), .Q ( new_AGEMA_signal_19603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C ( clk ), .D ( new_AGEMA_signal_19606 ), .Q ( new_AGEMA_signal_19607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C ( clk ), .D ( new_AGEMA_signal_19610 ), .Q ( new_AGEMA_signal_19611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C ( clk ), .D ( new_AGEMA_signal_19614 ), .Q ( new_AGEMA_signal_19615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C ( clk ), .D ( new_AGEMA_signal_19618 ), .Q ( new_AGEMA_signal_19619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C ( clk ), .D ( new_AGEMA_signal_19622 ), .Q ( new_AGEMA_signal_19623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C ( clk ), .D ( new_AGEMA_signal_19626 ), .Q ( new_AGEMA_signal_19627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C ( clk ), .D ( new_AGEMA_signal_19630 ), .Q ( new_AGEMA_signal_19631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C ( clk ), .D ( new_AGEMA_signal_19634 ), .Q ( new_AGEMA_signal_19635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C ( clk ), .D ( new_AGEMA_signal_19638 ), .Q ( new_AGEMA_signal_19639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C ( clk ), .D ( new_AGEMA_signal_19642 ), .Q ( new_AGEMA_signal_19643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C ( clk ), .D ( new_AGEMA_signal_19646 ), .Q ( new_AGEMA_signal_19647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C ( clk ), .D ( new_AGEMA_signal_19650 ), .Q ( new_AGEMA_signal_19651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C ( clk ), .D ( new_AGEMA_signal_19654 ), .Q ( new_AGEMA_signal_19655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C ( clk ), .D ( new_AGEMA_signal_19658 ), .Q ( new_AGEMA_signal_19659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C ( clk ), .D ( new_AGEMA_signal_19692 ), .Q ( new_AGEMA_signal_19693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C ( clk ), .D ( new_AGEMA_signal_19696 ), .Q ( new_AGEMA_signal_19697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C ( clk ), .D ( new_AGEMA_signal_19700 ), .Q ( new_AGEMA_signal_19701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C ( clk ), .D ( new_AGEMA_signal_19704 ), .Q ( new_AGEMA_signal_19705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C ( clk ), .D ( new_AGEMA_signal_19708 ), .Q ( new_AGEMA_signal_19709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C ( clk ), .D ( new_AGEMA_signal_19722 ), .Q ( new_AGEMA_signal_19723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C ( clk ), .D ( new_AGEMA_signal_19726 ), .Q ( new_AGEMA_signal_19727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C ( clk ), .D ( new_AGEMA_signal_19730 ), .Q ( new_AGEMA_signal_19731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C ( clk ), .D ( new_AGEMA_signal_19734 ), .Q ( new_AGEMA_signal_19735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C ( clk ), .D ( new_AGEMA_signal_19738 ), .Q ( new_AGEMA_signal_19739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C ( clk ), .D ( new_AGEMA_signal_19744 ), .Q ( new_AGEMA_signal_19745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C ( clk ), .D ( new_AGEMA_signal_19750 ), .Q ( new_AGEMA_signal_19751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C ( clk ), .D ( new_AGEMA_signal_19756 ), .Q ( new_AGEMA_signal_19757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C ( clk ), .D ( new_AGEMA_signal_19762 ), .Q ( new_AGEMA_signal_19763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C ( clk ), .D ( new_AGEMA_signal_19768 ), .Q ( new_AGEMA_signal_19769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C ( clk ), .D ( new_AGEMA_signal_19772 ), .Q ( new_AGEMA_signal_19773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C ( clk ), .D ( new_AGEMA_signal_19776 ), .Q ( new_AGEMA_signal_19777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C ( clk ), .D ( new_AGEMA_signal_19780 ), .Q ( new_AGEMA_signal_19781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C ( clk ), .D ( new_AGEMA_signal_19784 ), .Q ( new_AGEMA_signal_19785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C ( clk ), .D ( new_AGEMA_signal_19788 ), .Q ( new_AGEMA_signal_19789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C ( clk ), .D ( new_AGEMA_signal_19792 ), .Q ( new_AGEMA_signal_19793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C ( clk ), .D ( new_AGEMA_signal_19796 ), .Q ( new_AGEMA_signal_19797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C ( clk ), .D ( new_AGEMA_signal_19800 ), .Q ( new_AGEMA_signal_19801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C ( clk ), .D ( new_AGEMA_signal_19804 ), .Q ( new_AGEMA_signal_19805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C ( clk ), .D ( new_AGEMA_signal_19808 ), .Q ( new_AGEMA_signal_19809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C ( clk ), .D ( new_AGEMA_signal_19852 ), .Q ( new_AGEMA_signal_19853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C ( clk ), .D ( new_AGEMA_signal_19856 ), .Q ( new_AGEMA_signal_19857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C ( clk ), .D ( new_AGEMA_signal_19860 ), .Q ( new_AGEMA_signal_19861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C ( clk ), .D ( new_AGEMA_signal_19864 ), .Q ( new_AGEMA_signal_19865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C ( clk ), .D ( new_AGEMA_signal_19868 ), .Q ( new_AGEMA_signal_19869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C ( clk ), .D ( new_AGEMA_signal_19874 ), .Q ( new_AGEMA_signal_19875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C ( clk ), .D ( new_AGEMA_signal_19880 ), .Q ( new_AGEMA_signal_19881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C ( clk ), .D ( new_AGEMA_signal_19886 ), .Q ( new_AGEMA_signal_19887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C ( clk ), .D ( new_AGEMA_signal_19892 ), .Q ( new_AGEMA_signal_19893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C ( clk ), .D ( new_AGEMA_signal_19898 ), .Q ( new_AGEMA_signal_19899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C ( clk ), .D ( new_AGEMA_signal_19902 ), .Q ( new_AGEMA_signal_19903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C ( clk ), .D ( new_AGEMA_signal_19906 ), .Q ( new_AGEMA_signal_19907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C ( clk ), .D ( new_AGEMA_signal_19910 ), .Q ( new_AGEMA_signal_19911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C ( clk ), .D ( new_AGEMA_signal_19914 ), .Q ( new_AGEMA_signal_19915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C ( clk ), .D ( new_AGEMA_signal_19918 ), .Q ( new_AGEMA_signal_19919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C ( clk ), .D ( new_AGEMA_signal_19952 ), .Q ( new_AGEMA_signal_19953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C ( clk ), .D ( new_AGEMA_signal_19956 ), .Q ( new_AGEMA_signal_19957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C ( clk ), .D ( new_AGEMA_signal_19960 ), .Q ( new_AGEMA_signal_19961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C ( clk ), .D ( new_AGEMA_signal_19964 ), .Q ( new_AGEMA_signal_19965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C ( clk ), .D ( new_AGEMA_signal_19968 ), .Q ( new_AGEMA_signal_19969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C ( clk ), .D ( new_AGEMA_signal_19992 ), .Q ( new_AGEMA_signal_19993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C ( clk ), .D ( new_AGEMA_signal_19996 ), .Q ( new_AGEMA_signal_19997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C ( clk ), .D ( new_AGEMA_signal_20000 ), .Q ( new_AGEMA_signal_20001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C ( clk ), .D ( new_AGEMA_signal_20004 ), .Q ( new_AGEMA_signal_20005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C ( clk ), .D ( new_AGEMA_signal_20008 ), .Q ( new_AGEMA_signal_20009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C ( clk ), .D ( new_AGEMA_signal_20012 ), .Q ( new_AGEMA_signal_20013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C ( clk ), .D ( new_AGEMA_signal_20016 ), .Q ( new_AGEMA_signal_20017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C ( clk ), .D ( new_AGEMA_signal_20020 ), .Q ( new_AGEMA_signal_20021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C ( clk ), .D ( new_AGEMA_signal_20024 ), .Q ( new_AGEMA_signal_20025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C ( clk ), .D ( new_AGEMA_signal_20028 ), .Q ( new_AGEMA_signal_20029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C ( clk ), .D ( new_AGEMA_signal_20032 ), .Q ( new_AGEMA_signal_20033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C ( clk ), .D ( new_AGEMA_signal_20036 ), .Q ( new_AGEMA_signal_20037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C ( clk ), .D ( new_AGEMA_signal_20040 ), .Q ( new_AGEMA_signal_20041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C ( clk ), .D ( new_AGEMA_signal_20044 ), .Q ( new_AGEMA_signal_20045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C ( clk ), .D ( new_AGEMA_signal_20048 ), .Q ( new_AGEMA_signal_20049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C ( clk ), .D ( new_AGEMA_signal_20052 ), .Q ( new_AGEMA_signal_20053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C ( clk ), .D ( new_AGEMA_signal_20056 ), .Q ( new_AGEMA_signal_20057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C ( clk ), .D ( new_AGEMA_signal_20060 ), .Q ( new_AGEMA_signal_20061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C ( clk ), .D ( new_AGEMA_signal_20064 ), .Q ( new_AGEMA_signal_20065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C ( clk ), .D ( new_AGEMA_signal_20068 ), .Q ( new_AGEMA_signal_20069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C ( clk ), .D ( new_AGEMA_signal_20072 ), .Q ( new_AGEMA_signal_20073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C ( clk ), .D ( new_AGEMA_signal_20076 ), .Q ( new_AGEMA_signal_20077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C ( clk ), .D ( new_AGEMA_signal_20080 ), .Q ( new_AGEMA_signal_20081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C ( clk ), .D ( new_AGEMA_signal_20084 ), .Q ( new_AGEMA_signal_20085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C ( clk ), .D ( new_AGEMA_signal_20088 ), .Q ( new_AGEMA_signal_20089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C ( clk ), .D ( new_AGEMA_signal_20132 ), .Q ( new_AGEMA_signal_20133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C ( clk ), .D ( new_AGEMA_signal_20136 ), .Q ( new_AGEMA_signal_20137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C ( clk ), .D ( new_AGEMA_signal_20140 ), .Q ( new_AGEMA_signal_20141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C ( clk ), .D ( new_AGEMA_signal_20144 ), .Q ( new_AGEMA_signal_20145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C ( clk ), .D ( new_AGEMA_signal_20148 ), .Q ( new_AGEMA_signal_20149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C ( clk ), .D ( new_AGEMA_signal_20152 ), .Q ( new_AGEMA_signal_20153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C ( clk ), .D ( new_AGEMA_signal_20156 ), .Q ( new_AGEMA_signal_20157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C ( clk ), .D ( new_AGEMA_signal_20160 ), .Q ( new_AGEMA_signal_20161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C ( clk ), .D ( new_AGEMA_signal_20164 ), .Q ( new_AGEMA_signal_20165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C ( clk ), .D ( new_AGEMA_signal_20168 ), .Q ( new_AGEMA_signal_20169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C ( clk ), .D ( new_AGEMA_signal_20262 ), .Q ( new_AGEMA_signal_20263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C ( clk ), .D ( new_AGEMA_signal_20266 ), .Q ( new_AGEMA_signal_20267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C ( clk ), .D ( new_AGEMA_signal_20270 ), .Q ( new_AGEMA_signal_20271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C ( clk ), .D ( new_AGEMA_signal_20274 ), .Q ( new_AGEMA_signal_20275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C ( clk ), .D ( new_AGEMA_signal_20278 ), .Q ( new_AGEMA_signal_20279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C ( clk ), .D ( new_AGEMA_signal_20332 ), .Q ( new_AGEMA_signal_20333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C ( clk ), .D ( new_AGEMA_signal_20336 ), .Q ( new_AGEMA_signal_20337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C ( clk ), .D ( new_AGEMA_signal_20340 ), .Q ( new_AGEMA_signal_20341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C ( clk ), .D ( new_AGEMA_signal_20344 ), .Q ( new_AGEMA_signal_20345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C ( clk ), .D ( new_AGEMA_signal_20348 ), .Q ( new_AGEMA_signal_20349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C ( clk ), .D ( new_AGEMA_signal_20352 ), .Q ( new_AGEMA_signal_20353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C ( clk ), .D ( new_AGEMA_signal_20356 ), .Q ( new_AGEMA_signal_20357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C ( clk ), .D ( new_AGEMA_signal_20360 ), .Q ( new_AGEMA_signal_20361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C ( clk ), .D ( new_AGEMA_signal_20364 ), .Q ( new_AGEMA_signal_20365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C ( clk ), .D ( new_AGEMA_signal_20368 ), .Q ( new_AGEMA_signal_20369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C ( clk ), .D ( new_AGEMA_signal_20372 ), .Q ( new_AGEMA_signal_20373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C ( clk ), .D ( new_AGEMA_signal_20376 ), .Q ( new_AGEMA_signal_20377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C ( clk ), .D ( new_AGEMA_signal_20380 ), .Q ( new_AGEMA_signal_20381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C ( clk ), .D ( new_AGEMA_signal_20384 ), .Q ( new_AGEMA_signal_20385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C ( clk ), .D ( new_AGEMA_signal_20388 ), .Q ( new_AGEMA_signal_20389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C ( clk ), .D ( new_AGEMA_signal_20392 ), .Q ( new_AGEMA_signal_20393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C ( clk ), .D ( new_AGEMA_signal_20396 ), .Q ( new_AGEMA_signal_20397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C ( clk ), .D ( new_AGEMA_signal_20400 ), .Q ( new_AGEMA_signal_20401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C ( clk ), .D ( new_AGEMA_signal_20404 ), .Q ( new_AGEMA_signal_20405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C ( clk ), .D ( new_AGEMA_signal_20408 ), .Q ( new_AGEMA_signal_20409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C ( clk ), .D ( new_AGEMA_signal_20454 ), .Q ( new_AGEMA_signal_20455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C ( clk ), .D ( new_AGEMA_signal_20462 ), .Q ( new_AGEMA_signal_20463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C ( clk ), .D ( new_AGEMA_signal_20470 ), .Q ( new_AGEMA_signal_20471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C ( clk ), .D ( new_AGEMA_signal_20478 ), .Q ( new_AGEMA_signal_20479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C ( clk ), .D ( new_AGEMA_signal_20486 ), .Q ( new_AGEMA_signal_20487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C ( clk ), .D ( new_AGEMA_signal_20504 ), .Q ( new_AGEMA_signal_20505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C ( clk ), .D ( new_AGEMA_signal_20512 ), .Q ( new_AGEMA_signal_20513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C ( clk ), .D ( new_AGEMA_signal_20520 ), .Q ( new_AGEMA_signal_20521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C ( clk ), .D ( new_AGEMA_signal_20528 ), .Q ( new_AGEMA_signal_20529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C ( clk ), .D ( new_AGEMA_signal_20536 ), .Q ( new_AGEMA_signal_20537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C ( clk ), .D ( new_AGEMA_signal_20542 ), .Q ( new_AGEMA_signal_20543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C ( clk ), .D ( new_AGEMA_signal_20548 ), .Q ( new_AGEMA_signal_20549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C ( clk ), .D ( new_AGEMA_signal_20554 ), .Q ( new_AGEMA_signal_20555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C ( clk ), .D ( new_AGEMA_signal_20560 ), .Q ( new_AGEMA_signal_20561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C ( clk ), .D ( new_AGEMA_signal_20566 ), .Q ( new_AGEMA_signal_20567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C ( clk ), .D ( new_AGEMA_signal_20592 ), .Q ( new_AGEMA_signal_20593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C ( clk ), .D ( new_AGEMA_signal_20598 ), .Q ( new_AGEMA_signal_20599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C ( clk ), .D ( new_AGEMA_signal_20604 ), .Q ( new_AGEMA_signal_20605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C ( clk ), .D ( new_AGEMA_signal_20610 ), .Q ( new_AGEMA_signal_20611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C ( clk ), .D ( new_AGEMA_signal_20616 ), .Q ( new_AGEMA_signal_20617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C ( clk ), .D ( new_AGEMA_signal_20632 ), .Q ( new_AGEMA_signal_20633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C ( clk ), .D ( new_AGEMA_signal_20638 ), .Q ( new_AGEMA_signal_20639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C ( clk ), .D ( new_AGEMA_signal_20644 ), .Q ( new_AGEMA_signal_20645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C ( clk ), .D ( new_AGEMA_signal_20650 ), .Q ( new_AGEMA_signal_20651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C ( clk ), .D ( new_AGEMA_signal_20656 ), .Q ( new_AGEMA_signal_20657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C ( clk ), .D ( new_AGEMA_signal_20662 ), .Q ( new_AGEMA_signal_20663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C ( clk ), .D ( new_AGEMA_signal_20668 ), .Q ( new_AGEMA_signal_20669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C ( clk ), .D ( new_AGEMA_signal_20674 ), .Q ( new_AGEMA_signal_20675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C ( clk ), .D ( new_AGEMA_signal_20680 ), .Q ( new_AGEMA_signal_20681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C ( clk ), .D ( new_AGEMA_signal_20686 ), .Q ( new_AGEMA_signal_20687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C ( clk ), .D ( new_AGEMA_signal_20722 ), .Q ( new_AGEMA_signal_20723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C ( clk ), .D ( new_AGEMA_signal_20728 ), .Q ( new_AGEMA_signal_20729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C ( clk ), .D ( new_AGEMA_signal_20734 ), .Q ( new_AGEMA_signal_20735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C ( clk ), .D ( new_AGEMA_signal_20740 ), .Q ( new_AGEMA_signal_20741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C ( clk ), .D ( new_AGEMA_signal_20746 ), .Q ( new_AGEMA_signal_20747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C ( clk ), .D ( new_AGEMA_signal_20752 ), .Q ( new_AGEMA_signal_20753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C ( clk ), .D ( new_AGEMA_signal_20758 ), .Q ( new_AGEMA_signal_20759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C ( clk ), .D ( new_AGEMA_signal_20764 ), .Q ( new_AGEMA_signal_20765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C ( clk ), .D ( new_AGEMA_signal_20770 ), .Q ( new_AGEMA_signal_20771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C ( clk ), .D ( new_AGEMA_signal_20776 ), .Q ( new_AGEMA_signal_20777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C ( clk ), .D ( new_AGEMA_signal_20792 ), .Q ( new_AGEMA_signal_20793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C ( clk ), .D ( new_AGEMA_signal_20798 ), .Q ( new_AGEMA_signal_20799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C ( clk ), .D ( new_AGEMA_signal_20804 ), .Q ( new_AGEMA_signal_20805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C ( clk ), .D ( new_AGEMA_signal_20810 ), .Q ( new_AGEMA_signal_20811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C ( clk ), .D ( new_AGEMA_signal_20816 ), .Q ( new_AGEMA_signal_20817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C ( clk ), .D ( new_AGEMA_signal_20884 ), .Q ( new_AGEMA_signal_20885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C ( clk ), .D ( new_AGEMA_signal_20892 ), .Q ( new_AGEMA_signal_20893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C ( clk ), .D ( new_AGEMA_signal_20900 ), .Q ( new_AGEMA_signal_20901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C ( clk ), .D ( new_AGEMA_signal_20908 ), .Q ( new_AGEMA_signal_20909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C ( clk ), .D ( new_AGEMA_signal_20916 ), .Q ( new_AGEMA_signal_20917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C ( clk ), .D ( new_AGEMA_signal_20922 ), .Q ( new_AGEMA_signal_20923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C ( clk ), .D ( new_AGEMA_signal_20928 ), .Q ( new_AGEMA_signal_20929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C ( clk ), .D ( new_AGEMA_signal_20934 ), .Q ( new_AGEMA_signal_20935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C ( clk ), .D ( new_AGEMA_signal_20940 ), .Q ( new_AGEMA_signal_20941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C ( clk ), .D ( new_AGEMA_signal_20946 ), .Q ( new_AGEMA_signal_20947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C ( clk ), .D ( new_AGEMA_signal_21062 ), .Q ( new_AGEMA_signal_21063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C ( clk ), .D ( new_AGEMA_signal_21068 ), .Q ( new_AGEMA_signal_21069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C ( clk ), .D ( new_AGEMA_signal_21074 ), .Q ( new_AGEMA_signal_21075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C ( clk ), .D ( new_AGEMA_signal_21080 ), .Q ( new_AGEMA_signal_21081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C ( clk ), .D ( new_AGEMA_signal_21086 ), .Q ( new_AGEMA_signal_21087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C ( clk ), .D ( new_AGEMA_signal_21222 ), .Q ( new_AGEMA_signal_21223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C ( clk ), .D ( new_AGEMA_signal_21228 ), .Q ( new_AGEMA_signal_21229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C ( clk ), .D ( new_AGEMA_signal_21234 ), .Q ( new_AGEMA_signal_21235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C ( clk ), .D ( new_AGEMA_signal_21240 ), .Q ( new_AGEMA_signal_21241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C ( clk ), .D ( new_AGEMA_signal_21246 ), .Q ( new_AGEMA_signal_21247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C ( clk ), .D ( new_AGEMA_signal_21252 ), .Q ( new_AGEMA_signal_21253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C ( clk ), .D ( new_AGEMA_signal_21258 ), .Q ( new_AGEMA_signal_21259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C ( clk ), .D ( new_AGEMA_signal_21264 ), .Q ( new_AGEMA_signal_21265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C ( clk ), .D ( new_AGEMA_signal_21270 ), .Q ( new_AGEMA_signal_21271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C ( clk ), .D ( new_AGEMA_signal_21276 ), .Q ( new_AGEMA_signal_21277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C ( clk ), .D ( new_AGEMA_signal_21314 ), .Q ( new_AGEMA_signal_21315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C ( clk ), .D ( new_AGEMA_signal_21322 ), .Q ( new_AGEMA_signal_21323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C ( clk ), .D ( new_AGEMA_signal_21330 ), .Q ( new_AGEMA_signal_21331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C ( clk ), .D ( new_AGEMA_signal_21338 ), .Q ( new_AGEMA_signal_21339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C ( clk ), .D ( new_AGEMA_signal_21346 ), .Q ( new_AGEMA_signal_21347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C ( clk ), .D ( new_AGEMA_signal_21464 ), .Q ( new_AGEMA_signal_21465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C ( clk ), .D ( new_AGEMA_signal_21472 ), .Q ( new_AGEMA_signal_21473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C ( clk ), .D ( new_AGEMA_signal_21480 ), .Q ( new_AGEMA_signal_21481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C ( clk ), .D ( new_AGEMA_signal_21488 ), .Q ( new_AGEMA_signal_21489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C ( clk ), .D ( new_AGEMA_signal_21496 ), .Q ( new_AGEMA_signal_21497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C ( clk ), .D ( new_AGEMA_signal_21542 ), .Q ( new_AGEMA_signal_21543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C ( clk ), .D ( new_AGEMA_signal_21548 ), .Q ( new_AGEMA_signal_21549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C ( clk ), .D ( new_AGEMA_signal_21554 ), .Q ( new_AGEMA_signal_21555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C ( clk ), .D ( new_AGEMA_signal_21560 ), .Q ( new_AGEMA_signal_21561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C ( clk ), .D ( new_AGEMA_signal_21566 ), .Q ( new_AGEMA_signal_21567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C ( clk ), .D ( new_AGEMA_signal_21582 ), .Q ( new_AGEMA_signal_21583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C ( clk ), .D ( new_AGEMA_signal_21590 ), .Q ( new_AGEMA_signal_21591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C ( clk ), .D ( new_AGEMA_signal_21598 ), .Q ( new_AGEMA_signal_21599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C ( clk ), .D ( new_AGEMA_signal_21606 ), .Q ( new_AGEMA_signal_21607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C ( clk ), .D ( new_AGEMA_signal_21614 ), .Q ( new_AGEMA_signal_21615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C ( clk ), .D ( new_AGEMA_signal_21652 ), .Q ( new_AGEMA_signal_21653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C ( clk ), .D ( new_AGEMA_signal_21660 ), .Q ( new_AGEMA_signal_21661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C ( clk ), .D ( new_AGEMA_signal_21668 ), .Q ( new_AGEMA_signal_21669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C ( clk ), .D ( new_AGEMA_signal_21676 ), .Q ( new_AGEMA_signal_21677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C ( clk ), .D ( new_AGEMA_signal_21684 ), .Q ( new_AGEMA_signal_21685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C ( clk ), .D ( new_AGEMA_signal_21752 ), .Q ( new_AGEMA_signal_21753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C ( clk ), .D ( new_AGEMA_signal_21760 ), .Q ( new_AGEMA_signal_21761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C ( clk ), .D ( new_AGEMA_signal_21768 ), .Q ( new_AGEMA_signal_21769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C ( clk ), .D ( new_AGEMA_signal_21776 ), .Q ( new_AGEMA_signal_21777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C ( clk ), .D ( new_AGEMA_signal_21784 ), .Q ( new_AGEMA_signal_21785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C ( clk ), .D ( new_AGEMA_signal_21982 ), .Q ( new_AGEMA_signal_21983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C ( clk ), .D ( new_AGEMA_signal_21990 ), .Q ( new_AGEMA_signal_21991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C ( clk ), .D ( new_AGEMA_signal_21998 ), .Q ( new_AGEMA_signal_21999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C ( clk ), .D ( new_AGEMA_signal_22006 ), .Q ( new_AGEMA_signal_22007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C ( clk ), .D ( new_AGEMA_signal_22014 ), .Q ( new_AGEMA_signal_22015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C ( clk ), .D ( new_AGEMA_signal_22072 ), .Q ( new_AGEMA_signal_22073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C ( clk ), .D ( new_AGEMA_signal_22080 ), .Q ( new_AGEMA_signal_22081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C ( clk ), .D ( new_AGEMA_signal_22088 ), .Q ( new_AGEMA_signal_22089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C ( clk ), .D ( new_AGEMA_signal_22096 ), .Q ( new_AGEMA_signal_22097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C ( clk ), .D ( new_AGEMA_signal_22104 ), .Q ( new_AGEMA_signal_22105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C ( clk ), .D ( new_AGEMA_signal_22232 ), .Q ( new_AGEMA_signal_22233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C ( clk ), .D ( new_AGEMA_signal_22240 ), .Q ( new_AGEMA_signal_22241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C ( clk ), .D ( new_AGEMA_signal_22248 ), .Q ( new_AGEMA_signal_22249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C ( clk ), .D ( new_AGEMA_signal_22256 ), .Q ( new_AGEMA_signal_22257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C ( clk ), .D ( new_AGEMA_signal_22264 ), .Q ( new_AGEMA_signal_22265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C ( clk ), .D ( new_AGEMA_signal_22272 ), .Q ( new_AGEMA_signal_22273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C ( clk ), .D ( new_AGEMA_signal_22280 ), .Q ( new_AGEMA_signal_22281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C ( clk ), .D ( new_AGEMA_signal_22288 ), .Q ( new_AGEMA_signal_22289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C ( clk ), .D ( new_AGEMA_signal_22296 ), .Q ( new_AGEMA_signal_22297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C ( clk ), .D ( new_AGEMA_signal_22304 ), .Q ( new_AGEMA_signal_22305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C ( clk ), .D ( new_AGEMA_signal_22702 ), .Q ( new_AGEMA_signal_22703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C ( clk ), .D ( new_AGEMA_signal_22712 ), .Q ( new_AGEMA_signal_22713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C ( clk ), .D ( new_AGEMA_signal_22722 ), .Q ( new_AGEMA_signal_22723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C ( clk ), .D ( new_AGEMA_signal_22732 ), .Q ( new_AGEMA_signal_22733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C ( clk ), .D ( new_AGEMA_signal_22742 ), .Q ( new_AGEMA_signal_22743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C ( clk ), .D ( new_AGEMA_signal_22952 ), .Q ( new_AGEMA_signal_22953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C ( clk ), .D ( new_AGEMA_signal_22962 ), .Q ( new_AGEMA_signal_22963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C ( clk ), .D ( new_AGEMA_signal_22972 ), .Q ( new_AGEMA_signal_22973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C ( clk ), .D ( new_AGEMA_signal_22982 ), .Q ( new_AGEMA_signal_22983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C ( clk ), .D ( new_AGEMA_signal_22992 ), .Q ( new_AGEMA_signal_22993 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_2629 ( .C ( clk ), .D ( new_AGEMA_signal_19403 ), .Q ( new_AGEMA_signal_19404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C ( clk ), .D ( new_AGEMA_signal_19407 ), .Q ( new_AGEMA_signal_19408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C ( clk ), .D ( new_AGEMA_signal_19411 ), .Q ( new_AGEMA_signal_19412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C ( clk ), .D ( new_AGEMA_signal_19415 ), .Q ( new_AGEMA_signal_19416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C ( clk ), .D ( new_AGEMA_signal_19419 ), .Q ( new_AGEMA_signal_19420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C ( clk ), .D ( new_AGEMA_signal_19423 ), .Q ( new_AGEMA_signal_19424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C ( clk ), .D ( new_AGEMA_signal_19427 ), .Q ( new_AGEMA_signal_19428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C ( clk ), .D ( new_AGEMA_signal_19431 ), .Q ( new_AGEMA_signal_19432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C ( clk ), .D ( new_AGEMA_signal_19435 ), .Q ( new_AGEMA_signal_19436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C ( clk ), .D ( new_AGEMA_signal_19439 ), .Q ( new_AGEMA_signal_19440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C ( clk ), .D ( new_AGEMA_signal_19213 ), .Q ( new_AGEMA_signal_19442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C ( clk ), .D ( new_AGEMA_signal_19215 ), .Q ( new_AGEMA_signal_19444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C ( clk ), .D ( new_AGEMA_signal_19217 ), .Q ( new_AGEMA_signal_19446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C ( clk ), .D ( new_AGEMA_signal_19219 ), .Q ( new_AGEMA_signal_19448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C ( clk ), .D ( new_AGEMA_signal_19221 ), .Q ( new_AGEMA_signal_19450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_19452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C ( clk ), .D ( new_AGEMA_signal_2458 ), .Q ( new_AGEMA_signal_19454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C ( clk ), .D ( new_AGEMA_signal_2459 ), .Q ( new_AGEMA_signal_19456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C ( clk ), .D ( new_AGEMA_signal_2460 ), .Q ( new_AGEMA_signal_19458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C ( clk ), .D ( new_AGEMA_signal_2461 ), .Q ( new_AGEMA_signal_19460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C ( clk ), .D ( new_AGEMA_signal_19463 ), .Q ( new_AGEMA_signal_19464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C ( clk ), .D ( new_AGEMA_signal_19467 ), .Q ( new_AGEMA_signal_19468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C ( clk ), .D ( new_AGEMA_signal_19471 ), .Q ( new_AGEMA_signal_19472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C ( clk ), .D ( new_AGEMA_signal_19475 ), .Q ( new_AGEMA_signal_19476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C ( clk ), .D ( new_AGEMA_signal_19479 ), .Q ( new_AGEMA_signal_19480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C ( clk ), .D ( new_AGEMA_signal_19033 ), .Q ( new_AGEMA_signal_19482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C ( clk ), .D ( new_AGEMA_signal_19035 ), .Q ( new_AGEMA_signal_19484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C ( clk ), .D ( new_AGEMA_signal_19037 ), .Q ( new_AGEMA_signal_19486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C ( clk ), .D ( new_AGEMA_signal_19039 ), .Q ( new_AGEMA_signal_19488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C ( clk ), .D ( new_AGEMA_signal_19041 ), .Q ( new_AGEMA_signal_19490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C ( clk ), .D ( new_AGEMA_signal_19493 ), .Q ( new_AGEMA_signal_19494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C ( clk ), .D ( new_AGEMA_signal_19497 ), .Q ( new_AGEMA_signal_19498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C ( clk ), .D ( new_AGEMA_signal_19501 ), .Q ( new_AGEMA_signal_19502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C ( clk ), .D ( new_AGEMA_signal_19505 ), .Q ( new_AGEMA_signal_19506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C ( clk ), .D ( new_AGEMA_signal_19509 ), .Q ( new_AGEMA_signal_19510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_19512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C ( clk ), .D ( new_AGEMA_signal_2498 ), .Q ( new_AGEMA_signal_19514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C ( clk ), .D ( new_AGEMA_signal_2499 ), .Q ( new_AGEMA_signal_19516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C ( clk ), .D ( new_AGEMA_signal_2500 ), .Q ( new_AGEMA_signal_19518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C ( clk ), .D ( new_AGEMA_signal_2501 ), .Q ( new_AGEMA_signal_19520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C ( clk ), .D ( new_AGEMA_signal_19523 ), .Q ( new_AGEMA_signal_19524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C ( clk ), .D ( new_AGEMA_signal_19527 ), .Q ( new_AGEMA_signal_19528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C ( clk ), .D ( new_AGEMA_signal_19531 ), .Q ( new_AGEMA_signal_19532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C ( clk ), .D ( new_AGEMA_signal_19535 ), .Q ( new_AGEMA_signal_19536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C ( clk ), .D ( new_AGEMA_signal_19539 ), .Q ( new_AGEMA_signal_19540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C ( clk ), .D ( new_AGEMA_signal_19543 ), .Q ( new_AGEMA_signal_19544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C ( clk ), .D ( new_AGEMA_signal_19547 ), .Q ( new_AGEMA_signal_19548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C ( clk ), .D ( new_AGEMA_signal_19551 ), .Q ( new_AGEMA_signal_19552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C ( clk ), .D ( new_AGEMA_signal_19555 ), .Q ( new_AGEMA_signal_19556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C ( clk ), .D ( new_AGEMA_signal_19559 ), .Q ( new_AGEMA_signal_19560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_19562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C ( clk ), .D ( new_AGEMA_signal_2522 ), .Q ( new_AGEMA_signal_19564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C ( clk ), .D ( new_AGEMA_signal_2523 ), .Q ( new_AGEMA_signal_19566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C ( clk ), .D ( new_AGEMA_signal_2524 ), .Q ( new_AGEMA_signal_19568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C ( clk ), .D ( new_AGEMA_signal_2525 ), .Q ( new_AGEMA_signal_19570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C ( clk ), .D ( new_AGEMA_signal_18813 ), .Q ( new_AGEMA_signal_19572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C ( clk ), .D ( new_AGEMA_signal_18815 ), .Q ( new_AGEMA_signal_19574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C ( clk ), .D ( new_AGEMA_signal_18817 ), .Q ( new_AGEMA_signal_19576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C ( clk ), .D ( new_AGEMA_signal_18819 ), .Q ( new_AGEMA_signal_19578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C ( clk ), .D ( new_AGEMA_signal_18821 ), .Q ( new_AGEMA_signal_19580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C ( clk ), .D ( new_AGEMA_signal_18863 ), .Q ( new_AGEMA_signal_19582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C ( clk ), .D ( new_AGEMA_signal_18865 ), .Q ( new_AGEMA_signal_19584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C ( clk ), .D ( new_AGEMA_signal_18867 ), .Q ( new_AGEMA_signal_19586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C ( clk ), .D ( new_AGEMA_signal_18869 ), .Q ( new_AGEMA_signal_19588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C ( clk ), .D ( new_AGEMA_signal_18871 ), .Q ( new_AGEMA_signal_19590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C ( clk ), .D ( new_AGEMA_signal_19003 ), .Q ( new_AGEMA_signal_19592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C ( clk ), .D ( new_AGEMA_signal_19005 ), .Q ( new_AGEMA_signal_19594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C ( clk ), .D ( new_AGEMA_signal_19007 ), .Q ( new_AGEMA_signal_19596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C ( clk ), .D ( new_AGEMA_signal_19009 ), .Q ( new_AGEMA_signal_19598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C ( clk ), .D ( new_AGEMA_signal_19011 ), .Q ( new_AGEMA_signal_19600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C ( clk ), .D ( new_AGEMA_signal_19603 ), .Q ( new_AGEMA_signal_19604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C ( clk ), .D ( new_AGEMA_signal_19607 ), .Q ( new_AGEMA_signal_19608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C ( clk ), .D ( new_AGEMA_signal_19611 ), .Q ( new_AGEMA_signal_19612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C ( clk ), .D ( new_AGEMA_signal_19615 ), .Q ( new_AGEMA_signal_19616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C ( clk ), .D ( new_AGEMA_signal_19619 ), .Q ( new_AGEMA_signal_19620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C ( clk ), .D ( new_AGEMA_signal_19623 ), .Q ( new_AGEMA_signal_19624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C ( clk ), .D ( new_AGEMA_signal_19627 ), .Q ( new_AGEMA_signal_19628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C ( clk ), .D ( new_AGEMA_signal_19631 ), .Q ( new_AGEMA_signal_19632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C ( clk ), .D ( new_AGEMA_signal_19635 ), .Q ( new_AGEMA_signal_19636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C ( clk ), .D ( new_AGEMA_signal_19639 ), .Q ( new_AGEMA_signal_19640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C ( clk ), .D ( new_AGEMA_signal_19643 ), .Q ( new_AGEMA_signal_19644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C ( clk ), .D ( new_AGEMA_signal_19647 ), .Q ( new_AGEMA_signal_19648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C ( clk ), .D ( new_AGEMA_signal_19651 ), .Q ( new_AGEMA_signal_19652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C ( clk ), .D ( new_AGEMA_signal_19655 ), .Q ( new_AGEMA_signal_19656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C ( clk ), .D ( new_AGEMA_signal_19659 ), .Q ( new_AGEMA_signal_19660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_19662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C ( clk ), .D ( new_AGEMA_signal_2582 ), .Q ( new_AGEMA_signal_19664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C ( clk ), .D ( new_AGEMA_signal_2583 ), .Q ( new_AGEMA_signal_19666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C ( clk ), .D ( new_AGEMA_signal_2584 ), .Q ( new_AGEMA_signal_19668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C ( clk ), .D ( new_AGEMA_signal_2585 ), .Q ( new_AGEMA_signal_19670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_19672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C ( clk ), .D ( new_AGEMA_signal_2590 ), .Q ( new_AGEMA_signal_19674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C ( clk ), .D ( new_AGEMA_signal_2591 ), .Q ( new_AGEMA_signal_19676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C ( clk ), .D ( new_AGEMA_signal_2592 ), .Q ( new_AGEMA_signal_19678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C ( clk ), .D ( new_AGEMA_signal_2593 ), .Q ( new_AGEMA_signal_19680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_19682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C ( clk ), .D ( new_AGEMA_signal_1934 ), .Q ( new_AGEMA_signal_19684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C ( clk ), .D ( new_AGEMA_signal_1935 ), .Q ( new_AGEMA_signal_19686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C ( clk ), .D ( new_AGEMA_signal_1936 ), .Q ( new_AGEMA_signal_19688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C ( clk ), .D ( new_AGEMA_signal_1937 ), .Q ( new_AGEMA_signal_19690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C ( clk ), .D ( new_AGEMA_signal_19693 ), .Q ( new_AGEMA_signal_19694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C ( clk ), .D ( new_AGEMA_signal_19697 ), .Q ( new_AGEMA_signal_19698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C ( clk ), .D ( new_AGEMA_signal_19701 ), .Q ( new_AGEMA_signal_19702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C ( clk ), .D ( new_AGEMA_signal_19705 ), .Q ( new_AGEMA_signal_19706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C ( clk ), .D ( new_AGEMA_signal_19709 ), .Q ( new_AGEMA_signal_19710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_19712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C ( clk ), .D ( new_AGEMA_signal_2454 ), .Q ( new_AGEMA_signal_19714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C ( clk ), .D ( new_AGEMA_signal_2455 ), .Q ( new_AGEMA_signal_19716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C ( clk ), .D ( new_AGEMA_signal_2456 ), .Q ( new_AGEMA_signal_19718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C ( clk ), .D ( new_AGEMA_signal_2457 ), .Q ( new_AGEMA_signal_19720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C ( clk ), .D ( new_AGEMA_signal_19723 ), .Q ( new_AGEMA_signal_19724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C ( clk ), .D ( new_AGEMA_signal_19727 ), .Q ( new_AGEMA_signal_19728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C ( clk ), .D ( new_AGEMA_signal_19731 ), .Q ( new_AGEMA_signal_19732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C ( clk ), .D ( new_AGEMA_signal_19735 ), .Q ( new_AGEMA_signal_19736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C ( clk ), .D ( new_AGEMA_signal_19739 ), .Q ( new_AGEMA_signal_19740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C ( clk ), .D ( new_AGEMA_signal_19745 ), .Q ( new_AGEMA_signal_19746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C ( clk ), .D ( new_AGEMA_signal_19751 ), .Q ( new_AGEMA_signal_19752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C ( clk ), .D ( new_AGEMA_signal_19757 ), .Q ( new_AGEMA_signal_19758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C ( clk ), .D ( new_AGEMA_signal_19763 ), .Q ( new_AGEMA_signal_19764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C ( clk ), .D ( new_AGEMA_signal_19769 ), .Q ( new_AGEMA_signal_19770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C ( clk ), .D ( new_AGEMA_signal_19773 ), .Q ( new_AGEMA_signal_19774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C ( clk ), .D ( new_AGEMA_signal_19777 ), .Q ( new_AGEMA_signal_19778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C ( clk ), .D ( new_AGEMA_signal_19781 ), .Q ( new_AGEMA_signal_19782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C ( clk ), .D ( new_AGEMA_signal_19785 ), .Q ( new_AGEMA_signal_19786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C ( clk ), .D ( new_AGEMA_signal_19789 ), .Q ( new_AGEMA_signal_19790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C ( clk ), .D ( new_AGEMA_signal_19793 ), .Q ( new_AGEMA_signal_19794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C ( clk ), .D ( new_AGEMA_signal_19797 ), .Q ( new_AGEMA_signal_19798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C ( clk ), .D ( new_AGEMA_signal_19801 ), .Q ( new_AGEMA_signal_19802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C ( clk ), .D ( new_AGEMA_signal_19805 ), .Q ( new_AGEMA_signal_19806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C ( clk ), .D ( new_AGEMA_signal_19809 ), .Q ( new_AGEMA_signal_19810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_19812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C ( clk ), .D ( new_AGEMA_signal_2662 ), .Q ( new_AGEMA_signal_19814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C ( clk ), .D ( new_AGEMA_signal_2663 ), .Q ( new_AGEMA_signal_19816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C ( clk ), .D ( new_AGEMA_signal_2664 ), .Q ( new_AGEMA_signal_19818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C ( clk ), .D ( new_AGEMA_signal_2665 ), .Q ( new_AGEMA_signal_19820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_19822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C ( clk ), .D ( new_AGEMA_signal_3238 ), .Q ( new_AGEMA_signal_19824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C ( clk ), .D ( new_AGEMA_signal_3239 ), .Q ( new_AGEMA_signal_19826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C ( clk ), .D ( new_AGEMA_signal_3240 ), .Q ( new_AGEMA_signal_19828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C ( clk ), .D ( new_AGEMA_signal_3241 ), .Q ( new_AGEMA_signal_19830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_19832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C ( clk ), .D ( new_AGEMA_signal_2030 ), .Q ( new_AGEMA_signal_19834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C ( clk ), .D ( new_AGEMA_signal_2031 ), .Q ( new_AGEMA_signal_19836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C ( clk ), .D ( new_AGEMA_signal_2032 ), .Q ( new_AGEMA_signal_19838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C ( clk ), .D ( new_AGEMA_signal_2033 ), .Q ( new_AGEMA_signal_19840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_19842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C ( clk ), .D ( new_AGEMA_signal_2434 ), .Q ( new_AGEMA_signal_19844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C ( clk ), .D ( new_AGEMA_signal_2435 ), .Q ( new_AGEMA_signal_19846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C ( clk ), .D ( new_AGEMA_signal_2436 ), .Q ( new_AGEMA_signal_19848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C ( clk ), .D ( new_AGEMA_signal_2437 ), .Q ( new_AGEMA_signal_19850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C ( clk ), .D ( new_AGEMA_signal_19853 ), .Q ( new_AGEMA_signal_19854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C ( clk ), .D ( new_AGEMA_signal_19857 ), .Q ( new_AGEMA_signal_19858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C ( clk ), .D ( new_AGEMA_signal_19861 ), .Q ( new_AGEMA_signal_19862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C ( clk ), .D ( new_AGEMA_signal_19865 ), .Q ( new_AGEMA_signal_19866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C ( clk ), .D ( new_AGEMA_signal_19869 ), .Q ( new_AGEMA_signal_19870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C ( clk ), .D ( new_AGEMA_signal_19875 ), .Q ( new_AGEMA_signal_19876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C ( clk ), .D ( new_AGEMA_signal_19881 ), .Q ( new_AGEMA_signal_19882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C ( clk ), .D ( new_AGEMA_signal_19887 ), .Q ( new_AGEMA_signal_19888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C ( clk ), .D ( new_AGEMA_signal_19893 ), .Q ( new_AGEMA_signal_19894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C ( clk ), .D ( new_AGEMA_signal_19899 ), .Q ( new_AGEMA_signal_19900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C ( clk ), .D ( new_AGEMA_signal_19903 ), .Q ( new_AGEMA_signal_19904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C ( clk ), .D ( new_AGEMA_signal_19907 ), .Q ( new_AGEMA_signal_19908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C ( clk ), .D ( new_AGEMA_signal_19911 ), .Q ( new_AGEMA_signal_19912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C ( clk ), .D ( new_AGEMA_signal_19915 ), .Q ( new_AGEMA_signal_19916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C ( clk ), .D ( new_AGEMA_signal_19919 ), .Q ( new_AGEMA_signal_19920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_19922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C ( clk ), .D ( new_AGEMA_signal_3274 ), .Q ( new_AGEMA_signal_19924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C ( clk ), .D ( new_AGEMA_signal_3275 ), .Q ( new_AGEMA_signal_19926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C ( clk ), .D ( new_AGEMA_signal_3276 ), .Q ( new_AGEMA_signal_19928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C ( clk ), .D ( new_AGEMA_signal_3277 ), .Q ( new_AGEMA_signal_19930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C ( clk ), .D ( new_AGEMA_signal_19137 ), .Q ( new_AGEMA_signal_19932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C ( clk ), .D ( new_AGEMA_signal_19143 ), .Q ( new_AGEMA_signal_19934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C ( clk ), .D ( new_AGEMA_signal_19149 ), .Q ( new_AGEMA_signal_19936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C ( clk ), .D ( new_AGEMA_signal_19155 ), .Q ( new_AGEMA_signal_19938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C ( clk ), .D ( new_AGEMA_signal_19161 ), .Q ( new_AGEMA_signal_19940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_19942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C ( clk ), .D ( new_AGEMA_signal_2746 ), .Q ( new_AGEMA_signal_19944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C ( clk ), .D ( new_AGEMA_signal_2747 ), .Q ( new_AGEMA_signal_19946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C ( clk ), .D ( new_AGEMA_signal_2748 ), .Q ( new_AGEMA_signal_19948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C ( clk ), .D ( new_AGEMA_signal_2749 ), .Q ( new_AGEMA_signal_19950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C ( clk ), .D ( new_AGEMA_signal_19953 ), .Q ( new_AGEMA_signal_19954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C ( clk ), .D ( new_AGEMA_signal_19957 ), .Q ( new_AGEMA_signal_19958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C ( clk ), .D ( new_AGEMA_signal_19961 ), .Q ( new_AGEMA_signal_19962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C ( clk ), .D ( new_AGEMA_signal_19965 ), .Q ( new_AGEMA_signal_19966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C ( clk ), .D ( new_AGEMA_signal_19969 ), .Q ( new_AGEMA_signal_19970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_19972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C ( clk ), .D ( new_AGEMA_signal_2782 ), .Q ( new_AGEMA_signal_19974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C ( clk ), .D ( new_AGEMA_signal_2783 ), .Q ( new_AGEMA_signal_19976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C ( clk ), .D ( new_AGEMA_signal_2784 ), .Q ( new_AGEMA_signal_19978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C ( clk ), .D ( new_AGEMA_signal_2785 ), .Q ( new_AGEMA_signal_19980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_19982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C ( clk ), .D ( new_AGEMA_signal_2802 ), .Q ( new_AGEMA_signal_19984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C ( clk ), .D ( new_AGEMA_signal_2803 ), .Q ( new_AGEMA_signal_19986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C ( clk ), .D ( new_AGEMA_signal_2804 ), .Q ( new_AGEMA_signal_19988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C ( clk ), .D ( new_AGEMA_signal_2805 ), .Q ( new_AGEMA_signal_19990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C ( clk ), .D ( new_AGEMA_signal_19993 ), .Q ( new_AGEMA_signal_19994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C ( clk ), .D ( new_AGEMA_signal_19997 ), .Q ( new_AGEMA_signal_19998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C ( clk ), .D ( new_AGEMA_signal_20001 ), .Q ( new_AGEMA_signal_20002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C ( clk ), .D ( new_AGEMA_signal_20005 ), .Q ( new_AGEMA_signal_20006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C ( clk ), .D ( new_AGEMA_signal_20009 ), .Q ( new_AGEMA_signal_20010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C ( clk ), .D ( new_AGEMA_signal_20013 ), .Q ( new_AGEMA_signal_20014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C ( clk ), .D ( new_AGEMA_signal_20017 ), .Q ( new_AGEMA_signal_20018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C ( clk ), .D ( new_AGEMA_signal_20021 ), .Q ( new_AGEMA_signal_20022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C ( clk ), .D ( new_AGEMA_signal_20025 ), .Q ( new_AGEMA_signal_20026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C ( clk ), .D ( new_AGEMA_signal_20029 ), .Q ( new_AGEMA_signal_20030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C ( clk ), .D ( new_AGEMA_signal_20033 ), .Q ( new_AGEMA_signal_20034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C ( clk ), .D ( new_AGEMA_signal_20037 ), .Q ( new_AGEMA_signal_20038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C ( clk ), .D ( new_AGEMA_signal_20041 ), .Q ( new_AGEMA_signal_20042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C ( clk ), .D ( new_AGEMA_signal_20045 ), .Q ( new_AGEMA_signal_20046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C ( clk ), .D ( new_AGEMA_signal_20049 ), .Q ( new_AGEMA_signal_20050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C ( clk ), .D ( new_AGEMA_signal_20053 ), .Q ( new_AGEMA_signal_20054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C ( clk ), .D ( new_AGEMA_signal_20057 ), .Q ( new_AGEMA_signal_20058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C ( clk ), .D ( new_AGEMA_signal_20061 ), .Q ( new_AGEMA_signal_20062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C ( clk ), .D ( new_AGEMA_signal_20065 ), .Q ( new_AGEMA_signal_20066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C ( clk ), .D ( new_AGEMA_signal_20069 ), .Q ( new_AGEMA_signal_20070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C ( clk ), .D ( new_AGEMA_signal_20073 ), .Q ( new_AGEMA_signal_20074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C ( clk ), .D ( new_AGEMA_signal_20077 ), .Q ( new_AGEMA_signal_20078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C ( clk ), .D ( new_AGEMA_signal_20081 ), .Q ( new_AGEMA_signal_20082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C ( clk ), .D ( new_AGEMA_signal_20085 ), .Q ( new_AGEMA_signal_20086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C ( clk ), .D ( new_AGEMA_signal_20089 ), .Q ( new_AGEMA_signal_20090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_20092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C ( clk ), .D ( new_AGEMA_signal_2830 ), .Q ( new_AGEMA_signal_20094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C ( clk ), .D ( new_AGEMA_signal_2831 ), .Q ( new_AGEMA_signal_20096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C ( clk ), .D ( new_AGEMA_signal_2832 ), .Q ( new_AGEMA_signal_20098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C ( clk ), .D ( new_AGEMA_signal_2833 ), .Q ( new_AGEMA_signal_20100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C ( clk ), .D ( new_AGEMA_signal_18845 ), .Q ( new_AGEMA_signal_20102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C ( clk ), .D ( new_AGEMA_signal_18849 ), .Q ( new_AGEMA_signal_20104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C ( clk ), .D ( new_AGEMA_signal_18853 ), .Q ( new_AGEMA_signal_20106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C ( clk ), .D ( new_AGEMA_signal_18857 ), .Q ( new_AGEMA_signal_20108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C ( clk ), .D ( new_AGEMA_signal_18861 ), .Q ( new_AGEMA_signal_20110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_20112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C ( clk ), .D ( new_AGEMA_signal_2734 ), .Q ( new_AGEMA_signal_20114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C ( clk ), .D ( new_AGEMA_signal_2735 ), .Q ( new_AGEMA_signal_20116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C ( clk ), .D ( new_AGEMA_signal_2736 ), .Q ( new_AGEMA_signal_20118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C ( clk ), .D ( new_AGEMA_signal_2737 ), .Q ( new_AGEMA_signal_20120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_20122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C ( clk ), .D ( new_AGEMA_signal_2158 ), .Q ( new_AGEMA_signal_20124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C ( clk ), .D ( new_AGEMA_signal_2159 ), .Q ( new_AGEMA_signal_20126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C ( clk ), .D ( new_AGEMA_signal_2160 ), .Q ( new_AGEMA_signal_20128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C ( clk ), .D ( new_AGEMA_signal_2161 ), .Q ( new_AGEMA_signal_20130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C ( clk ), .D ( new_AGEMA_signal_20133 ), .Q ( new_AGEMA_signal_20134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C ( clk ), .D ( new_AGEMA_signal_20137 ), .Q ( new_AGEMA_signal_20138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C ( clk ), .D ( new_AGEMA_signal_20141 ), .Q ( new_AGEMA_signal_20142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C ( clk ), .D ( new_AGEMA_signal_20145 ), .Q ( new_AGEMA_signal_20146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C ( clk ), .D ( new_AGEMA_signal_20149 ), .Q ( new_AGEMA_signal_20150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C ( clk ), .D ( new_AGEMA_signal_20153 ), .Q ( new_AGEMA_signal_20154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C ( clk ), .D ( new_AGEMA_signal_20157 ), .Q ( new_AGEMA_signal_20158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C ( clk ), .D ( new_AGEMA_signal_20161 ), .Q ( new_AGEMA_signal_20162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C ( clk ), .D ( new_AGEMA_signal_20165 ), .Q ( new_AGEMA_signal_20166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C ( clk ), .D ( new_AGEMA_signal_20169 ), .Q ( new_AGEMA_signal_20170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_20172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C ( clk ), .D ( new_AGEMA_signal_2238 ), .Q ( new_AGEMA_signal_20174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C ( clk ), .D ( new_AGEMA_signal_2239 ), .Q ( new_AGEMA_signal_20176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C ( clk ), .D ( new_AGEMA_signal_2240 ), .Q ( new_AGEMA_signal_20178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C ( clk ), .D ( new_AGEMA_signal_2241 ), .Q ( new_AGEMA_signal_20180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_20182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C ( clk ), .D ( new_AGEMA_signal_2242 ), .Q ( new_AGEMA_signal_20184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C ( clk ), .D ( new_AGEMA_signal_2243 ), .Q ( new_AGEMA_signal_20186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C ( clk ), .D ( new_AGEMA_signal_2244 ), .Q ( new_AGEMA_signal_20188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C ( clk ), .D ( new_AGEMA_signal_2245 ), .Q ( new_AGEMA_signal_20190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_20192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C ( clk ), .D ( new_AGEMA_signal_2882 ), .Q ( new_AGEMA_signal_20194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C ( clk ), .D ( new_AGEMA_signal_2883 ), .Q ( new_AGEMA_signal_20196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C ( clk ), .D ( new_AGEMA_signal_2884 ), .Q ( new_AGEMA_signal_20198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C ( clk ), .D ( new_AGEMA_signal_2885 ), .Q ( new_AGEMA_signal_20200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_20202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C ( clk ), .D ( new_AGEMA_signal_2906 ), .Q ( new_AGEMA_signal_20204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C ( clk ), .D ( new_AGEMA_signal_2907 ), .Q ( new_AGEMA_signal_20206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C ( clk ), .D ( new_AGEMA_signal_2908 ), .Q ( new_AGEMA_signal_20208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C ( clk ), .D ( new_AGEMA_signal_2909 ), .Q ( new_AGEMA_signal_20210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_20212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C ( clk ), .D ( new_AGEMA_signal_2918 ), .Q ( new_AGEMA_signal_20214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C ( clk ), .D ( new_AGEMA_signal_2919 ), .Q ( new_AGEMA_signal_20216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C ( clk ), .D ( new_AGEMA_signal_2920 ), .Q ( new_AGEMA_signal_20218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C ( clk ), .D ( new_AGEMA_signal_2921 ), .Q ( new_AGEMA_signal_20220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_20222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C ( clk ), .D ( new_AGEMA_signal_2926 ), .Q ( new_AGEMA_signal_20224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C ( clk ), .D ( new_AGEMA_signal_2927 ), .Q ( new_AGEMA_signal_20226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C ( clk ), .D ( new_AGEMA_signal_2928 ), .Q ( new_AGEMA_signal_20228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C ( clk ), .D ( new_AGEMA_signal_2929 ), .Q ( new_AGEMA_signal_20230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_20232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C ( clk ), .D ( new_AGEMA_signal_2278 ), .Q ( new_AGEMA_signal_20234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C ( clk ), .D ( new_AGEMA_signal_2279 ), .Q ( new_AGEMA_signal_20236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C ( clk ), .D ( new_AGEMA_signal_2280 ), .Q ( new_AGEMA_signal_20238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C ( clk ), .D ( new_AGEMA_signal_2281 ), .Q ( new_AGEMA_signal_20240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_20242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C ( clk ), .D ( new_AGEMA_signal_2958 ), .Q ( new_AGEMA_signal_20244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C ( clk ), .D ( new_AGEMA_signal_2959 ), .Q ( new_AGEMA_signal_20246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C ( clk ), .D ( new_AGEMA_signal_2960 ), .Q ( new_AGEMA_signal_20248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C ( clk ), .D ( new_AGEMA_signal_2961 ), .Q ( new_AGEMA_signal_20250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_20252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C ( clk ), .D ( new_AGEMA_signal_2962 ), .Q ( new_AGEMA_signal_20254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C ( clk ), .D ( new_AGEMA_signal_2963 ), .Q ( new_AGEMA_signal_20256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C ( clk ), .D ( new_AGEMA_signal_2964 ), .Q ( new_AGEMA_signal_20258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C ( clk ), .D ( new_AGEMA_signal_2965 ), .Q ( new_AGEMA_signal_20260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C ( clk ), .D ( new_AGEMA_signal_20263 ), .Q ( new_AGEMA_signal_20264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C ( clk ), .D ( new_AGEMA_signal_20267 ), .Q ( new_AGEMA_signal_20268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C ( clk ), .D ( new_AGEMA_signal_20271 ), .Q ( new_AGEMA_signal_20272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C ( clk ), .D ( new_AGEMA_signal_20275 ), .Q ( new_AGEMA_signal_20276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C ( clk ), .D ( new_AGEMA_signal_20279 ), .Q ( new_AGEMA_signal_20280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_20282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C ( clk ), .D ( new_AGEMA_signal_2330 ), .Q ( new_AGEMA_signal_20284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C ( clk ), .D ( new_AGEMA_signal_2331 ), .Q ( new_AGEMA_signal_20286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C ( clk ), .D ( new_AGEMA_signal_2332 ), .Q ( new_AGEMA_signal_20288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C ( clk ), .D ( new_AGEMA_signal_2333 ), .Q ( new_AGEMA_signal_20290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_20292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C ( clk ), .D ( new_AGEMA_signal_2426 ), .Q ( new_AGEMA_signal_20294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C ( clk ), .D ( new_AGEMA_signal_2427 ), .Q ( new_AGEMA_signal_20296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C ( clk ), .D ( new_AGEMA_signal_2428 ), .Q ( new_AGEMA_signal_20298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C ( clk ), .D ( new_AGEMA_signal_2429 ), .Q ( new_AGEMA_signal_20300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_20302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C ( clk ), .D ( new_AGEMA_signal_2342 ), .Q ( new_AGEMA_signal_20304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C ( clk ), .D ( new_AGEMA_signal_2343 ), .Q ( new_AGEMA_signal_20306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C ( clk ), .D ( new_AGEMA_signal_2344 ), .Q ( new_AGEMA_signal_20308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C ( clk ), .D ( new_AGEMA_signal_2345 ), .Q ( new_AGEMA_signal_20310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_20312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C ( clk ), .D ( new_AGEMA_signal_2998 ), .Q ( new_AGEMA_signal_20314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C ( clk ), .D ( new_AGEMA_signal_2999 ), .Q ( new_AGEMA_signal_20316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C ( clk ), .D ( new_AGEMA_signal_3000 ), .Q ( new_AGEMA_signal_20318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C ( clk ), .D ( new_AGEMA_signal_3001 ), .Q ( new_AGEMA_signal_20320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_20322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C ( clk ), .D ( new_AGEMA_signal_3478 ), .Q ( new_AGEMA_signal_20324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C ( clk ), .D ( new_AGEMA_signal_3479 ), .Q ( new_AGEMA_signal_20326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C ( clk ), .D ( new_AGEMA_signal_3480 ), .Q ( new_AGEMA_signal_20328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C ( clk ), .D ( new_AGEMA_signal_3481 ), .Q ( new_AGEMA_signal_20330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C ( clk ), .D ( new_AGEMA_signal_20333 ), .Q ( new_AGEMA_signal_20334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C ( clk ), .D ( new_AGEMA_signal_20337 ), .Q ( new_AGEMA_signal_20338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C ( clk ), .D ( new_AGEMA_signal_20341 ), .Q ( new_AGEMA_signal_20342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C ( clk ), .D ( new_AGEMA_signal_20345 ), .Q ( new_AGEMA_signal_20346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C ( clk ), .D ( new_AGEMA_signal_20349 ), .Q ( new_AGEMA_signal_20350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C ( clk ), .D ( new_AGEMA_signal_20353 ), .Q ( new_AGEMA_signal_20354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C ( clk ), .D ( new_AGEMA_signal_20357 ), .Q ( new_AGEMA_signal_20358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C ( clk ), .D ( new_AGEMA_signal_20361 ), .Q ( new_AGEMA_signal_20362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C ( clk ), .D ( new_AGEMA_signal_20365 ), .Q ( new_AGEMA_signal_20366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C ( clk ), .D ( new_AGEMA_signal_20369 ), .Q ( new_AGEMA_signal_20370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C ( clk ), .D ( new_AGEMA_signal_20373 ), .Q ( new_AGEMA_signal_20374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C ( clk ), .D ( new_AGEMA_signal_20377 ), .Q ( new_AGEMA_signal_20378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C ( clk ), .D ( new_AGEMA_signal_20381 ), .Q ( new_AGEMA_signal_20382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C ( clk ), .D ( new_AGEMA_signal_20385 ), .Q ( new_AGEMA_signal_20386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C ( clk ), .D ( new_AGEMA_signal_20389 ), .Q ( new_AGEMA_signal_20390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C ( clk ), .D ( new_AGEMA_signal_20393 ), .Q ( new_AGEMA_signal_20394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C ( clk ), .D ( new_AGEMA_signal_20397 ), .Q ( new_AGEMA_signal_20398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C ( clk ), .D ( new_AGEMA_signal_20401 ), .Q ( new_AGEMA_signal_20402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C ( clk ), .D ( new_AGEMA_signal_20405 ), .Q ( new_AGEMA_signal_20406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C ( clk ), .D ( new_AGEMA_signal_20409 ), .Q ( new_AGEMA_signal_20410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C ( clk ), .D ( new_AGEMA_signal_19073 ), .Q ( new_AGEMA_signal_20412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C ( clk ), .D ( new_AGEMA_signal_19075 ), .Q ( new_AGEMA_signal_20416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C ( clk ), .D ( new_AGEMA_signal_19077 ), .Q ( new_AGEMA_signal_20420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C ( clk ), .D ( new_AGEMA_signal_19079 ), .Q ( new_AGEMA_signal_20424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C ( clk ), .D ( new_AGEMA_signal_19081 ), .Q ( new_AGEMA_signal_20428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_20432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C ( clk ), .D ( new_AGEMA_signal_2442 ), .Q ( new_AGEMA_signal_20436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C ( clk ), .D ( new_AGEMA_signal_2443 ), .Q ( new_AGEMA_signal_20440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C ( clk ), .D ( new_AGEMA_signal_2444 ), .Q ( new_AGEMA_signal_20444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C ( clk ), .D ( new_AGEMA_signal_2445 ), .Q ( new_AGEMA_signal_20448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C ( clk ), .D ( new_AGEMA_signal_20455 ), .Q ( new_AGEMA_signal_20456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C ( clk ), .D ( new_AGEMA_signal_20463 ), .Q ( new_AGEMA_signal_20464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C ( clk ), .D ( new_AGEMA_signal_20471 ), .Q ( new_AGEMA_signal_20472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C ( clk ), .D ( new_AGEMA_signal_20479 ), .Q ( new_AGEMA_signal_20480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C ( clk ), .D ( new_AGEMA_signal_20487 ), .Q ( new_AGEMA_signal_20488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C ( clk ), .D ( new_AGEMA_signal_20505 ), .Q ( new_AGEMA_signal_20506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C ( clk ), .D ( new_AGEMA_signal_20513 ), .Q ( new_AGEMA_signal_20514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C ( clk ), .D ( new_AGEMA_signal_20521 ), .Q ( new_AGEMA_signal_20522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C ( clk ), .D ( new_AGEMA_signal_20529 ), .Q ( new_AGEMA_signal_20530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C ( clk ), .D ( new_AGEMA_signal_20537 ), .Q ( new_AGEMA_signal_20538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C ( clk ), .D ( new_AGEMA_signal_20543 ), .Q ( new_AGEMA_signal_20544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C ( clk ), .D ( new_AGEMA_signal_20549 ), .Q ( new_AGEMA_signal_20550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C ( clk ), .D ( new_AGEMA_signal_20555 ), .Q ( new_AGEMA_signal_20556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C ( clk ), .D ( new_AGEMA_signal_20561 ), .Q ( new_AGEMA_signal_20562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C ( clk ), .D ( new_AGEMA_signal_20567 ), .Q ( new_AGEMA_signal_20568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_20572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C ( clk ), .D ( new_AGEMA_signal_1838 ), .Q ( new_AGEMA_signal_20576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C ( clk ), .D ( new_AGEMA_signal_1839 ), .Q ( new_AGEMA_signal_20580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C ( clk ), .D ( new_AGEMA_signal_1840 ), .Q ( new_AGEMA_signal_20584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C ( clk ), .D ( new_AGEMA_signal_1841 ), .Q ( new_AGEMA_signal_20588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C ( clk ), .D ( new_AGEMA_signal_20593 ), .Q ( new_AGEMA_signal_20594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C ( clk ), .D ( new_AGEMA_signal_20599 ), .Q ( new_AGEMA_signal_20600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C ( clk ), .D ( new_AGEMA_signal_20605 ), .Q ( new_AGEMA_signal_20606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C ( clk ), .D ( new_AGEMA_signal_20611 ), .Q ( new_AGEMA_signal_20612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C ( clk ), .D ( new_AGEMA_signal_20617 ), .Q ( new_AGEMA_signal_20618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C ( clk ), .D ( new_AGEMA_signal_20633 ), .Q ( new_AGEMA_signal_20634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C ( clk ), .D ( new_AGEMA_signal_20639 ), .Q ( new_AGEMA_signal_20640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C ( clk ), .D ( new_AGEMA_signal_20645 ), .Q ( new_AGEMA_signal_20646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C ( clk ), .D ( new_AGEMA_signal_20651 ), .Q ( new_AGEMA_signal_20652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C ( clk ), .D ( new_AGEMA_signal_20657 ), .Q ( new_AGEMA_signal_20658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C ( clk ), .D ( new_AGEMA_signal_20663 ), .Q ( new_AGEMA_signal_20664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C ( clk ), .D ( new_AGEMA_signal_20669 ), .Q ( new_AGEMA_signal_20670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C ( clk ), .D ( new_AGEMA_signal_20675 ), .Q ( new_AGEMA_signal_20676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C ( clk ), .D ( new_AGEMA_signal_20681 ), .Q ( new_AGEMA_signal_20682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C ( clk ), .D ( new_AGEMA_signal_20687 ), .Q ( new_AGEMA_signal_20688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_20702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C ( clk ), .D ( new_AGEMA_signal_2594 ), .Q ( new_AGEMA_signal_20706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C ( clk ), .D ( new_AGEMA_signal_2595 ), .Q ( new_AGEMA_signal_20710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C ( clk ), .D ( new_AGEMA_signal_2596 ), .Q ( new_AGEMA_signal_20714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C ( clk ), .D ( new_AGEMA_signal_2597 ), .Q ( new_AGEMA_signal_20718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C ( clk ), .D ( new_AGEMA_signal_20723 ), .Q ( new_AGEMA_signal_20724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C ( clk ), .D ( new_AGEMA_signal_20729 ), .Q ( new_AGEMA_signal_20730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C ( clk ), .D ( new_AGEMA_signal_20735 ), .Q ( new_AGEMA_signal_20736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C ( clk ), .D ( new_AGEMA_signal_20741 ), .Q ( new_AGEMA_signal_20742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C ( clk ), .D ( new_AGEMA_signal_20747 ), .Q ( new_AGEMA_signal_20748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C ( clk ), .D ( new_AGEMA_signal_20753 ), .Q ( new_AGEMA_signal_20754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C ( clk ), .D ( new_AGEMA_signal_20759 ), .Q ( new_AGEMA_signal_20760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C ( clk ), .D ( new_AGEMA_signal_20765 ), .Q ( new_AGEMA_signal_20766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C ( clk ), .D ( new_AGEMA_signal_20771 ), .Q ( new_AGEMA_signal_20772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C ( clk ), .D ( new_AGEMA_signal_20777 ), .Q ( new_AGEMA_signal_20778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C ( clk ), .D ( new_AGEMA_signal_20793 ), .Q ( new_AGEMA_signal_20794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C ( clk ), .D ( new_AGEMA_signal_20799 ), .Q ( new_AGEMA_signal_20800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C ( clk ), .D ( new_AGEMA_signal_20805 ), .Q ( new_AGEMA_signal_20806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C ( clk ), .D ( new_AGEMA_signal_20811 ), .Q ( new_AGEMA_signal_20812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C ( clk ), .D ( new_AGEMA_signal_20817 ), .Q ( new_AGEMA_signal_20818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_20832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C ( clk ), .D ( new_AGEMA_signal_2650 ), .Q ( new_AGEMA_signal_20836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C ( clk ), .D ( new_AGEMA_signal_2651 ), .Q ( new_AGEMA_signal_20840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C ( clk ), .D ( new_AGEMA_signal_2652 ), .Q ( new_AGEMA_signal_20844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C ( clk ), .D ( new_AGEMA_signal_2653 ), .Q ( new_AGEMA_signal_20848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_20852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C ( clk ), .D ( new_AGEMA_signal_2658 ), .Q ( new_AGEMA_signal_20856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C ( clk ), .D ( new_AGEMA_signal_2659 ), .Q ( new_AGEMA_signal_20860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C ( clk ), .D ( new_AGEMA_signal_2660 ), .Q ( new_AGEMA_signal_20864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C ( clk ), .D ( new_AGEMA_signal_2661 ), .Q ( new_AGEMA_signal_20868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C ( clk ), .D ( new_AGEMA_signal_20885 ), .Q ( new_AGEMA_signal_20886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C ( clk ), .D ( new_AGEMA_signal_20893 ), .Q ( new_AGEMA_signal_20894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C ( clk ), .D ( new_AGEMA_signal_20901 ), .Q ( new_AGEMA_signal_20902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C ( clk ), .D ( new_AGEMA_signal_20909 ), .Q ( new_AGEMA_signal_20910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C ( clk ), .D ( new_AGEMA_signal_20917 ), .Q ( new_AGEMA_signal_20918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C ( clk ), .D ( new_AGEMA_signal_20923 ), .Q ( new_AGEMA_signal_20924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C ( clk ), .D ( new_AGEMA_signal_20929 ), .Q ( new_AGEMA_signal_20930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C ( clk ), .D ( new_AGEMA_signal_20935 ), .Q ( new_AGEMA_signal_20936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C ( clk ), .D ( new_AGEMA_signal_20941 ), .Q ( new_AGEMA_signal_20942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C ( clk ), .D ( new_AGEMA_signal_20947 ), .Q ( new_AGEMA_signal_20948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_20952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C ( clk ), .D ( new_AGEMA_signal_2034 ), .Q ( new_AGEMA_signal_20956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C ( clk ), .D ( new_AGEMA_signal_2035 ), .Q ( new_AGEMA_signal_20960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C ( clk ), .D ( new_AGEMA_signal_2036 ), .Q ( new_AGEMA_signal_20964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C ( clk ), .D ( new_AGEMA_signal_2037 ), .Q ( new_AGEMA_signal_20968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_20972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C ( clk ), .D ( new_AGEMA_signal_2694 ), .Q ( new_AGEMA_signal_20976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C ( clk ), .D ( new_AGEMA_signal_2695 ), .Q ( new_AGEMA_signal_20980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C ( clk ), .D ( new_AGEMA_signal_2696 ), .Q ( new_AGEMA_signal_20984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C ( clk ), .D ( new_AGEMA_signal_2697 ), .Q ( new_AGEMA_signal_20988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_21012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C ( clk ), .D ( new_AGEMA_signal_2094 ), .Q ( new_AGEMA_signal_21016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C ( clk ), .D ( new_AGEMA_signal_2095 ), .Q ( new_AGEMA_signal_21020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C ( clk ), .D ( new_AGEMA_signal_2096 ), .Q ( new_AGEMA_signal_21024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C ( clk ), .D ( new_AGEMA_signal_2097 ), .Q ( new_AGEMA_signal_21028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_21032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C ( clk ), .D ( new_AGEMA_signal_2754 ), .Q ( new_AGEMA_signal_21036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C ( clk ), .D ( new_AGEMA_signal_2755 ), .Q ( new_AGEMA_signal_21040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C ( clk ), .D ( new_AGEMA_signal_2756 ), .Q ( new_AGEMA_signal_21044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C ( clk ), .D ( new_AGEMA_signal_2757 ), .Q ( new_AGEMA_signal_21048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C ( clk ), .D ( new_AGEMA_signal_21063 ), .Q ( new_AGEMA_signal_21064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C ( clk ), .D ( new_AGEMA_signal_21069 ), .Q ( new_AGEMA_signal_21070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C ( clk ), .D ( new_AGEMA_signal_21075 ), .Q ( new_AGEMA_signal_21076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C ( clk ), .D ( new_AGEMA_signal_21081 ), .Q ( new_AGEMA_signal_21082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C ( clk ), .D ( new_AGEMA_signal_21087 ), .Q ( new_AGEMA_signal_21088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_21092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C ( clk ), .D ( new_AGEMA_signal_2786 ), .Q ( new_AGEMA_signal_21096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C ( clk ), .D ( new_AGEMA_signal_2787 ), .Q ( new_AGEMA_signal_21100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C ( clk ), .D ( new_AGEMA_signal_2788 ), .Q ( new_AGEMA_signal_21104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C ( clk ), .D ( new_AGEMA_signal_2789 ), .Q ( new_AGEMA_signal_21108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_21122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C ( clk ), .D ( new_AGEMA_signal_2170 ), .Q ( new_AGEMA_signal_21126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C ( clk ), .D ( new_AGEMA_signal_2171 ), .Q ( new_AGEMA_signal_21130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C ( clk ), .D ( new_AGEMA_signal_2172 ), .Q ( new_AGEMA_signal_21134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C ( clk ), .D ( new_AGEMA_signal_2173 ), .Q ( new_AGEMA_signal_21138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_21142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C ( clk ), .D ( new_AGEMA_signal_2810 ), .Q ( new_AGEMA_signal_21146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C ( clk ), .D ( new_AGEMA_signal_2811 ), .Q ( new_AGEMA_signal_21150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C ( clk ), .D ( new_AGEMA_signal_2812 ), .Q ( new_AGEMA_signal_21154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C ( clk ), .D ( new_AGEMA_signal_2813 ), .Q ( new_AGEMA_signal_21158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C ( clk ), .D ( new_AGEMA_signal_18573 ), .Q ( new_AGEMA_signal_21162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C ( clk ), .D ( new_AGEMA_signal_18575 ), .Q ( new_AGEMA_signal_21166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C ( clk ), .D ( new_AGEMA_signal_18577 ), .Q ( new_AGEMA_signal_21170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C ( clk ), .D ( new_AGEMA_signal_18579 ), .Q ( new_AGEMA_signal_21174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C ( clk ), .D ( new_AGEMA_signal_18581 ), .Q ( new_AGEMA_signal_21178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C ( clk ), .D ( new_AGEMA_signal_18583 ), .Q ( new_AGEMA_signal_21192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C ( clk ), .D ( new_AGEMA_signal_18585 ), .Q ( new_AGEMA_signal_21196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C ( clk ), .D ( new_AGEMA_signal_18587 ), .Q ( new_AGEMA_signal_21200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C ( clk ), .D ( new_AGEMA_signal_18589 ), .Q ( new_AGEMA_signal_21204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C ( clk ), .D ( new_AGEMA_signal_18591 ), .Q ( new_AGEMA_signal_21208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C ( clk ), .D ( new_AGEMA_signal_21223 ), .Q ( new_AGEMA_signal_21224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C ( clk ), .D ( new_AGEMA_signal_21229 ), .Q ( new_AGEMA_signal_21230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C ( clk ), .D ( new_AGEMA_signal_21235 ), .Q ( new_AGEMA_signal_21236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C ( clk ), .D ( new_AGEMA_signal_21241 ), .Q ( new_AGEMA_signal_21242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C ( clk ), .D ( new_AGEMA_signal_21247 ), .Q ( new_AGEMA_signal_21248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C ( clk ), .D ( new_AGEMA_signal_21253 ), .Q ( new_AGEMA_signal_21254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C ( clk ), .D ( new_AGEMA_signal_21259 ), .Q ( new_AGEMA_signal_21260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C ( clk ), .D ( new_AGEMA_signal_21265 ), .Q ( new_AGEMA_signal_21266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C ( clk ), .D ( new_AGEMA_signal_21271 ), .Q ( new_AGEMA_signal_21272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C ( clk ), .D ( new_AGEMA_signal_21277 ), .Q ( new_AGEMA_signal_21278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_21282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C ( clk ), .D ( new_AGEMA_signal_2250 ), .Q ( new_AGEMA_signal_21286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C ( clk ), .D ( new_AGEMA_signal_2251 ), .Q ( new_AGEMA_signal_21290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C ( clk ), .D ( new_AGEMA_signal_2252 ), .Q ( new_AGEMA_signal_21294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C ( clk ), .D ( new_AGEMA_signal_2253 ), .Q ( new_AGEMA_signal_21298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C ( clk ), .D ( new_AGEMA_signal_21315 ), .Q ( new_AGEMA_signal_21316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C ( clk ), .D ( new_AGEMA_signal_21323 ), .Q ( new_AGEMA_signal_21324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C ( clk ), .D ( new_AGEMA_signal_21331 ), .Q ( new_AGEMA_signal_21332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C ( clk ), .D ( new_AGEMA_signal_21339 ), .Q ( new_AGEMA_signal_21340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C ( clk ), .D ( new_AGEMA_signal_21347 ), .Q ( new_AGEMA_signal_21348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_21362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C ( clk ), .D ( new_AGEMA_signal_2946 ), .Q ( new_AGEMA_signal_21366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C ( clk ), .D ( new_AGEMA_signal_2947 ), .Q ( new_AGEMA_signal_21370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C ( clk ), .D ( new_AGEMA_signal_2948 ), .Q ( new_AGEMA_signal_21374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C ( clk ), .D ( new_AGEMA_signal_2949 ), .Q ( new_AGEMA_signal_21378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_21382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C ( clk ), .D ( new_AGEMA_signal_2954 ), .Q ( new_AGEMA_signal_21386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C ( clk ), .D ( new_AGEMA_signal_2955 ), .Q ( new_AGEMA_signal_21390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C ( clk ), .D ( new_AGEMA_signal_2956 ), .Q ( new_AGEMA_signal_21394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C ( clk ), .D ( new_AGEMA_signal_2957 ), .Q ( new_AGEMA_signal_21398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_21402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C ( clk ), .D ( new_AGEMA_signal_2318 ), .Q ( new_AGEMA_signal_21406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C ( clk ), .D ( new_AGEMA_signal_2319 ), .Q ( new_AGEMA_signal_21410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C ( clk ), .D ( new_AGEMA_signal_2320 ), .Q ( new_AGEMA_signal_21414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C ( clk ), .D ( new_AGEMA_signal_2321 ), .Q ( new_AGEMA_signal_21418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_21422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C ( clk ), .D ( new_AGEMA_signal_2982 ), .Q ( new_AGEMA_signal_21426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C ( clk ), .D ( new_AGEMA_signal_2983 ), .Q ( new_AGEMA_signal_21430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C ( clk ), .D ( new_AGEMA_signal_2984 ), .Q ( new_AGEMA_signal_21434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C ( clk ), .D ( new_AGEMA_signal_2985 ), .Q ( new_AGEMA_signal_21438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_21442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C ( clk ), .D ( new_AGEMA_signal_2994 ), .Q ( new_AGEMA_signal_21446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C ( clk ), .D ( new_AGEMA_signal_2995 ), .Q ( new_AGEMA_signal_21450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C ( clk ), .D ( new_AGEMA_signal_2996 ), .Q ( new_AGEMA_signal_21454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C ( clk ), .D ( new_AGEMA_signal_2997 ), .Q ( new_AGEMA_signal_21458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C ( clk ), .D ( new_AGEMA_signal_21465 ), .Q ( new_AGEMA_signal_21466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C ( clk ), .D ( new_AGEMA_signal_21473 ), .Q ( new_AGEMA_signal_21474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C ( clk ), .D ( new_AGEMA_signal_21481 ), .Q ( new_AGEMA_signal_21482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C ( clk ), .D ( new_AGEMA_signal_21489 ), .Q ( new_AGEMA_signal_21490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C ( clk ), .D ( new_AGEMA_signal_21497 ), .Q ( new_AGEMA_signal_21498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_21512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C ( clk ), .D ( new_AGEMA_signal_3026 ), .Q ( new_AGEMA_signal_21516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C ( clk ), .D ( new_AGEMA_signal_3027 ), .Q ( new_AGEMA_signal_21520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C ( clk ), .D ( new_AGEMA_signal_3028 ), .Q ( new_AGEMA_signal_21524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C ( clk ), .D ( new_AGEMA_signal_3029 ), .Q ( new_AGEMA_signal_21528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C ( clk ), .D ( new_AGEMA_signal_21543 ), .Q ( new_AGEMA_signal_21544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C ( clk ), .D ( new_AGEMA_signal_21549 ), .Q ( new_AGEMA_signal_21550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C ( clk ), .D ( new_AGEMA_signal_21555 ), .Q ( new_AGEMA_signal_21556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C ( clk ), .D ( new_AGEMA_signal_21561 ), .Q ( new_AGEMA_signal_21562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C ( clk ), .D ( new_AGEMA_signal_21567 ), .Q ( new_AGEMA_signal_21568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C ( clk ), .D ( new_AGEMA_signal_21583 ), .Q ( new_AGEMA_signal_21584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C ( clk ), .D ( new_AGEMA_signal_21591 ), .Q ( new_AGEMA_signal_21592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C ( clk ), .D ( new_AGEMA_signal_21599 ), .Q ( new_AGEMA_signal_21600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C ( clk ), .D ( new_AGEMA_signal_21607 ), .Q ( new_AGEMA_signal_21608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C ( clk ), .D ( new_AGEMA_signal_21615 ), .Q ( new_AGEMA_signal_21616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C ( clk ), .D ( new_AGEMA_signal_21653 ), .Q ( new_AGEMA_signal_21654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C ( clk ), .D ( new_AGEMA_signal_21661 ), .Q ( new_AGEMA_signal_21662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C ( clk ), .D ( new_AGEMA_signal_21669 ), .Q ( new_AGEMA_signal_21670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C ( clk ), .D ( new_AGEMA_signal_21677 ), .Q ( new_AGEMA_signal_21678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C ( clk ), .D ( new_AGEMA_signal_21685 ), .Q ( new_AGEMA_signal_21686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_21702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C ( clk ), .D ( new_AGEMA_signal_1858 ), .Q ( new_AGEMA_signal_21708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C ( clk ), .D ( new_AGEMA_signal_1859 ), .Q ( new_AGEMA_signal_21714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C ( clk ), .D ( new_AGEMA_signal_1860 ), .Q ( new_AGEMA_signal_21720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C ( clk ), .D ( new_AGEMA_signal_1861 ), .Q ( new_AGEMA_signal_21726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C ( clk ), .D ( new_AGEMA_signal_21753 ), .Q ( new_AGEMA_signal_21754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C ( clk ), .D ( new_AGEMA_signal_21761 ), .Q ( new_AGEMA_signal_21762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C ( clk ), .D ( new_AGEMA_signal_21769 ), .Q ( new_AGEMA_signal_21770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C ( clk ), .D ( new_AGEMA_signal_21777 ), .Q ( new_AGEMA_signal_21778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C ( clk ), .D ( new_AGEMA_signal_21785 ), .Q ( new_AGEMA_signal_21786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_21812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C ( clk ), .D ( new_AGEMA_signal_1518 ), .Q ( new_AGEMA_signal_21818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C ( clk ), .D ( new_AGEMA_signal_1519 ), .Q ( new_AGEMA_signal_21824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C ( clk ), .D ( new_AGEMA_signal_1520 ), .Q ( new_AGEMA_signal_21830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C ( clk ), .D ( new_AGEMA_signal_1521 ), .Q ( new_AGEMA_signal_21836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_21842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C ( clk ), .D ( new_AGEMA_signal_2010 ), .Q ( new_AGEMA_signal_21848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C ( clk ), .D ( new_AGEMA_signal_2011 ), .Q ( new_AGEMA_signal_21854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C ( clk ), .D ( new_AGEMA_signal_2012 ), .Q ( new_AGEMA_signal_21860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C ( clk ), .D ( new_AGEMA_signal_2013 ), .Q ( new_AGEMA_signal_21866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_21872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C ( clk ), .D ( new_AGEMA_signal_2038 ), .Q ( new_AGEMA_signal_21878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C ( clk ), .D ( new_AGEMA_signal_2039 ), .Q ( new_AGEMA_signal_21884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C ( clk ), .D ( new_AGEMA_signal_2040 ), .Q ( new_AGEMA_signal_21890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C ( clk ), .D ( new_AGEMA_signal_2041 ), .Q ( new_AGEMA_signal_21896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_21902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C ( clk ), .D ( new_AGEMA_signal_2702 ), .Q ( new_AGEMA_signal_21908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C ( clk ), .D ( new_AGEMA_signal_2703 ), .Q ( new_AGEMA_signal_21914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C ( clk ), .D ( new_AGEMA_signal_2704 ), .Q ( new_AGEMA_signal_21920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C ( clk ), .D ( new_AGEMA_signal_2705 ), .Q ( new_AGEMA_signal_21926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_21932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C ( clk ), .D ( new_AGEMA_signal_3270 ), .Q ( new_AGEMA_signal_21938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C ( clk ), .D ( new_AGEMA_signal_3271 ), .Q ( new_AGEMA_signal_21944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C ( clk ), .D ( new_AGEMA_signal_3272 ), .Q ( new_AGEMA_signal_21950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C ( clk ), .D ( new_AGEMA_signal_3273 ), .Q ( new_AGEMA_signal_21956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C ( clk ), .D ( new_AGEMA_signal_21983 ), .Q ( new_AGEMA_signal_21984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C ( clk ), .D ( new_AGEMA_signal_21991 ), .Q ( new_AGEMA_signal_21992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C ( clk ), .D ( new_AGEMA_signal_21999 ), .Q ( new_AGEMA_signal_22000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C ( clk ), .D ( new_AGEMA_signal_22007 ), .Q ( new_AGEMA_signal_22008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C ( clk ), .D ( new_AGEMA_signal_22015 ), .Q ( new_AGEMA_signal_22016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_22042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C ( clk ), .D ( new_AGEMA_signal_2134 ), .Q ( new_AGEMA_signal_22048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C ( clk ), .D ( new_AGEMA_signal_2135 ), .Q ( new_AGEMA_signal_22054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C ( clk ), .D ( new_AGEMA_signal_2136 ), .Q ( new_AGEMA_signal_22060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C ( clk ), .D ( new_AGEMA_signal_2137 ), .Q ( new_AGEMA_signal_22066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C ( clk ), .D ( new_AGEMA_signal_22073 ), .Q ( new_AGEMA_signal_22074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C ( clk ), .D ( new_AGEMA_signal_22081 ), .Q ( new_AGEMA_signal_22082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C ( clk ), .D ( new_AGEMA_signal_22089 ), .Q ( new_AGEMA_signal_22090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C ( clk ), .D ( new_AGEMA_signal_22097 ), .Q ( new_AGEMA_signal_22098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C ( clk ), .D ( new_AGEMA_signal_22105 ), .Q ( new_AGEMA_signal_22106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_22122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C ( clk ), .D ( new_AGEMA_signal_2178 ), .Q ( new_AGEMA_signal_22128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C ( clk ), .D ( new_AGEMA_signal_2179 ), .Q ( new_AGEMA_signal_22134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C ( clk ), .D ( new_AGEMA_signal_2180 ), .Q ( new_AGEMA_signal_22140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5371 ( .C ( clk ), .D ( new_AGEMA_signal_2181 ), .Q ( new_AGEMA_signal_22146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_22172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C ( clk ), .D ( new_AGEMA_signal_2842 ), .Q ( new_AGEMA_signal_22178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C ( clk ), .D ( new_AGEMA_signal_2843 ), .Q ( new_AGEMA_signal_22184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C ( clk ), .D ( new_AGEMA_signal_2844 ), .Q ( new_AGEMA_signal_22190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C ( clk ), .D ( new_AGEMA_signal_2845 ), .Q ( new_AGEMA_signal_22196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_22202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C ( clk ), .D ( new_AGEMA_signal_2218 ), .Q ( new_AGEMA_signal_22208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C ( clk ), .D ( new_AGEMA_signal_2219 ), .Q ( new_AGEMA_signal_22214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C ( clk ), .D ( new_AGEMA_signal_2220 ), .Q ( new_AGEMA_signal_22220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C ( clk ), .D ( new_AGEMA_signal_2221 ), .Q ( new_AGEMA_signal_22226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C ( clk ), .D ( new_AGEMA_signal_22233 ), .Q ( new_AGEMA_signal_22234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C ( clk ), .D ( new_AGEMA_signal_22241 ), .Q ( new_AGEMA_signal_22242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C ( clk ), .D ( new_AGEMA_signal_22249 ), .Q ( new_AGEMA_signal_22250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C ( clk ), .D ( new_AGEMA_signal_22257 ), .Q ( new_AGEMA_signal_22258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C ( clk ), .D ( new_AGEMA_signal_22265 ), .Q ( new_AGEMA_signal_22266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C ( clk ), .D ( new_AGEMA_signal_22273 ), .Q ( new_AGEMA_signal_22274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C ( clk ), .D ( new_AGEMA_signal_22281 ), .Q ( new_AGEMA_signal_22282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C ( clk ), .D ( new_AGEMA_signal_22289 ), .Q ( new_AGEMA_signal_22290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C ( clk ), .D ( new_AGEMA_signal_22297 ), .Q ( new_AGEMA_signal_22298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C ( clk ), .D ( new_AGEMA_signal_22305 ), .Q ( new_AGEMA_signal_22306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_22312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C ( clk ), .D ( new_AGEMA_signal_2938 ), .Q ( new_AGEMA_signal_22318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C ( clk ), .D ( new_AGEMA_signal_2939 ), .Q ( new_AGEMA_signal_22324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C ( clk ), .D ( new_AGEMA_signal_2940 ), .Q ( new_AGEMA_signal_22330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C ( clk ), .D ( new_AGEMA_signal_2941 ), .Q ( new_AGEMA_signal_22336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_22342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C ( clk ), .D ( new_AGEMA_signal_2290 ), .Q ( new_AGEMA_signal_22348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C ( clk ), .D ( new_AGEMA_signal_2291 ), .Q ( new_AGEMA_signal_22354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C ( clk ), .D ( new_AGEMA_signal_2292 ), .Q ( new_AGEMA_signal_22360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C ( clk ), .D ( new_AGEMA_signal_2293 ), .Q ( new_AGEMA_signal_22366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_22512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C ( clk ), .D ( new_AGEMA_signal_2514 ), .Q ( new_AGEMA_signal_22520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C ( clk ), .D ( new_AGEMA_signal_2515 ), .Q ( new_AGEMA_signal_22528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C ( clk ), .D ( new_AGEMA_signal_2516 ), .Q ( new_AGEMA_signal_22536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C ( clk ), .D ( new_AGEMA_signal_2517 ), .Q ( new_AGEMA_signal_22544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_22552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C ( clk ), .D ( new_AGEMA_signal_1458 ), .Q ( new_AGEMA_signal_22560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C ( clk ), .D ( new_AGEMA_signal_1459 ), .Q ( new_AGEMA_signal_22568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C ( clk ), .D ( new_AGEMA_signal_1460 ), .Q ( new_AGEMA_signal_22576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C ( clk ), .D ( new_AGEMA_signal_1461 ), .Q ( new_AGEMA_signal_22584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_22592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C ( clk ), .D ( new_AGEMA_signal_2538 ), .Q ( new_AGEMA_signal_22600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C ( clk ), .D ( new_AGEMA_signal_2539 ), .Q ( new_AGEMA_signal_22608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C ( clk ), .D ( new_AGEMA_signal_2540 ), .Q ( new_AGEMA_signal_22616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C ( clk ), .D ( new_AGEMA_signal_2541 ), .Q ( new_AGEMA_signal_22624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_22632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C ( clk ), .D ( new_AGEMA_signal_2558 ), .Q ( new_AGEMA_signal_22640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C ( clk ), .D ( new_AGEMA_signal_2559 ), .Q ( new_AGEMA_signal_22648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C ( clk ), .D ( new_AGEMA_signal_2560 ), .Q ( new_AGEMA_signal_22656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C ( clk ), .D ( new_AGEMA_signal_2561 ), .Q ( new_AGEMA_signal_22664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C ( clk ), .D ( new_AGEMA_signal_22703 ), .Q ( new_AGEMA_signal_22704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C ( clk ), .D ( new_AGEMA_signal_22713 ), .Q ( new_AGEMA_signal_22714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C ( clk ), .D ( new_AGEMA_signal_22723 ), .Q ( new_AGEMA_signal_22724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C ( clk ), .D ( new_AGEMA_signal_22733 ), .Q ( new_AGEMA_signal_22734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C ( clk ), .D ( new_AGEMA_signal_22743 ), .Q ( new_AGEMA_signal_22744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_22752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C ( clk ), .D ( new_AGEMA_signal_2626 ), .Q ( new_AGEMA_signal_22760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C ( clk ), .D ( new_AGEMA_signal_2627 ), .Q ( new_AGEMA_signal_22768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C ( clk ), .D ( new_AGEMA_signal_2628 ), .Q ( new_AGEMA_signal_22776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C ( clk ), .D ( new_AGEMA_signal_2629 ), .Q ( new_AGEMA_signal_22784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_22792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C ( clk ), .D ( new_AGEMA_signal_2634 ), .Q ( new_AGEMA_signal_22800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C ( clk ), .D ( new_AGEMA_signal_2635 ), .Q ( new_AGEMA_signal_22808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C ( clk ), .D ( new_AGEMA_signal_2636 ), .Q ( new_AGEMA_signal_22816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C ( clk ), .D ( new_AGEMA_signal_2637 ), .Q ( new_AGEMA_signal_22824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_22832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C ( clk ), .D ( new_AGEMA_signal_1510 ), .Q ( new_AGEMA_signal_22840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C ( clk ), .D ( new_AGEMA_signal_1511 ), .Q ( new_AGEMA_signal_22848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C ( clk ), .D ( new_AGEMA_signal_1512 ), .Q ( new_AGEMA_signal_22856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C ( clk ), .D ( new_AGEMA_signal_1513 ), .Q ( new_AGEMA_signal_22864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C ( clk ), .D ( new_AGEMA_signal_22953 ), .Q ( new_AGEMA_signal_22954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C ( clk ), .D ( new_AGEMA_signal_22963 ), .Q ( new_AGEMA_signal_22964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C ( clk ), .D ( new_AGEMA_signal_22973 ), .Q ( new_AGEMA_signal_22974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C ( clk ), .D ( new_AGEMA_signal_22983 ), .Q ( new_AGEMA_signal_22984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C ( clk ), .D ( new_AGEMA_signal_22993 ), .Q ( new_AGEMA_signal_22994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C ( clk ), .D ( new_AGEMA_signal_19223 ), .Q ( new_AGEMA_signal_23002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C ( clk ), .D ( new_AGEMA_signal_19225 ), .Q ( new_AGEMA_signal_23010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C ( clk ), .D ( new_AGEMA_signal_19227 ), .Q ( new_AGEMA_signal_23018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C ( clk ), .D ( new_AGEMA_signal_19229 ), .Q ( new_AGEMA_signal_23026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C ( clk ), .D ( new_AGEMA_signal_19231 ), .Q ( new_AGEMA_signal_23034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_23072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C ( clk ), .D ( new_AGEMA_signal_2914 ), .Q ( new_AGEMA_signal_23080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C ( clk ), .D ( new_AGEMA_signal_2915 ), .Q ( new_AGEMA_signal_23088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C ( clk ), .D ( new_AGEMA_signal_2916 ), .Q ( new_AGEMA_signal_23096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C ( clk ), .D ( new_AGEMA_signal_2917 ), .Q ( new_AGEMA_signal_23104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_23112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C ( clk ), .D ( new_AGEMA_signal_2950 ), .Q ( new_AGEMA_signal_23120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C ( clk ), .D ( new_AGEMA_signal_2951 ), .Q ( new_AGEMA_signal_23128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C ( clk ), .D ( new_AGEMA_signal_2952 ), .Q ( new_AGEMA_signal_23136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C ( clk ), .D ( new_AGEMA_signal_2953 ), .Q ( new_AGEMA_signal_23144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_23202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C ( clk ), .D ( new_AGEMA_signal_2346 ), .Q ( new_AGEMA_signal_23210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C ( clk ), .D ( new_AGEMA_signal_2347 ), .Q ( new_AGEMA_signal_23218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C ( clk ), .D ( new_AGEMA_signal_2348 ), .Q ( new_AGEMA_signal_23226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C ( clk ), .D ( new_AGEMA_signal_2349 ), .Q ( new_AGEMA_signal_23234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_23532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C ( clk ), .D ( new_AGEMA_signal_2646 ), .Q ( new_AGEMA_signal_23542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C ( clk ), .D ( new_AGEMA_signal_2647 ), .Q ( new_AGEMA_signal_23552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C ( clk ), .D ( new_AGEMA_signal_2648 ), .Q ( new_AGEMA_signal_23562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C ( clk ), .D ( new_AGEMA_signal_2649 ), .Q ( new_AGEMA_signal_23572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7737 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_24512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7751 ( .C ( clk ), .D ( new_AGEMA_signal_1962 ), .Q ( new_AGEMA_signal_24526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7765 ( .C ( clk ), .D ( new_AGEMA_signal_1963 ), .Q ( new_AGEMA_signal_24540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7779 ( .C ( clk ), .D ( new_AGEMA_signal_1964 ), .Q ( new_AGEMA_signal_24554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7793 ( .C ( clk ), .D ( new_AGEMA_signal_1965 ), .Q ( new_AGEMA_signal_24568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7847 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_24622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7861 ( .C ( clk ), .D ( new_AGEMA_signal_3334 ), .Q ( new_AGEMA_signal_24636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7875 ( .C ( clk ), .D ( new_AGEMA_signal_3335 ), .Q ( new_AGEMA_signal_24650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7889 ( .C ( clk ), .D ( new_AGEMA_signal_3336 ), .Q ( new_AGEMA_signal_24664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7903 ( .C ( clk ), .D ( new_AGEMA_signal_3337 ), .Q ( new_AGEMA_signal_24678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8027 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_24802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8043 ( .C ( clk ), .D ( new_AGEMA_signal_2630 ), .Q ( new_AGEMA_signal_24818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8059 ( .C ( clk ), .D ( new_AGEMA_signal_2631 ), .Q ( new_AGEMA_signal_24834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8075 ( .C ( clk ), .D ( new_AGEMA_signal_2632 ), .Q ( new_AGEMA_signal_24850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8091 ( .C ( clk ), .D ( new_AGEMA_signal_2633 ), .Q ( new_AGEMA_signal_24866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8137 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_24912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8153 ( .C ( clk ), .D ( new_AGEMA_signal_2790 ), .Q ( new_AGEMA_signal_24928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8169 ( .C ( clk ), .D ( new_AGEMA_signal_2791 ), .Q ( new_AGEMA_signal_24944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8185 ( .C ( clk ), .D ( new_AGEMA_signal_2792 ), .Q ( new_AGEMA_signal_24960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8201 ( .C ( clk ), .D ( new_AGEMA_signal_2793 ), .Q ( new_AGEMA_signal_24976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8517 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_25292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8535 ( .C ( clk ), .D ( new_AGEMA_signal_2138 ), .Q ( new_AGEMA_signal_25310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8553 ( .C ( clk ), .D ( new_AGEMA_signal_2139 ), .Q ( new_AGEMA_signal_25328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8571 ( .C ( clk ), .D ( new_AGEMA_signal_2140 ), .Q ( new_AGEMA_signal_25346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8589 ( .C ( clk ), .D ( new_AGEMA_signal_2141 ), .Q ( new_AGEMA_signal_25364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8767 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_25542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8787 ( .C ( clk ), .D ( new_AGEMA_signal_2794 ), .Q ( new_AGEMA_signal_25562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8807 ( .C ( clk ), .D ( new_AGEMA_signal_2795 ), .Q ( new_AGEMA_signal_25582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8827 ( .C ( clk ), .D ( new_AGEMA_signal_2796 ), .Q ( new_AGEMA_signal_25602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8847 ( .C ( clk ), .D ( new_AGEMA_signal_2797 ), .Q ( new_AGEMA_signal_25622 ) ) ;

    /* cells in depth 8 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1968 ( .ina ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, n1924}), .inb ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, n1923}), .clk ( clk ), .rnd ({Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770], Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765]}), .outt ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n1936}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1982 ( .ina ({new_AGEMA_signal_18541, new_AGEMA_signal_18539, new_AGEMA_signal_18537, new_AGEMA_signal_18535, new_AGEMA_signal_18533}), .inb ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n1927}), .clk ( clk ), .rnd ({Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790], Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780]}), .outt ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, n1928}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U1994 ( .ina ({new_AGEMA_signal_18551, new_AGEMA_signal_18549, new_AGEMA_signal_18547, new_AGEMA_signal_18545, new_AGEMA_signal_18543}), .inb ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, n1929}), .clk ( clk ), .rnd ({Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800], Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795]}), .outt ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, n1931}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2012 ( .ina ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, n2665}), .inb ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n1938}), .clk ( clk ), .rnd ({Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820], Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810]}), .outt ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n1939}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2024 ( .ina ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, n2235}), .inb ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n1943}), .clk ( clk ), .rnd ({Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830], Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825]}), .outt ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, n1948}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2032 ( .ina ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, n1946}), .inb ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, n1945}), .clk ( clk ), .rnd ({Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850], Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840]}), .outt ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, n1947}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2041 ( .ina ({new_AGEMA_signal_18571, new_AGEMA_signal_18567, new_AGEMA_signal_18563, new_AGEMA_signal_18559, new_AGEMA_signal_18555}), .inb ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, n1951}), .clk ( clk ), .rnd ({Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860], Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855]}), .outt ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n1954}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2049 ( .ina ({new_AGEMA_signal_18581, new_AGEMA_signal_18579, new_AGEMA_signal_18577, new_AGEMA_signal_18575, new_AGEMA_signal_18573}), .inb ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, n1952}), .clk ( clk ), .rnd ({Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880], Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870]}), .outt ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, n1953}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2058 ( .ina ({new_AGEMA_signal_18591, new_AGEMA_signal_18589, new_AGEMA_signal_18587, new_AGEMA_signal_18585, new_AGEMA_signal_18583}), .inb ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2687}), .clk ( clk ), .rnd ({Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890], Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885]}), .outt ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, n2658}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2065 ( .ina ({new_AGEMA_signal_18601, new_AGEMA_signal_18599, new_AGEMA_signal_18597, new_AGEMA_signal_18595, new_AGEMA_signal_18593}), .inb ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n1963}), .clk ( clk ), .rnd ({Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910], Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900]}), .outt ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, n1965}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2078 ( .ina ({new_AGEMA_signal_18611, new_AGEMA_signal_18609, new_AGEMA_signal_18607, new_AGEMA_signal_18605, new_AGEMA_signal_18603}), .inb ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, n1968}), .clk ( clk ), .rnd ({Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920], Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915]}), .outt ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, n1970}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2084 ( .ina ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, n2684}), .inb ({new_AGEMA_signal_18621, new_AGEMA_signal_18619, new_AGEMA_signal_18617, new_AGEMA_signal_18615, new_AGEMA_signal_18613}), .clk ( clk ), .rnd ({Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940], Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930]}), .outt ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, n1969}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2093 ( .ina ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n1972}), .inb ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n1971}), .clk ( clk ), .rnd ({Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950], Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945]}), .outt ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n1978}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2102 ( .ina ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, n1974}), .inb ({new_AGEMA_signal_18631, new_AGEMA_signal_18629, new_AGEMA_signal_18627, new_AGEMA_signal_18625, new_AGEMA_signal_18623}), .clk ( clk ), .rnd ({Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970], Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960]}), .outt ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, n1975}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2107 ( .ina ({new_AGEMA_signal_18641, new_AGEMA_signal_18639, new_AGEMA_signal_18637, new_AGEMA_signal_18635, new_AGEMA_signal_18633}), .inb ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, n1979}), .clk ( clk ), .rnd ({Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980], Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975]}), .outt ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, n1980}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2114 ( .ina ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n1985}), .inb ({new_AGEMA_signal_18651, new_AGEMA_signal_18649, new_AGEMA_signal_18647, new_AGEMA_signal_18645, new_AGEMA_signal_18643}), .clk ( clk ), .rnd ({Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000], Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990]}), .outt ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n1986}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2124 ( .ina ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, n1994}), .inb ({new_AGEMA_signal_18661, new_AGEMA_signal_18659, new_AGEMA_signal_18657, new_AGEMA_signal_18655, new_AGEMA_signal_18653}), .clk ( clk ), .rnd ({Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010], Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005]}), .outt ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, n1997}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2137 ( .ina ({new_AGEMA_signal_18671, new_AGEMA_signal_18669, new_AGEMA_signal_18667, new_AGEMA_signal_18665, new_AGEMA_signal_18663}), .inb ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2137}), .clk ( clk ), .rnd ({Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030], Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020]}), .outt ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, n2012}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2145 ( .ina ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, n2006}), .inb ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, n2005}), .clk ( clk ), .rnd ({Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040], Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035]}), .outt ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n2007}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2161 ( .ins ({new_AGEMA_signal_18681, new_AGEMA_signal_18679, new_AGEMA_signal_18677, new_AGEMA_signal_18675, new_AGEMA_signal_18673}), .inb ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, new_AGEMA_signal_1834, n2020}), .ina ({new_AGEMA_signal_18701, new_AGEMA_signal_18697, new_AGEMA_signal_18693, new_AGEMA_signal_18689, new_AGEMA_signal_18685}), .clk ( clk ), .rnd ({Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060], Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050]}), .outt ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, n2021}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2176 ( .ina ({new_AGEMA_signal_18711, new_AGEMA_signal_18709, new_AGEMA_signal_18707, new_AGEMA_signal_18705, new_AGEMA_signal_18703}), .inb ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n2031}), .clk ( clk ), .rnd ({Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070], Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065]}), .outt ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, n2032}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2185 ( .ina ({new_AGEMA_signal_18721, new_AGEMA_signal_18719, new_AGEMA_signal_18717, new_AGEMA_signal_18715, new_AGEMA_signal_18713}), .inb ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, n2040}), .clk ( clk ), .rnd ({Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090], Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080]}), .outt ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2041}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2189 ( .ina ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, n2665}), .inb ({new_AGEMA_signal_18731, new_AGEMA_signal_18729, new_AGEMA_signal_18727, new_AGEMA_signal_18725, new_AGEMA_signal_18723}), .clk ( clk ), .rnd ({Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100], Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095]}), .outt ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, n2043}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2194 ( .ina ({new_AGEMA_signal_18741, new_AGEMA_signal_18739, new_AGEMA_signal_18737, new_AGEMA_signal_18735, new_AGEMA_signal_18733}), .inb ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, n2045}), .clk ( clk ), .rnd ({Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120], Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110]}), .outt ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, new_AGEMA_signal_3146, n2046}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2204 ( .ins ({new_AGEMA_signal_18681, new_AGEMA_signal_18679, new_AGEMA_signal_18677, new_AGEMA_signal_18675, new_AGEMA_signal_18673}), .inb ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, n2056}), .ina ({new_AGEMA_signal_18751, new_AGEMA_signal_18749, new_AGEMA_signal_18747, new_AGEMA_signal_18745, new_AGEMA_signal_18743}), .clk ( clk ), .rnd ({Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130], Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125]}), .outt ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2058}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2210 ( .ina ({new_AGEMA_signal_18761, new_AGEMA_signal_18759, new_AGEMA_signal_18757, new_AGEMA_signal_18755, new_AGEMA_signal_18753}), .inb ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, n2060}), .clk ( clk ), .rnd ({Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150], Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140]}), .outt ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, n2063}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2218 ( .ina ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2066}), .inb ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, n2065}), .clk ( clk ), .rnd ({Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160], Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155]}), .outt ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, new_AGEMA_signal_3158, n2652}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2227 ( .ina ({new_AGEMA_signal_18771, new_AGEMA_signal_18769, new_AGEMA_signal_18767, new_AGEMA_signal_18765, new_AGEMA_signal_18763}), .inb ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n2074}), .clk ( clk ), .rnd ({Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180], Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170]}), .outt ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2076}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2236 ( .ina ({new_AGEMA_signal_18791, new_AGEMA_signal_18787, new_AGEMA_signal_18783, new_AGEMA_signal_18779, new_AGEMA_signal_18775}), .inb ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, n2082}), .clk ( clk ), .rnd ({Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190], Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185]}), .outt ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, n2105}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2241 ( .ina ({new_AGEMA_signal_18801, new_AGEMA_signal_18799, new_AGEMA_signal_18797, new_AGEMA_signal_18795, new_AGEMA_signal_18793}), .inb ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, n2084}), .clk ( clk ), .rnd ({Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210], Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200]}), .outt ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, new_AGEMA_signal_3170, n2099}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2243 ( .ina ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n2085}), .inb ({new_AGEMA_signal_18811, new_AGEMA_signal_18809, new_AGEMA_signal_18807, new_AGEMA_signal_18805, new_AGEMA_signal_18803}), .clk ( clk ), .rnd ({Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220], Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215]}), .outt ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2091}) ) ;
    and_HPC1 #(.security_order(4), .pipeline(1)) U2246 ( .ina ({new_AGEMA_signal_18821, new_AGEMA_signal_18819, new_AGEMA_signal_18817, new_AGEMA_signal_18815, new_AGEMA_signal_18813}), .inb ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, n2131}), .clk ( clk ), .rnd ({Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240], Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230]}), .outt ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, n2090}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2253 ( .ina ({new_AGEMA_signal_18831, new_AGEMA_signal_18829, new_AGEMA_signal_18827, new_AGEMA_signal_18825, new_AGEMA_signal_18823}), .inb ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2330}), .clk ( clk ), .rnd ({Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250], Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245]}), .outt ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, n2093}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2262 ( .ina ({new_AGEMA_signal_18841, new_AGEMA_signal_18839, new_AGEMA_signal_18837, new_AGEMA_signal_18835, new_AGEMA_signal_18833}), .inb ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2160}), .clk ( clk ), .rnd ({Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270], Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260]}), .outt ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2102}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2266 ( .ina ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, n2504}), .inb ({new_AGEMA_signal_18861, new_AGEMA_signal_18857, new_AGEMA_signal_18853, new_AGEMA_signal_18849, new_AGEMA_signal_18845}), .clk ( clk ), .rnd ({Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280], Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275]}), .outt ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, n2106}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2272 ( .ina ({new_AGEMA_signal_18871, new_AGEMA_signal_18869, new_AGEMA_signal_18867, new_AGEMA_signal_18865, new_AGEMA_signal_18863}), .inb ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, n2114}), .clk ( clk ), .rnd ({Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300], Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290]}), .outt ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, n2116}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2282 ( .ina ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, n2291}), .inb ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, new_AGEMA_signal_1942, n2119}), .clk ( clk ), .rnd ({Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310], Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305]}), .outt ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, n2120}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2293 ( .ina ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, n2130}), .inb ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, n2129}), .clk ( clk ), .rnd ({Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330], Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320]}), .outt ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2155}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2296 ( .ina ({new_AGEMA_signal_18881, new_AGEMA_signal_18879, new_AGEMA_signal_18877, new_AGEMA_signal_18875, new_AGEMA_signal_18873}), .inb ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, n2131}), .clk ( clk ), .rnd ({Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340], Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335]}), .outt ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2543}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2299 ( .ina ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, n2133}), .inb ({new_AGEMA_signal_18891, new_AGEMA_signal_18889, new_AGEMA_signal_18887, new_AGEMA_signal_18885, new_AGEMA_signal_18883}), .clk ( clk ), .rnd ({Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360], Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350]}), .outt ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, n2134}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2303 ( .ina ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2137}), .inb ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, n2136}), .clk ( clk ), .rnd ({Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370], Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365]}), .outt ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, n2143}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2308 ( .ina ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2139}), .inb ({new_AGEMA_signal_18911, new_AGEMA_signal_18907, new_AGEMA_signal_18903, new_AGEMA_signal_18899, new_AGEMA_signal_18895}), .clk ( clk ), .rnd ({Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390], Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380]}), .outt ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2140}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2324 ( .ina ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, n2157}), .inb ({new_AGEMA_signal_18921, new_AGEMA_signal_18919, new_AGEMA_signal_18917, new_AGEMA_signal_18915, new_AGEMA_signal_18913}), .clk ( clk ), .rnd ({Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400], Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395]}), .outt ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, n2159}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2326 ( .ina ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2160}), .inb ({new_AGEMA_signal_18931, new_AGEMA_signal_18929, new_AGEMA_signal_18927, new_AGEMA_signal_18925, new_AGEMA_signal_18923}), .clk ( clk ), .rnd ({Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420], Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410]}), .outt ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, n2161}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2330 ( .ina ({new_AGEMA_signal_18571, new_AGEMA_signal_18567, new_AGEMA_signal_18563, new_AGEMA_signal_18559, new_AGEMA_signal_18555}), .inb ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2163}), .clk ( clk ), .rnd ({Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430], Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425]}), .outt ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, n2164}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2345 ( .ina ({new_AGEMA_signal_18941, new_AGEMA_signal_18939, new_AGEMA_signal_18937, new_AGEMA_signal_18935, new_AGEMA_signal_18933}), .inb ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, n2177}), .clk ( clk ), .rnd ({Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450], Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440]}), .outt ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, n2179}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2359 ( .ina ({new_AGEMA_signal_18961, new_AGEMA_signal_18957, new_AGEMA_signal_18953, new_AGEMA_signal_18949, new_AGEMA_signal_18945}), .inb ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, n2191}), .clk ( clk ), .rnd ({Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460], Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455]}), .outt ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, n2192}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2370 ( .ina ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2201}), .inb ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2200}), .clk ( clk ), .rnd ({Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480], Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470]}), .outt ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, n2203}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2382 ( .ina ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, n2217}), .inb ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, new_AGEMA_signal_2014, n2216}), .clk ( clk ), .rnd ({Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490], Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485]}), .outt ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, n2224}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2388 ( .ina ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2222}), .inb ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, n2221}), .clk ( clk ), .rnd ({Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510], Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500]}), .outt ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2223}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2392 ( .ina ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, n2504}), .inb ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, n2226}), .clk ( clk ), .rnd ({Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520], Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515]}), .outt ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, n2229}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2399 ( .ina ({new_AGEMA_signal_18581, new_AGEMA_signal_18579, new_AGEMA_signal_18577, new_AGEMA_signal_18575, new_AGEMA_signal_18573}), .inb ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, new_AGEMA_signal_3254, n2233}), .clk ( clk ), .rnd ({Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540], Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530]}), .outt ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, n2234}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2410 ( .ina ({new_AGEMA_signal_18591, new_AGEMA_signal_18589, new_AGEMA_signal_18587, new_AGEMA_signal_18585, new_AGEMA_signal_18583}), .inb ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, n2244}), .clk ( clk ), .rnd ({Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550], Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545]}), .outt ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2246}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2418 ( .ina ({new_AGEMA_signal_18971, new_AGEMA_signal_18969, new_AGEMA_signal_18967, new_AGEMA_signal_18965, new_AGEMA_signal_18963}), .inb ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2253}), .clk ( clk ), .rnd ({Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570], Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560]}), .outt ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, n2254}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2425 ( .ina ({new_AGEMA_signal_18981, new_AGEMA_signal_18979, new_AGEMA_signal_18977, new_AGEMA_signal_18975, new_AGEMA_signal_18973}), .inb ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, n2260}), .clk ( clk ), .rnd ({Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580], Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575]}), .outt ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, new_AGEMA_signal_3266, n2263}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2434 ( .ina ({new_AGEMA_signal_18991, new_AGEMA_signal_18989, new_AGEMA_signal_18987, new_AGEMA_signal_18985, new_AGEMA_signal_18983}), .inb ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, n2265}), .clk ( clk ), .rnd ({Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600], Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590]}), .outt ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, n2267}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2438 ( .ina ({new_AGEMA_signal_18581, new_AGEMA_signal_18579, new_AGEMA_signal_18577, new_AGEMA_signal_18575, new_AGEMA_signal_18573}), .inb ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n2269}), .clk ( clk ), .rnd ({Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610], Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605]}), .outt ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2270}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2445 ( .ina ({new_AGEMA_signal_19001, new_AGEMA_signal_18999, new_AGEMA_signal_18997, new_AGEMA_signal_18995, new_AGEMA_signal_18993}), .inb ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, n2277}), .clk ( clk ), .rnd ({Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630], Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620]}), .outt ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, n2279}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2450 ( .ina ({new_AGEMA_signal_18701, new_AGEMA_signal_18697, new_AGEMA_signal_18693, new_AGEMA_signal_18689, new_AGEMA_signal_18685}), .inb ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n2282}), .clk ( clk ), .rnd ({Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640], Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635]}), .outt ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, n2283}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2453 ( .ina ({new_AGEMA_signal_18801, new_AGEMA_signal_18799, new_AGEMA_signal_18797, new_AGEMA_signal_18795, new_AGEMA_signal_18793}), .inb ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2284}), .clk ( clk ), .rnd ({Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660], Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650]}), .outt ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, n2285}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2457 ( .ina ({new_AGEMA_signal_18571, new_AGEMA_signal_18567, new_AGEMA_signal_18563, new_AGEMA_signal_18559, new_AGEMA_signal_18555}), .inb ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, n2459}), .clk ( clk ), .rnd ({Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670], Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665]}), .outt ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, n2686}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2460 ( .ina ({new_AGEMA_signal_18591, new_AGEMA_signal_18589, new_AGEMA_signal_18587, new_AGEMA_signal_18585, new_AGEMA_signal_18583}), .inb ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, n2288}), .clk ( clk ), .rnd ({Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690], Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680]}), .outt ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n2289}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2463 ( .ina ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2458}), .inb ({new_AGEMA_signal_19011, new_AGEMA_signal_19009, new_AGEMA_signal_19007, new_AGEMA_signal_19005, new_AGEMA_signal_19003}), .clk ( clk ), .rnd ({Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700], Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695]}), .outt ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, n2297}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2465 ( .ina ({new_AGEMA_signal_19021, new_AGEMA_signal_19019, new_AGEMA_signal_19017, new_AGEMA_signal_19015, new_AGEMA_signal_19013}), .inb ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, n2291}), .clk ( clk ), .rnd ({Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720], Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710]}), .outt ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, n2292}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2473 ( .ina ({new_AGEMA_signal_19031, new_AGEMA_signal_19029, new_AGEMA_signal_19027, new_AGEMA_signal_19025, new_AGEMA_signal_19023}), .inb ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, n2300}), .clk ( clk ), .rnd ({Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730], Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725]}), .outt ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2301}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2483 ( .ina ({new_AGEMA_signal_19041, new_AGEMA_signal_19039, new_AGEMA_signal_19037, new_AGEMA_signal_19035, new_AGEMA_signal_19033}), .inb ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, n2314}), .clk ( clk ), .rnd ({Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750], Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740]}), .outt ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, n2321}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2487 ( .ina ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, n2319}), .inb ({new_AGEMA_signal_19051, new_AGEMA_signal_19049, new_AGEMA_signal_19047, new_AGEMA_signal_19045, new_AGEMA_signal_19043}), .clk ( clk ), .rnd ({Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760], Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755]}), .outt ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n2320}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2493 ( .ina ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, n2326}), .inb ({new_AGEMA_signal_19061, new_AGEMA_signal_19059, new_AGEMA_signal_19057, new_AGEMA_signal_19055, new_AGEMA_signal_19053}), .clk ( clk ), .rnd ({Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780], Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770]}), .outt ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, new_AGEMA_signal_2762, n2334}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2497 ( .ina ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2329}), .inb ({new_AGEMA_signal_18701, new_AGEMA_signal_18697, new_AGEMA_signal_18693, new_AGEMA_signal_18689, new_AGEMA_signal_18685}), .clk ( clk ), .rnd ({Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790], Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785]}), .outt ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, n2332}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2498 ( .ina ({new_AGEMA_signal_19071, new_AGEMA_signal_19069, new_AGEMA_signal_19067, new_AGEMA_signal_19065, new_AGEMA_signal_19063}), .inb ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2330}), .clk ( clk ), .rnd ({Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810], Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800]}), .outt ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2331}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2502 ( .ina ({new_AGEMA_signal_19081, new_AGEMA_signal_19079, new_AGEMA_signal_19077, new_AGEMA_signal_19075, new_AGEMA_signal_19073}), .inb ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, n2335}), .clk ( clk ), .rnd ({Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820], Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815]}), .outt ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2336}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2508 ( .ina ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, n2341}), .inb ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, n2340}), .clk ( clk ), .rnd ({Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840], Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830]}), .outt ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, n2342}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2519 ( .ina ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2352}), .inb ({new_AGEMA_signal_19091, new_AGEMA_signal_19089, new_AGEMA_signal_19087, new_AGEMA_signal_19085, new_AGEMA_signal_19083}), .clk ( clk ), .rnd ({Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850], Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845]}), .outt ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, n2367}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2523 ( .ina ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2354}), .inb ({new_AGEMA_signal_19101, new_AGEMA_signal_19099, new_AGEMA_signal_19097, new_AGEMA_signal_19095, new_AGEMA_signal_19093}), .clk ( clk ), .rnd ({Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870], Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860]}), .outt ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2358}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2547 ( .ina ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, n2385}), .inb ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2384}), .clk ( clk ), .rnd ({Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880], Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875]}), .outt ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, n2387}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2555 ( .ina ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, n2391}), .inb ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, n2390}), .clk ( clk ), .rnd ({Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900], Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890]}), .outt ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2392}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2566 ( .ina ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, n2403}), .inb ({new_AGEMA_signal_19111, new_AGEMA_signal_19109, new_AGEMA_signal_19107, new_AGEMA_signal_19105, new_AGEMA_signal_19103}), .clk ( clk ), .rnd ({Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910], Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905]}), .outt ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2404}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2570 ( .ina ({new_AGEMA_signal_18761, new_AGEMA_signal_18759, new_AGEMA_signal_18757, new_AGEMA_signal_18755, new_AGEMA_signal_18753}), .inb ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, n2408}), .clk ( clk ), .rnd ({Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930], Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920]}), .outt ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, n2409}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2575 ( .ina ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, n2574}), .inb ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, n2413}), .clk ( clk ), .rnd ({Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940], Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935]}), .outt ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2414}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2578 ( .ina ({new_AGEMA_signal_19121, new_AGEMA_signal_19119, new_AGEMA_signal_19117, new_AGEMA_signal_19115, new_AGEMA_signal_19113}), .inb ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2416}), .clk ( clk ), .rnd ({Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960], Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950]}), .outt ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2418}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2589 ( .ina ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, n2689}), .inb ({new_AGEMA_signal_19131, new_AGEMA_signal_19129, new_AGEMA_signal_19127, new_AGEMA_signal_19125, new_AGEMA_signal_19123}), .clk ( clk ), .rnd ({Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970], Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965]}), .outt ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, new_AGEMA_signal_3362, n2432}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2592 ( .ina ({new_AGEMA_signal_19161, new_AGEMA_signal_19155, new_AGEMA_signal_19149, new_AGEMA_signal_19143, new_AGEMA_signal_19137}), .inb ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2434}), .clk ( clk ), .rnd ({Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990], Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980]}), .outt ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2435}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2601 ( .ina ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, n2445}), .inb ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2444}), .clk ( clk ), .rnd ({Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000], Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995]}), .outt ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2449}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2603 ( .ina ({new_AGEMA_signal_19041, new_AGEMA_signal_19039, new_AGEMA_signal_19037, new_AGEMA_signal_19035, new_AGEMA_signal_19033}), .inb ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, n2447}), .clk ( clk ), .rnd ({Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020], Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010]}), .outt ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, n2448}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2609 ( .ina ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, n2454}), .inb ({new_AGEMA_signal_19171, new_AGEMA_signal_19169, new_AGEMA_signal_19167, new_AGEMA_signal_19165, new_AGEMA_signal_19163}), .clk ( clk ), .rnd ({Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030], Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025]}), .outt ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, n2455}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2612 ( .ina ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2687}), .inb ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2458}), .clk ( clk ), .rnd ({Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050], Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040]}), .outt ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2460}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2618 ( .ina ({new_AGEMA_signal_19021, new_AGEMA_signal_19019, new_AGEMA_signal_19017, new_AGEMA_signal_19015, new_AGEMA_signal_19013}), .inb ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2465}), .clk ( clk ), .rnd ({Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060], Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055]}), .outt ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2466}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2629 ( .ina ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, n2476}), .inb ({new_AGEMA_signal_19181, new_AGEMA_signal_19179, new_AGEMA_signal_19177, new_AGEMA_signal_19175, new_AGEMA_signal_19173}), .clk ( clk ), .rnd ({Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080], Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070]}), .outt ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, n2477}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2634 ( .ina ({new_AGEMA_signal_18751, new_AGEMA_signal_18749, new_AGEMA_signal_18747, new_AGEMA_signal_18745, new_AGEMA_signal_18743}), .inb ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, n2481}), .clk ( clk ), .rnd ({Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090], Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085]}), .outt ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2482}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2640 ( .ina ({new_AGEMA_signal_19191, new_AGEMA_signal_19189, new_AGEMA_signal_19187, new_AGEMA_signal_19185, new_AGEMA_signal_19183}), .inb ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, n2486}), .clk ( clk ), .rnd ({Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110], Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100]}), .outt ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n2490}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2648 ( .ina ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, n2495}), .inb ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, n2494}), .clk ( clk ), .rnd ({Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120], Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115]}), .outt ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, n2496}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2654 ( .ina ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, n2504}), .inb ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2503}), .clk ( clk ), .rnd ({Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140], Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130]}), .outt ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, new_AGEMA_signal_3746, n2507}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2664 ( .ina ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n2518}), .inb ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, n2517}), .clk ( clk ), .rnd ({Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150], Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145]}), .outt ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, n2525}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2669 ( .ina ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, n2523}), .inb ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, n2522}), .clk ( clk ), .rnd ({Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170], Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160]}), .outt ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, n2524}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2676 ( .ina ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n2532}), .inb ({new_AGEMA_signal_19211, new_AGEMA_signal_19207, new_AGEMA_signal_19203, new_AGEMA_signal_19199, new_AGEMA_signal_19195}), .clk ( clk ), .rnd ({Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180], Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175]}), .outt ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2537}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2678 ( .ina ({new_AGEMA_signal_18761, new_AGEMA_signal_18759, new_AGEMA_signal_18757, new_AGEMA_signal_18755, new_AGEMA_signal_18753}), .inb ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, n2534}), .clk ( clk ), .rnd ({Fresh[8204], Fresh[8203], Fresh[8202], Fresh[8201], Fresh[8200], Fresh[8199], Fresh[8198], Fresh[8197], Fresh[8196], Fresh[8195], Fresh[8194], Fresh[8193], Fresh[8192], Fresh[8191], Fresh[8190]}), .outt ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, n2536}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2684 ( .ina ({new_AGEMA_signal_19221, new_AGEMA_signal_19219, new_AGEMA_signal_19217, new_AGEMA_signal_19215, new_AGEMA_signal_19213}), .inb ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2546}), .clk ( clk ), .rnd ({Fresh[8219], Fresh[8218], Fresh[8217], Fresh[8216], Fresh[8215], Fresh[8214], Fresh[8213], Fresh[8212], Fresh[8211], Fresh[8210], Fresh[8209], Fresh[8208], Fresh[8207], Fresh[8206], Fresh[8205]}), .outt ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, n2547}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2693 ( .ina ({new_AGEMA_signal_19231, new_AGEMA_signal_19229, new_AGEMA_signal_19227, new_AGEMA_signal_19225, new_AGEMA_signal_19223}), .inb ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2556}), .clk ( clk ), .rnd ({Fresh[8234], Fresh[8233], Fresh[8232], Fresh[8231], Fresh[8230], Fresh[8229], Fresh[8228], Fresh[8227], Fresh[8226], Fresh[8225], Fresh[8224], Fresh[8223], Fresh[8222], Fresh[8221], Fresh[8220]}), .outt ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, n2557}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2699 ( .ina ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, n2715}), .inb ({new_AGEMA_signal_19241, new_AGEMA_signal_19239, new_AGEMA_signal_19237, new_AGEMA_signal_19235, new_AGEMA_signal_19233}), .clk ( clk ), .rnd ({Fresh[8249], Fresh[8248], Fresh[8247], Fresh[8246], Fresh[8245], Fresh[8244], Fresh[8243], Fresh[8242], Fresh[8241], Fresh[8240], Fresh[8239], Fresh[8238], Fresh[8237], Fresh[8236], Fresh[8235]}), .outt ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n2565}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2704 ( .ina ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, n2574}), .inb ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2573}), .clk ( clk ), .rnd ({Fresh[8264], Fresh[8263], Fresh[8262], Fresh[8261], Fresh[8260], Fresh[8259], Fresh[8258], Fresh[8257], Fresh[8256], Fresh[8255], Fresh[8254], Fresh[8253], Fresh[8252], Fresh[8251], Fresh[8250]}), .outt ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, n2591}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2709 ( .ina ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, n2579}), .inb ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, n2578}), .clk ( clk ), .rnd ({Fresh[8279], Fresh[8278], Fresh[8277], Fresh[8276], Fresh[8275], Fresh[8274], Fresh[8273], Fresh[8272], Fresh[8271], Fresh[8270], Fresh[8269], Fresh[8268], Fresh[8267], Fresh[8266], Fresh[8265]}), .outt ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, n2580}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2727 ( .ina ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, n2601}), .inb ({new_AGEMA_signal_19261, new_AGEMA_signal_19257, new_AGEMA_signal_19253, new_AGEMA_signal_19249, new_AGEMA_signal_19245}), .clk ( clk ), .rnd ({Fresh[8294], Fresh[8293], Fresh[8292], Fresh[8291], Fresh[8290], Fresh[8289], Fresh[8288], Fresh[8287], Fresh[8286], Fresh[8285], Fresh[8284], Fresh[8283], Fresh[8282], Fresh[8281], Fresh[8280]}), .outt ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, n2602}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2738 ( .ina ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, n2618}), .inb ({new_AGEMA_signal_19271, new_AGEMA_signal_19269, new_AGEMA_signal_19267, new_AGEMA_signal_19265, new_AGEMA_signal_19263}), .clk ( clk ), .rnd ({Fresh[8309], Fresh[8308], Fresh[8307], Fresh[8306], Fresh[8305], Fresh[8304], Fresh[8303], Fresh[8302], Fresh[8301], Fresh[8300], Fresh[8299], Fresh[8298], Fresh[8297], Fresh[8296], Fresh[8295]}), .outt ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, n2619}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2744 ( .ina ({new_AGEMA_signal_18811, new_AGEMA_signal_18809, new_AGEMA_signal_18807, new_AGEMA_signal_18805, new_AGEMA_signal_18803}), .inb ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2626}), .clk ( clk ), .rnd ({Fresh[8324], Fresh[8323], Fresh[8322], Fresh[8321], Fresh[8320], Fresh[8319], Fresh[8318], Fresh[8317], Fresh[8316], Fresh[8315], Fresh[8314], Fresh[8313], Fresh[8312], Fresh[8311], Fresh[8310]}), .outt ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, n2628}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2753 ( .ina ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, n2644}), .inb ({new_AGEMA_signal_18881, new_AGEMA_signal_18879, new_AGEMA_signal_18877, new_AGEMA_signal_18875, new_AGEMA_signal_18873}), .clk ( clk ), .rnd ({Fresh[8339], Fresh[8338], Fresh[8337], Fresh[8336], Fresh[8335], Fresh[8334], Fresh[8333], Fresh[8332], Fresh[8331], Fresh[8330], Fresh[8329], Fresh[8328], Fresh[8327], Fresh[8326], Fresh[8325]}), .outt ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2649}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2755 ( .ina ({new_AGEMA_signal_19281, new_AGEMA_signal_19279, new_AGEMA_signal_19277, new_AGEMA_signal_19275, new_AGEMA_signal_19273}), .inb ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, n2646}), .clk ( clk ), .rnd ({Fresh[8354], Fresh[8353], Fresh[8352], Fresh[8351], Fresh[8350], Fresh[8349], Fresh[8348], Fresh[8347], Fresh[8346], Fresh[8345], Fresh[8344], Fresh[8343], Fresh[8342], Fresh[8341], Fresh[8340]}), .outt ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, n2648}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2765 ( .ina ({new_AGEMA_signal_18591, new_AGEMA_signal_18589, new_AGEMA_signal_18587, new_AGEMA_signal_18585, new_AGEMA_signal_18583}), .inb ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, n2663}), .clk ( clk ), .rnd ({Fresh[8369], Fresh[8368], Fresh[8367], Fresh[8366], Fresh[8365], Fresh[8364], Fresh[8363], Fresh[8362], Fresh[8361], Fresh[8360], Fresh[8359], Fresh[8358], Fresh[8357], Fresh[8356], Fresh[8355]}), .outt ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, n2664}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2771 ( .ina ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2675}), .inb ({new_AGEMA_signal_19291, new_AGEMA_signal_19289, new_AGEMA_signal_19287, new_AGEMA_signal_19285, new_AGEMA_signal_19283}), .clk ( clk ), .rnd ({Fresh[8384], Fresh[8383], Fresh[8382], Fresh[8381], Fresh[8380], Fresh[8379], Fresh[8378], Fresh[8377], Fresh[8376], Fresh[8375], Fresh[8374], Fresh[8373], Fresh[8372], Fresh[8371], Fresh[8370]}), .outt ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, n2681}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2773 ( .ina ({new_AGEMA_signal_18921, new_AGEMA_signal_18919, new_AGEMA_signal_18917, new_AGEMA_signal_18915, new_AGEMA_signal_18913}), .inb ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, n2678}), .clk ( clk ), .rnd ({Fresh[8399], Fresh[8398], Fresh[8397], Fresh[8396], Fresh[8395], Fresh[8394], Fresh[8393], Fresh[8392], Fresh[8391], Fresh[8390], Fresh[8389], Fresh[8388], Fresh[8387], Fresh[8386], Fresh[8385]}), .outt ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, n2680}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2776 ( .ina ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, n2684}), .inb ({new_AGEMA_signal_19301, new_AGEMA_signal_19299, new_AGEMA_signal_19297, new_AGEMA_signal_19295, new_AGEMA_signal_19293}), .clk ( clk ), .rnd ({Fresh[8414], Fresh[8413], Fresh[8412], Fresh[8411], Fresh[8410], Fresh[8409], Fresh[8408], Fresh[8407], Fresh[8406], Fresh[8405], Fresh[8404], Fresh[8403], Fresh[8402], Fresh[8401], Fresh[8400]}), .outt ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2685}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2778 ( .ina ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2687}), .inb ({new_AGEMA_signal_19221, new_AGEMA_signal_19219, new_AGEMA_signal_19217, new_AGEMA_signal_19215, new_AGEMA_signal_19213}), .clk ( clk ), .rnd ({Fresh[8429], Fresh[8428], Fresh[8427], Fresh[8426], Fresh[8425], Fresh[8424], Fresh[8423], Fresh[8422], Fresh[8421], Fresh[8420], Fresh[8419], Fresh[8418], Fresh[8417], Fresh[8416], Fresh[8415]}), .outt ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, n2698}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2779 ( .ina ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, n2689}), .inb ({new_AGEMA_signal_19231, new_AGEMA_signal_19229, new_AGEMA_signal_19227, new_AGEMA_signal_19225, new_AGEMA_signal_19223}), .clk ( clk ), .rnd ({Fresh[8444], Fresh[8443], Fresh[8442], Fresh[8441], Fresh[8440], Fresh[8439], Fresh[8438], Fresh[8437], Fresh[8436], Fresh[8435], Fresh[8434], Fresh[8433], Fresh[8432], Fresh[8431], Fresh[8430]}), .outt ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, n2692}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2793 ( .ina ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, n2715}), .inb ({new_AGEMA_signal_19311, new_AGEMA_signal_19309, new_AGEMA_signal_19307, new_AGEMA_signal_19305, new_AGEMA_signal_19303}), .clk ( clk ), .rnd ({Fresh[8459], Fresh[8458], Fresh[8457], Fresh[8456], Fresh[8455], Fresh[8454], Fresh[8453], Fresh[8452], Fresh[8451], Fresh[8450], Fresh[8449], Fresh[8448], Fresh[8447], Fresh[8446], Fresh[8445]}), .outt ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2716}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2800 ( .ina ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2727}), .inb ({new_AGEMA_signal_19321, new_AGEMA_signal_19319, new_AGEMA_signal_19317, new_AGEMA_signal_19315, new_AGEMA_signal_19313}), .clk ( clk ), .rnd ({Fresh[8474], Fresh[8473], Fresh[8472], Fresh[8471], Fresh[8470], Fresh[8469], Fresh[8468], Fresh[8467], Fresh[8466], Fresh[8465], Fresh[8464], Fresh[8463], Fresh[8462], Fresh[8461], Fresh[8460]}), .outt ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, n2728}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2804 ( .ina ({new_AGEMA_signal_19331, new_AGEMA_signal_19329, new_AGEMA_signal_19327, new_AGEMA_signal_19325, new_AGEMA_signal_19323}), .inb ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2733}), .clk ( clk ), .rnd ({Fresh[8489], Fresh[8488], Fresh[8487], Fresh[8486], Fresh[8485], Fresh[8484], Fresh[8483], Fresh[8482], Fresh[8481], Fresh[8480], Fresh[8479], Fresh[8478], Fresh[8477], Fresh[8476], Fresh[8475]}), .outt ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, n2735}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2808 ( .ina ({new_AGEMA_signal_18651, new_AGEMA_signal_18649, new_AGEMA_signal_18647, new_AGEMA_signal_18645, new_AGEMA_signal_18643}), .inb ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, n2740}), .clk ( clk ), .rnd ({Fresh[8504], Fresh[8503], Fresh[8502], Fresh[8501], Fresh[8500], Fresh[8499], Fresh[8498], Fresh[8497], Fresh[8496], Fresh[8495], Fresh[8494], Fresh[8493], Fresh[8492], Fresh[8491], Fresh[8490]}), .outt ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2743}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2813 ( .ina ({new_AGEMA_signal_19351, new_AGEMA_signal_19347, new_AGEMA_signal_19343, new_AGEMA_signal_19339, new_AGEMA_signal_19335}), .inb ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2749}), .clk ( clk ), .rnd ({Fresh[8519], Fresh[8518], Fresh[8517], Fresh[8516], Fresh[8515], Fresh[8514], Fresh[8513], Fresh[8512], Fresh[8511], Fresh[8510], Fresh[8509], Fresh[8508], Fresh[8507], Fresh[8506], Fresh[8505]}), .outt ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, n2751}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2817 ( .ina ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2757}), .inb ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, n2756}), .clk ( clk ), .rnd ({Fresh[8534], Fresh[8533], Fresh[8532], Fresh[8531], Fresh[8530], Fresh[8529], Fresh[8528], Fresh[8527], Fresh[8526], Fresh[8525], Fresh[8524], Fresh[8523], Fresh[8522], Fresh[8521], Fresh[8520]}), .outt ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, n2758}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2820 ( .ina ({new_AGEMA_signal_19361, new_AGEMA_signal_19359, new_AGEMA_signal_19357, new_AGEMA_signal_19355, new_AGEMA_signal_19353}), .inb ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, n2762}), .clk ( clk ), .rnd ({Fresh[8549], Fresh[8548], Fresh[8547], Fresh[8546], Fresh[8545], Fresh[8544], Fresh[8543], Fresh[8542], Fresh[8541], Fresh[8540], Fresh[8539], Fresh[8538], Fresh[8537], Fresh[8536], Fresh[8535]}), .outt ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, n2764}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2827 ( .ina ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2776}), .inb ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, n2775}), .clk ( clk ), .rnd ({Fresh[8564], Fresh[8563], Fresh[8562], Fresh[8561], Fresh[8560], Fresh[8559], Fresh[8558], Fresh[8557], Fresh[8556], Fresh[8555], Fresh[8554], Fresh[8553], Fresh[8552], Fresh[8551], Fresh[8550]}), .outt ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2800}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2831 ( .ina ({new_AGEMA_signal_19371, new_AGEMA_signal_19369, new_AGEMA_signal_19367, new_AGEMA_signal_19365, new_AGEMA_signal_19363}), .inb ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2783}), .clk ( clk ), .rnd ({Fresh[8579], Fresh[8578], Fresh[8577], Fresh[8576], Fresh[8575], Fresh[8574], Fresh[8573], Fresh[8572], Fresh[8571], Fresh[8570], Fresh[8569], Fresh[8568], Fresh[8567], Fresh[8566], Fresh[8565]}), .outt ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, new_AGEMA_signal_3038, n2788}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2837 ( .ina ({new_AGEMA_signal_19391, new_AGEMA_signal_19387, new_AGEMA_signal_19383, new_AGEMA_signal_19379, new_AGEMA_signal_19375}), .inb ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2795}), .clk ( clk ), .rnd ({Fresh[8594], Fresh[8593], Fresh[8592], Fresh[8591], Fresh[8590], Fresh[8589], Fresh[8588], Fresh[8587], Fresh[8586], Fresh[8585], Fresh[8584], Fresh[8583], Fresh[8582], Fresh[8581], Fresh[8580]}), .outt ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507, new_AGEMA_signal_3506, n2797}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2846 ( .ina ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, n2814}), .inb ({new_AGEMA_signal_18681, new_AGEMA_signal_18679, new_AGEMA_signal_18677, new_AGEMA_signal_18675, new_AGEMA_signal_18673}), .clk ( clk ), .rnd ({Fresh[8609], Fresh[8608], Fresh[8607], Fresh[8606], Fresh[8605], Fresh[8604], Fresh[8603], Fresh[8602], Fresh[8601], Fresh[8600], Fresh[8599], Fresh[8598], Fresh[8597], Fresh[8596], Fresh[8595]}), .outt ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2822}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2849 ( .ina ({new_AGEMA_signal_19401, new_AGEMA_signal_19399, new_AGEMA_signal_19397, new_AGEMA_signal_19395, new_AGEMA_signal_19393}), .inb ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, n2819}), .clk ( clk ), .rnd ({Fresh[8624], Fresh[8623], Fresh[8622], Fresh[8621], Fresh[8620], Fresh[8619], Fresh[8618], Fresh[8617], Fresh[8616], Fresh[8615], Fresh[8614], Fresh[8613], Fresh[8612], Fresh[8611], Fresh[8610]}), .outt ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C ( clk ), .D ( new_AGEMA_signal_19404 ), .Q ( new_AGEMA_signal_19405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C ( clk ), .D ( new_AGEMA_signal_19408 ), .Q ( new_AGEMA_signal_19409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C ( clk ), .D ( new_AGEMA_signal_19412 ), .Q ( new_AGEMA_signal_19413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C ( clk ), .D ( new_AGEMA_signal_19416 ), .Q ( new_AGEMA_signal_19417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C ( clk ), .D ( new_AGEMA_signal_19420 ), .Q ( new_AGEMA_signal_19421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C ( clk ), .D ( new_AGEMA_signal_19424 ), .Q ( new_AGEMA_signal_19425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C ( clk ), .D ( new_AGEMA_signal_19428 ), .Q ( new_AGEMA_signal_19429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C ( clk ), .D ( new_AGEMA_signal_19432 ), .Q ( new_AGEMA_signal_19433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C ( clk ), .D ( new_AGEMA_signal_19436 ), .Q ( new_AGEMA_signal_19437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C ( clk ), .D ( new_AGEMA_signal_19440 ), .Q ( new_AGEMA_signal_19441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C ( clk ), .D ( new_AGEMA_signal_19442 ), .Q ( new_AGEMA_signal_19443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C ( clk ), .D ( new_AGEMA_signal_19444 ), .Q ( new_AGEMA_signal_19445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C ( clk ), .D ( new_AGEMA_signal_19446 ), .Q ( new_AGEMA_signal_19447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C ( clk ), .D ( new_AGEMA_signal_19448 ), .Q ( new_AGEMA_signal_19449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C ( clk ), .D ( new_AGEMA_signal_19450 ), .Q ( new_AGEMA_signal_19451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C ( clk ), .D ( new_AGEMA_signal_19452 ), .Q ( new_AGEMA_signal_19453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C ( clk ), .D ( new_AGEMA_signal_19454 ), .Q ( new_AGEMA_signal_19455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C ( clk ), .D ( new_AGEMA_signal_19456 ), .Q ( new_AGEMA_signal_19457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C ( clk ), .D ( new_AGEMA_signal_19458 ), .Q ( new_AGEMA_signal_19459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C ( clk ), .D ( new_AGEMA_signal_19460 ), .Q ( new_AGEMA_signal_19461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C ( clk ), .D ( new_AGEMA_signal_19464 ), .Q ( new_AGEMA_signal_19465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C ( clk ), .D ( new_AGEMA_signal_19468 ), .Q ( new_AGEMA_signal_19469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C ( clk ), .D ( new_AGEMA_signal_19472 ), .Q ( new_AGEMA_signal_19473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C ( clk ), .D ( new_AGEMA_signal_19476 ), .Q ( new_AGEMA_signal_19477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C ( clk ), .D ( new_AGEMA_signal_19480 ), .Q ( new_AGEMA_signal_19481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C ( clk ), .D ( new_AGEMA_signal_19482 ), .Q ( new_AGEMA_signal_19483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C ( clk ), .D ( new_AGEMA_signal_19484 ), .Q ( new_AGEMA_signal_19485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C ( clk ), .D ( new_AGEMA_signal_19486 ), .Q ( new_AGEMA_signal_19487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C ( clk ), .D ( new_AGEMA_signal_19488 ), .Q ( new_AGEMA_signal_19489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C ( clk ), .D ( new_AGEMA_signal_19490 ), .Q ( new_AGEMA_signal_19491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C ( clk ), .D ( new_AGEMA_signal_19494 ), .Q ( new_AGEMA_signal_19495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C ( clk ), .D ( new_AGEMA_signal_19498 ), .Q ( new_AGEMA_signal_19499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C ( clk ), .D ( new_AGEMA_signal_19502 ), .Q ( new_AGEMA_signal_19503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C ( clk ), .D ( new_AGEMA_signal_19506 ), .Q ( new_AGEMA_signal_19507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C ( clk ), .D ( new_AGEMA_signal_19510 ), .Q ( new_AGEMA_signal_19511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C ( clk ), .D ( new_AGEMA_signal_19512 ), .Q ( new_AGEMA_signal_19513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C ( clk ), .D ( new_AGEMA_signal_19514 ), .Q ( new_AGEMA_signal_19515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C ( clk ), .D ( new_AGEMA_signal_19516 ), .Q ( new_AGEMA_signal_19517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C ( clk ), .D ( new_AGEMA_signal_19518 ), .Q ( new_AGEMA_signal_19519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C ( clk ), .D ( new_AGEMA_signal_19520 ), .Q ( new_AGEMA_signal_19521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C ( clk ), .D ( new_AGEMA_signal_19524 ), .Q ( new_AGEMA_signal_19525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C ( clk ), .D ( new_AGEMA_signal_19528 ), .Q ( new_AGEMA_signal_19529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C ( clk ), .D ( new_AGEMA_signal_19532 ), .Q ( new_AGEMA_signal_19533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C ( clk ), .D ( new_AGEMA_signal_19536 ), .Q ( new_AGEMA_signal_19537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C ( clk ), .D ( new_AGEMA_signal_19540 ), .Q ( new_AGEMA_signal_19541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C ( clk ), .D ( new_AGEMA_signal_19544 ), .Q ( new_AGEMA_signal_19545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C ( clk ), .D ( new_AGEMA_signal_19548 ), .Q ( new_AGEMA_signal_19549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C ( clk ), .D ( new_AGEMA_signal_19552 ), .Q ( new_AGEMA_signal_19553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C ( clk ), .D ( new_AGEMA_signal_19556 ), .Q ( new_AGEMA_signal_19557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C ( clk ), .D ( new_AGEMA_signal_19560 ), .Q ( new_AGEMA_signal_19561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C ( clk ), .D ( new_AGEMA_signal_19562 ), .Q ( new_AGEMA_signal_19563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C ( clk ), .D ( new_AGEMA_signal_19564 ), .Q ( new_AGEMA_signal_19565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C ( clk ), .D ( new_AGEMA_signal_19566 ), .Q ( new_AGEMA_signal_19567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C ( clk ), .D ( new_AGEMA_signal_19568 ), .Q ( new_AGEMA_signal_19569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C ( clk ), .D ( new_AGEMA_signal_19570 ), .Q ( new_AGEMA_signal_19571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C ( clk ), .D ( new_AGEMA_signal_19572 ), .Q ( new_AGEMA_signal_19573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C ( clk ), .D ( new_AGEMA_signal_19574 ), .Q ( new_AGEMA_signal_19575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C ( clk ), .D ( new_AGEMA_signal_19576 ), .Q ( new_AGEMA_signal_19577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C ( clk ), .D ( new_AGEMA_signal_19578 ), .Q ( new_AGEMA_signal_19579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C ( clk ), .D ( new_AGEMA_signal_19580 ), .Q ( new_AGEMA_signal_19581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C ( clk ), .D ( new_AGEMA_signal_19582 ), .Q ( new_AGEMA_signal_19583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C ( clk ), .D ( new_AGEMA_signal_19584 ), .Q ( new_AGEMA_signal_19585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C ( clk ), .D ( new_AGEMA_signal_19586 ), .Q ( new_AGEMA_signal_19587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C ( clk ), .D ( new_AGEMA_signal_19588 ), .Q ( new_AGEMA_signal_19589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C ( clk ), .D ( new_AGEMA_signal_19590 ), .Q ( new_AGEMA_signal_19591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C ( clk ), .D ( new_AGEMA_signal_19592 ), .Q ( new_AGEMA_signal_19593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C ( clk ), .D ( new_AGEMA_signal_19594 ), .Q ( new_AGEMA_signal_19595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C ( clk ), .D ( new_AGEMA_signal_19596 ), .Q ( new_AGEMA_signal_19597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C ( clk ), .D ( new_AGEMA_signal_19598 ), .Q ( new_AGEMA_signal_19599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C ( clk ), .D ( new_AGEMA_signal_19600 ), .Q ( new_AGEMA_signal_19601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C ( clk ), .D ( new_AGEMA_signal_19604 ), .Q ( new_AGEMA_signal_19605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C ( clk ), .D ( new_AGEMA_signal_19608 ), .Q ( new_AGEMA_signal_19609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C ( clk ), .D ( new_AGEMA_signal_19612 ), .Q ( new_AGEMA_signal_19613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C ( clk ), .D ( new_AGEMA_signal_19616 ), .Q ( new_AGEMA_signal_19617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C ( clk ), .D ( new_AGEMA_signal_19620 ), .Q ( new_AGEMA_signal_19621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C ( clk ), .D ( new_AGEMA_signal_19624 ), .Q ( new_AGEMA_signal_19625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C ( clk ), .D ( new_AGEMA_signal_19628 ), .Q ( new_AGEMA_signal_19629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C ( clk ), .D ( new_AGEMA_signal_19632 ), .Q ( new_AGEMA_signal_19633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C ( clk ), .D ( new_AGEMA_signal_19636 ), .Q ( new_AGEMA_signal_19637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C ( clk ), .D ( new_AGEMA_signal_19640 ), .Q ( new_AGEMA_signal_19641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C ( clk ), .D ( new_AGEMA_signal_19644 ), .Q ( new_AGEMA_signal_19645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C ( clk ), .D ( new_AGEMA_signal_19648 ), .Q ( new_AGEMA_signal_19649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C ( clk ), .D ( new_AGEMA_signal_19652 ), .Q ( new_AGEMA_signal_19653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C ( clk ), .D ( new_AGEMA_signal_19656 ), .Q ( new_AGEMA_signal_19657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C ( clk ), .D ( new_AGEMA_signal_19660 ), .Q ( new_AGEMA_signal_19661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C ( clk ), .D ( new_AGEMA_signal_19662 ), .Q ( new_AGEMA_signal_19663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C ( clk ), .D ( new_AGEMA_signal_19664 ), .Q ( new_AGEMA_signal_19665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C ( clk ), .D ( new_AGEMA_signal_19666 ), .Q ( new_AGEMA_signal_19667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C ( clk ), .D ( new_AGEMA_signal_19668 ), .Q ( new_AGEMA_signal_19669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C ( clk ), .D ( new_AGEMA_signal_19670 ), .Q ( new_AGEMA_signal_19671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C ( clk ), .D ( new_AGEMA_signal_19672 ), .Q ( new_AGEMA_signal_19673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C ( clk ), .D ( new_AGEMA_signal_19674 ), .Q ( new_AGEMA_signal_19675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C ( clk ), .D ( new_AGEMA_signal_19676 ), .Q ( new_AGEMA_signal_19677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C ( clk ), .D ( new_AGEMA_signal_19678 ), .Q ( new_AGEMA_signal_19679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C ( clk ), .D ( new_AGEMA_signal_19680 ), .Q ( new_AGEMA_signal_19681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C ( clk ), .D ( new_AGEMA_signal_19682 ), .Q ( new_AGEMA_signal_19683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C ( clk ), .D ( new_AGEMA_signal_19684 ), .Q ( new_AGEMA_signal_19685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C ( clk ), .D ( new_AGEMA_signal_19686 ), .Q ( new_AGEMA_signal_19687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C ( clk ), .D ( new_AGEMA_signal_19688 ), .Q ( new_AGEMA_signal_19689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C ( clk ), .D ( new_AGEMA_signal_19690 ), .Q ( new_AGEMA_signal_19691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C ( clk ), .D ( new_AGEMA_signal_19694 ), .Q ( new_AGEMA_signal_19695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C ( clk ), .D ( new_AGEMA_signal_19698 ), .Q ( new_AGEMA_signal_19699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C ( clk ), .D ( new_AGEMA_signal_19702 ), .Q ( new_AGEMA_signal_19703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C ( clk ), .D ( new_AGEMA_signal_19706 ), .Q ( new_AGEMA_signal_19707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C ( clk ), .D ( new_AGEMA_signal_19710 ), .Q ( new_AGEMA_signal_19711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C ( clk ), .D ( new_AGEMA_signal_19712 ), .Q ( new_AGEMA_signal_19713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C ( clk ), .D ( new_AGEMA_signal_19714 ), .Q ( new_AGEMA_signal_19715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C ( clk ), .D ( new_AGEMA_signal_19716 ), .Q ( new_AGEMA_signal_19717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C ( clk ), .D ( new_AGEMA_signal_19718 ), .Q ( new_AGEMA_signal_19719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C ( clk ), .D ( new_AGEMA_signal_19720 ), .Q ( new_AGEMA_signal_19721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C ( clk ), .D ( new_AGEMA_signal_19724 ), .Q ( new_AGEMA_signal_19725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C ( clk ), .D ( new_AGEMA_signal_19728 ), .Q ( new_AGEMA_signal_19729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C ( clk ), .D ( new_AGEMA_signal_19732 ), .Q ( new_AGEMA_signal_19733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C ( clk ), .D ( new_AGEMA_signal_19736 ), .Q ( new_AGEMA_signal_19737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C ( clk ), .D ( new_AGEMA_signal_19740 ), .Q ( new_AGEMA_signal_19741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C ( clk ), .D ( new_AGEMA_signal_19746 ), .Q ( new_AGEMA_signal_19747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C ( clk ), .D ( new_AGEMA_signal_19752 ), .Q ( new_AGEMA_signal_19753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C ( clk ), .D ( new_AGEMA_signal_19758 ), .Q ( new_AGEMA_signal_19759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C ( clk ), .D ( new_AGEMA_signal_19764 ), .Q ( new_AGEMA_signal_19765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C ( clk ), .D ( new_AGEMA_signal_19770 ), .Q ( new_AGEMA_signal_19771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C ( clk ), .D ( new_AGEMA_signal_19774 ), .Q ( new_AGEMA_signal_19775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C ( clk ), .D ( new_AGEMA_signal_19778 ), .Q ( new_AGEMA_signal_19779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C ( clk ), .D ( new_AGEMA_signal_19782 ), .Q ( new_AGEMA_signal_19783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C ( clk ), .D ( new_AGEMA_signal_19786 ), .Q ( new_AGEMA_signal_19787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C ( clk ), .D ( new_AGEMA_signal_19790 ), .Q ( new_AGEMA_signal_19791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C ( clk ), .D ( new_AGEMA_signal_19794 ), .Q ( new_AGEMA_signal_19795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C ( clk ), .D ( new_AGEMA_signal_19798 ), .Q ( new_AGEMA_signal_19799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C ( clk ), .D ( new_AGEMA_signal_19802 ), .Q ( new_AGEMA_signal_19803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C ( clk ), .D ( new_AGEMA_signal_19806 ), .Q ( new_AGEMA_signal_19807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C ( clk ), .D ( new_AGEMA_signal_19810 ), .Q ( new_AGEMA_signal_19811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C ( clk ), .D ( new_AGEMA_signal_19812 ), .Q ( new_AGEMA_signal_19813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C ( clk ), .D ( new_AGEMA_signal_19814 ), .Q ( new_AGEMA_signal_19815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C ( clk ), .D ( new_AGEMA_signal_19816 ), .Q ( new_AGEMA_signal_19817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C ( clk ), .D ( new_AGEMA_signal_19818 ), .Q ( new_AGEMA_signal_19819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C ( clk ), .D ( new_AGEMA_signal_19820 ), .Q ( new_AGEMA_signal_19821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C ( clk ), .D ( new_AGEMA_signal_19822 ), .Q ( new_AGEMA_signal_19823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C ( clk ), .D ( new_AGEMA_signal_19824 ), .Q ( new_AGEMA_signal_19825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C ( clk ), .D ( new_AGEMA_signal_19826 ), .Q ( new_AGEMA_signal_19827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C ( clk ), .D ( new_AGEMA_signal_19828 ), .Q ( new_AGEMA_signal_19829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C ( clk ), .D ( new_AGEMA_signal_19830 ), .Q ( new_AGEMA_signal_19831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C ( clk ), .D ( new_AGEMA_signal_19832 ), .Q ( new_AGEMA_signal_19833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C ( clk ), .D ( new_AGEMA_signal_19834 ), .Q ( new_AGEMA_signal_19835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C ( clk ), .D ( new_AGEMA_signal_19836 ), .Q ( new_AGEMA_signal_19837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C ( clk ), .D ( new_AGEMA_signal_19838 ), .Q ( new_AGEMA_signal_19839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C ( clk ), .D ( new_AGEMA_signal_19840 ), .Q ( new_AGEMA_signal_19841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C ( clk ), .D ( new_AGEMA_signal_19842 ), .Q ( new_AGEMA_signal_19843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C ( clk ), .D ( new_AGEMA_signal_19844 ), .Q ( new_AGEMA_signal_19845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C ( clk ), .D ( new_AGEMA_signal_19846 ), .Q ( new_AGEMA_signal_19847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C ( clk ), .D ( new_AGEMA_signal_19848 ), .Q ( new_AGEMA_signal_19849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C ( clk ), .D ( new_AGEMA_signal_19850 ), .Q ( new_AGEMA_signal_19851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C ( clk ), .D ( new_AGEMA_signal_19854 ), .Q ( new_AGEMA_signal_19855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C ( clk ), .D ( new_AGEMA_signal_19858 ), .Q ( new_AGEMA_signal_19859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C ( clk ), .D ( new_AGEMA_signal_19862 ), .Q ( new_AGEMA_signal_19863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C ( clk ), .D ( new_AGEMA_signal_19866 ), .Q ( new_AGEMA_signal_19867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C ( clk ), .D ( new_AGEMA_signal_19870 ), .Q ( new_AGEMA_signal_19871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C ( clk ), .D ( new_AGEMA_signal_19876 ), .Q ( new_AGEMA_signal_19877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C ( clk ), .D ( new_AGEMA_signal_19882 ), .Q ( new_AGEMA_signal_19883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C ( clk ), .D ( new_AGEMA_signal_19888 ), .Q ( new_AGEMA_signal_19889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C ( clk ), .D ( new_AGEMA_signal_19894 ), .Q ( new_AGEMA_signal_19895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C ( clk ), .D ( new_AGEMA_signal_19900 ), .Q ( new_AGEMA_signal_19901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C ( clk ), .D ( new_AGEMA_signal_19904 ), .Q ( new_AGEMA_signal_19905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C ( clk ), .D ( new_AGEMA_signal_19908 ), .Q ( new_AGEMA_signal_19909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C ( clk ), .D ( new_AGEMA_signal_19912 ), .Q ( new_AGEMA_signal_19913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C ( clk ), .D ( new_AGEMA_signal_19916 ), .Q ( new_AGEMA_signal_19917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C ( clk ), .D ( new_AGEMA_signal_19920 ), .Q ( new_AGEMA_signal_19921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C ( clk ), .D ( new_AGEMA_signal_19922 ), .Q ( new_AGEMA_signal_19923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C ( clk ), .D ( new_AGEMA_signal_19924 ), .Q ( new_AGEMA_signal_19925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C ( clk ), .D ( new_AGEMA_signal_19926 ), .Q ( new_AGEMA_signal_19927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C ( clk ), .D ( new_AGEMA_signal_19928 ), .Q ( new_AGEMA_signal_19929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C ( clk ), .D ( new_AGEMA_signal_19930 ), .Q ( new_AGEMA_signal_19931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C ( clk ), .D ( new_AGEMA_signal_19932 ), .Q ( new_AGEMA_signal_19933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C ( clk ), .D ( new_AGEMA_signal_19934 ), .Q ( new_AGEMA_signal_19935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C ( clk ), .D ( new_AGEMA_signal_19936 ), .Q ( new_AGEMA_signal_19937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C ( clk ), .D ( new_AGEMA_signal_19938 ), .Q ( new_AGEMA_signal_19939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C ( clk ), .D ( new_AGEMA_signal_19940 ), .Q ( new_AGEMA_signal_19941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C ( clk ), .D ( new_AGEMA_signal_19942 ), .Q ( new_AGEMA_signal_19943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C ( clk ), .D ( new_AGEMA_signal_19944 ), .Q ( new_AGEMA_signal_19945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C ( clk ), .D ( new_AGEMA_signal_19946 ), .Q ( new_AGEMA_signal_19947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C ( clk ), .D ( new_AGEMA_signal_19948 ), .Q ( new_AGEMA_signal_19949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C ( clk ), .D ( new_AGEMA_signal_19950 ), .Q ( new_AGEMA_signal_19951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C ( clk ), .D ( new_AGEMA_signal_19954 ), .Q ( new_AGEMA_signal_19955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C ( clk ), .D ( new_AGEMA_signal_19958 ), .Q ( new_AGEMA_signal_19959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C ( clk ), .D ( new_AGEMA_signal_19962 ), .Q ( new_AGEMA_signal_19963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C ( clk ), .D ( new_AGEMA_signal_19966 ), .Q ( new_AGEMA_signal_19967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C ( clk ), .D ( new_AGEMA_signal_19970 ), .Q ( new_AGEMA_signal_19971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C ( clk ), .D ( new_AGEMA_signal_19972 ), .Q ( new_AGEMA_signal_19973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C ( clk ), .D ( new_AGEMA_signal_19974 ), .Q ( new_AGEMA_signal_19975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C ( clk ), .D ( new_AGEMA_signal_19976 ), .Q ( new_AGEMA_signal_19977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C ( clk ), .D ( new_AGEMA_signal_19978 ), .Q ( new_AGEMA_signal_19979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C ( clk ), .D ( new_AGEMA_signal_19980 ), .Q ( new_AGEMA_signal_19981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C ( clk ), .D ( new_AGEMA_signal_19982 ), .Q ( new_AGEMA_signal_19983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C ( clk ), .D ( new_AGEMA_signal_19984 ), .Q ( new_AGEMA_signal_19985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C ( clk ), .D ( new_AGEMA_signal_19986 ), .Q ( new_AGEMA_signal_19987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C ( clk ), .D ( new_AGEMA_signal_19988 ), .Q ( new_AGEMA_signal_19989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C ( clk ), .D ( new_AGEMA_signal_19990 ), .Q ( new_AGEMA_signal_19991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C ( clk ), .D ( new_AGEMA_signal_19994 ), .Q ( new_AGEMA_signal_19995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C ( clk ), .D ( new_AGEMA_signal_19998 ), .Q ( new_AGEMA_signal_19999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C ( clk ), .D ( new_AGEMA_signal_20002 ), .Q ( new_AGEMA_signal_20003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C ( clk ), .D ( new_AGEMA_signal_20006 ), .Q ( new_AGEMA_signal_20007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C ( clk ), .D ( new_AGEMA_signal_20010 ), .Q ( new_AGEMA_signal_20011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C ( clk ), .D ( new_AGEMA_signal_20014 ), .Q ( new_AGEMA_signal_20015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C ( clk ), .D ( new_AGEMA_signal_20018 ), .Q ( new_AGEMA_signal_20019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C ( clk ), .D ( new_AGEMA_signal_20022 ), .Q ( new_AGEMA_signal_20023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C ( clk ), .D ( new_AGEMA_signal_20026 ), .Q ( new_AGEMA_signal_20027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C ( clk ), .D ( new_AGEMA_signal_20030 ), .Q ( new_AGEMA_signal_20031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C ( clk ), .D ( new_AGEMA_signal_20034 ), .Q ( new_AGEMA_signal_20035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C ( clk ), .D ( new_AGEMA_signal_20038 ), .Q ( new_AGEMA_signal_20039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C ( clk ), .D ( new_AGEMA_signal_20042 ), .Q ( new_AGEMA_signal_20043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C ( clk ), .D ( new_AGEMA_signal_20046 ), .Q ( new_AGEMA_signal_20047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C ( clk ), .D ( new_AGEMA_signal_20050 ), .Q ( new_AGEMA_signal_20051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C ( clk ), .D ( new_AGEMA_signal_20054 ), .Q ( new_AGEMA_signal_20055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C ( clk ), .D ( new_AGEMA_signal_20058 ), .Q ( new_AGEMA_signal_20059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C ( clk ), .D ( new_AGEMA_signal_20062 ), .Q ( new_AGEMA_signal_20063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C ( clk ), .D ( new_AGEMA_signal_20066 ), .Q ( new_AGEMA_signal_20067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C ( clk ), .D ( new_AGEMA_signal_20070 ), .Q ( new_AGEMA_signal_20071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C ( clk ), .D ( new_AGEMA_signal_20074 ), .Q ( new_AGEMA_signal_20075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C ( clk ), .D ( new_AGEMA_signal_20078 ), .Q ( new_AGEMA_signal_20079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C ( clk ), .D ( new_AGEMA_signal_20082 ), .Q ( new_AGEMA_signal_20083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C ( clk ), .D ( new_AGEMA_signal_20086 ), .Q ( new_AGEMA_signal_20087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C ( clk ), .D ( new_AGEMA_signal_20090 ), .Q ( new_AGEMA_signal_20091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C ( clk ), .D ( new_AGEMA_signal_20092 ), .Q ( new_AGEMA_signal_20093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C ( clk ), .D ( new_AGEMA_signal_20094 ), .Q ( new_AGEMA_signal_20095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C ( clk ), .D ( new_AGEMA_signal_20096 ), .Q ( new_AGEMA_signal_20097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C ( clk ), .D ( new_AGEMA_signal_20098 ), .Q ( new_AGEMA_signal_20099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C ( clk ), .D ( new_AGEMA_signal_20100 ), .Q ( new_AGEMA_signal_20101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C ( clk ), .D ( new_AGEMA_signal_20102 ), .Q ( new_AGEMA_signal_20103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C ( clk ), .D ( new_AGEMA_signal_20104 ), .Q ( new_AGEMA_signal_20105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C ( clk ), .D ( new_AGEMA_signal_20106 ), .Q ( new_AGEMA_signal_20107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C ( clk ), .D ( new_AGEMA_signal_20108 ), .Q ( new_AGEMA_signal_20109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C ( clk ), .D ( new_AGEMA_signal_20110 ), .Q ( new_AGEMA_signal_20111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C ( clk ), .D ( new_AGEMA_signal_20112 ), .Q ( new_AGEMA_signal_20113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C ( clk ), .D ( new_AGEMA_signal_20114 ), .Q ( new_AGEMA_signal_20115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C ( clk ), .D ( new_AGEMA_signal_20116 ), .Q ( new_AGEMA_signal_20117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C ( clk ), .D ( new_AGEMA_signal_20118 ), .Q ( new_AGEMA_signal_20119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C ( clk ), .D ( new_AGEMA_signal_20120 ), .Q ( new_AGEMA_signal_20121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C ( clk ), .D ( new_AGEMA_signal_20122 ), .Q ( new_AGEMA_signal_20123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C ( clk ), .D ( new_AGEMA_signal_20124 ), .Q ( new_AGEMA_signal_20125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C ( clk ), .D ( new_AGEMA_signal_20126 ), .Q ( new_AGEMA_signal_20127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C ( clk ), .D ( new_AGEMA_signal_20128 ), .Q ( new_AGEMA_signal_20129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C ( clk ), .D ( new_AGEMA_signal_20130 ), .Q ( new_AGEMA_signal_20131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C ( clk ), .D ( new_AGEMA_signal_20134 ), .Q ( new_AGEMA_signal_20135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C ( clk ), .D ( new_AGEMA_signal_20138 ), .Q ( new_AGEMA_signal_20139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C ( clk ), .D ( new_AGEMA_signal_20142 ), .Q ( new_AGEMA_signal_20143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C ( clk ), .D ( new_AGEMA_signal_20146 ), .Q ( new_AGEMA_signal_20147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C ( clk ), .D ( new_AGEMA_signal_20150 ), .Q ( new_AGEMA_signal_20151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C ( clk ), .D ( new_AGEMA_signal_20154 ), .Q ( new_AGEMA_signal_20155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C ( clk ), .D ( new_AGEMA_signal_20158 ), .Q ( new_AGEMA_signal_20159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C ( clk ), .D ( new_AGEMA_signal_20162 ), .Q ( new_AGEMA_signal_20163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C ( clk ), .D ( new_AGEMA_signal_20166 ), .Q ( new_AGEMA_signal_20167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C ( clk ), .D ( new_AGEMA_signal_20170 ), .Q ( new_AGEMA_signal_20171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C ( clk ), .D ( new_AGEMA_signal_20172 ), .Q ( new_AGEMA_signal_20173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C ( clk ), .D ( new_AGEMA_signal_20174 ), .Q ( new_AGEMA_signal_20175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C ( clk ), .D ( new_AGEMA_signal_20176 ), .Q ( new_AGEMA_signal_20177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C ( clk ), .D ( new_AGEMA_signal_20178 ), .Q ( new_AGEMA_signal_20179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C ( clk ), .D ( new_AGEMA_signal_20180 ), .Q ( new_AGEMA_signal_20181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C ( clk ), .D ( new_AGEMA_signal_20182 ), .Q ( new_AGEMA_signal_20183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C ( clk ), .D ( new_AGEMA_signal_20184 ), .Q ( new_AGEMA_signal_20185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C ( clk ), .D ( new_AGEMA_signal_20186 ), .Q ( new_AGEMA_signal_20187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C ( clk ), .D ( new_AGEMA_signal_20188 ), .Q ( new_AGEMA_signal_20189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C ( clk ), .D ( new_AGEMA_signal_20190 ), .Q ( new_AGEMA_signal_20191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C ( clk ), .D ( new_AGEMA_signal_20192 ), .Q ( new_AGEMA_signal_20193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C ( clk ), .D ( new_AGEMA_signal_20194 ), .Q ( new_AGEMA_signal_20195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C ( clk ), .D ( new_AGEMA_signal_20196 ), .Q ( new_AGEMA_signal_20197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C ( clk ), .D ( new_AGEMA_signal_20198 ), .Q ( new_AGEMA_signal_20199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C ( clk ), .D ( new_AGEMA_signal_20200 ), .Q ( new_AGEMA_signal_20201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C ( clk ), .D ( new_AGEMA_signal_20202 ), .Q ( new_AGEMA_signal_20203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C ( clk ), .D ( new_AGEMA_signal_20204 ), .Q ( new_AGEMA_signal_20205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C ( clk ), .D ( new_AGEMA_signal_20206 ), .Q ( new_AGEMA_signal_20207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C ( clk ), .D ( new_AGEMA_signal_20208 ), .Q ( new_AGEMA_signal_20209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C ( clk ), .D ( new_AGEMA_signal_20210 ), .Q ( new_AGEMA_signal_20211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C ( clk ), .D ( new_AGEMA_signal_20212 ), .Q ( new_AGEMA_signal_20213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C ( clk ), .D ( new_AGEMA_signal_20214 ), .Q ( new_AGEMA_signal_20215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C ( clk ), .D ( new_AGEMA_signal_20216 ), .Q ( new_AGEMA_signal_20217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C ( clk ), .D ( new_AGEMA_signal_20218 ), .Q ( new_AGEMA_signal_20219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C ( clk ), .D ( new_AGEMA_signal_20220 ), .Q ( new_AGEMA_signal_20221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C ( clk ), .D ( new_AGEMA_signal_20222 ), .Q ( new_AGEMA_signal_20223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C ( clk ), .D ( new_AGEMA_signal_20224 ), .Q ( new_AGEMA_signal_20225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C ( clk ), .D ( new_AGEMA_signal_20226 ), .Q ( new_AGEMA_signal_20227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C ( clk ), .D ( new_AGEMA_signal_20228 ), .Q ( new_AGEMA_signal_20229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C ( clk ), .D ( new_AGEMA_signal_20230 ), .Q ( new_AGEMA_signal_20231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C ( clk ), .D ( new_AGEMA_signal_20232 ), .Q ( new_AGEMA_signal_20233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C ( clk ), .D ( new_AGEMA_signal_20234 ), .Q ( new_AGEMA_signal_20235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C ( clk ), .D ( new_AGEMA_signal_20236 ), .Q ( new_AGEMA_signal_20237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C ( clk ), .D ( new_AGEMA_signal_20238 ), .Q ( new_AGEMA_signal_20239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C ( clk ), .D ( new_AGEMA_signal_20240 ), .Q ( new_AGEMA_signal_20241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C ( clk ), .D ( new_AGEMA_signal_20242 ), .Q ( new_AGEMA_signal_20243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C ( clk ), .D ( new_AGEMA_signal_20244 ), .Q ( new_AGEMA_signal_20245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C ( clk ), .D ( new_AGEMA_signal_20246 ), .Q ( new_AGEMA_signal_20247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C ( clk ), .D ( new_AGEMA_signal_20248 ), .Q ( new_AGEMA_signal_20249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C ( clk ), .D ( new_AGEMA_signal_20250 ), .Q ( new_AGEMA_signal_20251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C ( clk ), .D ( new_AGEMA_signal_20252 ), .Q ( new_AGEMA_signal_20253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C ( clk ), .D ( new_AGEMA_signal_20254 ), .Q ( new_AGEMA_signal_20255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C ( clk ), .D ( new_AGEMA_signal_20256 ), .Q ( new_AGEMA_signal_20257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C ( clk ), .D ( new_AGEMA_signal_20258 ), .Q ( new_AGEMA_signal_20259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C ( clk ), .D ( new_AGEMA_signal_20260 ), .Q ( new_AGEMA_signal_20261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C ( clk ), .D ( new_AGEMA_signal_20264 ), .Q ( new_AGEMA_signal_20265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C ( clk ), .D ( new_AGEMA_signal_20268 ), .Q ( new_AGEMA_signal_20269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C ( clk ), .D ( new_AGEMA_signal_20272 ), .Q ( new_AGEMA_signal_20273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C ( clk ), .D ( new_AGEMA_signal_20276 ), .Q ( new_AGEMA_signal_20277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C ( clk ), .D ( new_AGEMA_signal_20280 ), .Q ( new_AGEMA_signal_20281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C ( clk ), .D ( new_AGEMA_signal_20282 ), .Q ( new_AGEMA_signal_20283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C ( clk ), .D ( new_AGEMA_signal_20284 ), .Q ( new_AGEMA_signal_20285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C ( clk ), .D ( new_AGEMA_signal_20286 ), .Q ( new_AGEMA_signal_20287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C ( clk ), .D ( new_AGEMA_signal_20288 ), .Q ( new_AGEMA_signal_20289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C ( clk ), .D ( new_AGEMA_signal_20290 ), .Q ( new_AGEMA_signal_20291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C ( clk ), .D ( new_AGEMA_signal_20292 ), .Q ( new_AGEMA_signal_20293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C ( clk ), .D ( new_AGEMA_signal_20294 ), .Q ( new_AGEMA_signal_20295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C ( clk ), .D ( new_AGEMA_signal_20296 ), .Q ( new_AGEMA_signal_20297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C ( clk ), .D ( new_AGEMA_signal_20298 ), .Q ( new_AGEMA_signal_20299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C ( clk ), .D ( new_AGEMA_signal_20300 ), .Q ( new_AGEMA_signal_20301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C ( clk ), .D ( new_AGEMA_signal_20302 ), .Q ( new_AGEMA_signal_20303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C ( clk ), .D ( new_AGEMA_signal_20304 ), .Q ( new_AGEMA_signal_20305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C ( clk ), .D ( new_AGEMA_signal_20306 ), .Q ( new_AGEMA_signal_20307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C ( clk ), .D ( new_AGEMA_signal_20308 ), .Q ( new_AGEMA_signal_20309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C ( clk ), .D ( new_AGEMA_signal_20310 ), .Q ( new_AGEMA_signal_20311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C ( clk ), .D ( new_AGEMA_signal_20312 ), .Q ( new_AGEMA_signal_20313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C ( clk ), .D ( new_AGEMA_signal_20314 ), .Q ( new_AGEMA_signal_20315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C ( clk ), .D ( new_AGEMA_signal_20316 ), .Q ( new_AGEMA_signal_20317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C ( clk ), .D ( new_AGEMA_signal_20318 ), .Q ( new_AGEMA_signal_20319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C ( clk ), .D ( new_AGEMA_signal_20320 ), .Q ( new_AGEMA_signal_20321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C ( clk ), .D ( new_AGEMA_signal_20322 ), .Q ( new_AGEMA_signal_20323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C ( clk ), .D ( new_AGEMA_signal_20324 ), .Q ( new_AGEMA_signal_20325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C ( clk ), .D ( new_AGEMA_signal_20326 ), .Q ( new_AGEMA_signal_20327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C ( clk ), .D ( new_AGEMA_signal_20328 ), .Q ( new_AGEMA_signal_20329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C ( clk ), .D ( new_AGEMA_signal_20330 ), .Q ( new_AGEMA_signal_20331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C ( clk ), .D ( new_AGEMA_signal_20334 ), .Q ( new_AGEMA_signal_20335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C ( clk ), .D ( new_AGEMA_signal_20338 ), .Q ( new_AGEMA_signal_20339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C ( clk ), .D ( new_AGEMA_signal_20342 ), .Q ( new_AGEMA_signal_20343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C ( clk ), .D ( new_AGEMA_signal_20346 ), .Q ( new_AGEMA_signal_20347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C ( clk ), .D ( new_AGEMA_signal_20350 ), .Q ( new_AGEMA_signal_20351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C ( clk ), .D ( new_AGEMA_signal_20354 ), .Q ( new_AGEMA_signal_20355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C ( clk ), .D ( new_AGEMA_signal_20358 ), .Q ( new_AGEMA_signal_20359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C ( clk ), .D ( new_AGEMA_signal_20362 ), .Q ( new_AGEMA_signal_20363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C ( clk ), .D ( new_AGEMA_signal_20366 ), .Q ( new_AGEMA_signal_20367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C ( clk ), .D ( new_AGEMA_signal_20370 ), .Q ( new_AGEMA_signal_20371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C ( clk ), .D ( new_AGEMA_signal_20374 ), .Q ( new_AGEMA_signal_20375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C ( clk ), .D ( new_AGEMA_signal_20378 ), .Q ( new_AGEMA_signal_20379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C ( clk ), .D ( new_AGEMA_signal_20382 ), .Q ( new_AGEMA_signal_20383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C ( clk ), .D ( new_AGEMA_signal_20386 ), .Q ( new_AGEMA_signal_20387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C ( clk ), .D ( new_AGEMA_signal_20390 ), .Q ( new_AGEMA_signal_20391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C ( clk ), .D ( new_AGEMA_signal_20394 ), .Q ( new_AGEMA_signal_20395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C ( clk ), .D ( new_AGEMA_signal_20398 ), .Q ( new_AGEMA_signal_20399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C ( clk ), .D ( new_AGEMA_signal_20402 ), .Q ( new_AGEMA_signal_20403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C ( clk ), .D ( new_AGEMA_signal_20406 ), .Q ( new_AGEMA_signal_20407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C ( clk ), .D ( new_AGEMA_signal_20410 ), .Q ( new_AGEMA_signal_20411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C ( clk ), .D ( new_AGEMA_signal_20412 ), .Q ( new_AGEMA_signal_20413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C ( clk ), .D ( new_AGEMA_signal_20416 ), .Q ( new_AGEMA_signal_20417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C ( clk ), .D ( new_AGEMA_signal_20420 ), .Q ( new_AGEMA_signal_20421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C ( clk ), .D ( new_AGEMA_signal_20424 ), .Q ( new_AGEMA_signal_20425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C ( clk ), .D ( new_AGEMA_signal_20428 ), .Q ( new_AGEMA_signal_20429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C ( clk ), .D ( new_AGEMA_signal_20432 ), .Q ( new_AGEMA_signal_20433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C ( clk ), .D ( new_AGEMA_signal_20436 ), .Q ( new_AGEMA_signal_20437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C ( clk ), .D ( new_AGEMA_signal_20440 ), .Q ( new_AGEMA_signal_20441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C ( clk ), .D ( new_AGEMA_signal_20444 ), .Q ( new_AGEMA_signal_20445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C ( clk ), .D ( new_AGEMA_signal_20448 ), .Q ( new_AGEMA_signal_20449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C ( clk ), .D ( new_AGEMA_signal_20456 ), .Q ( new_AGEMA_signal_20457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C ( clk ), .D ( new_AGEMA_signal_20464 ), .Q ( new_AGEMA_signal_20465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C ( clk ), .D ( new_AGEMA_signal_20472 ), .Q ( new_AGEMA_signal_20473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C ( clk ), .D ( new_AGEMA_signal_20480 ), .Q ( new_AGEMA_signal_20481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C ( clk ), .D ( new_AGEMA_signal_20488 ), .Q ( new_AGEMA_signal_20489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C ( clk ), .D ( new_AGEMA_signal_20506 ), .Q ( new_AGEMA_signal_20507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C ( clk ), .D ( new_AGEMA_signal_20514 ), .Q ( new_AGEMA_signal_20515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C ( clk ), .D ( new_AGEMA_signal_20522 ), .Q ( new_AGEMA_signal_20523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C ( clk ), .D ( new_AGEMA_signal_20530 ), .Q ( new_AGEMA_signal_20531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C ( clk ), .D ( new_AGEMA_signal_20538 ), .Q ( new_AGEMA_signal_20539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C ( clk ), .D ( new_AGEMA_signal_20544 ), .Q ( new_AGEMA_signal_20545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C ( clk ), .D ( new_AGEMA_signal_20550 ), .Q ( new_AGEMA_signal_20551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C ( clk ), .D ( new_AGEMA_signal_20556 ), .Q ( new_AGEMA_signal_20557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C ( clk ), .D ( new_AGEMA_signal_20562 ), .Q ( new_AGEMA_signal_20563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C ( clk ), .D ( new_AGEMA_signal_20568 ), .Q ( new_AGEMA_signal_20569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C ( clk ), .D ( new_AGEMA_signal_20572 ), .Q ( new_AGEMA_signal_20573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C ( clk ), .D ( new_AGEMA_signal_20576 ), .Q ( new_AGEMA_signal_20577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C ( clk ), .D ( new_AGEMA_signal_20580 ), .Q ( new_AGEMA_signal_20581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C ( clk ), .D ( new_AGEMA_signal_20584 ), .Q ( new_AGEMA_signal_20585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C ( clk ), .D ( new_AGEMA_signal_20588 ), .Q ( new_AGEMA_signal_20589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C ( clk ), .D ( new_AGEMA_signal_20594 ), .Q ( new_AGEMA_signal_20595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C ( clk ), .D ( new_AGEMA_signal_20600 ), .Q ( new_AGEMA_signal_20601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C ( clk ), .D ( new_AGEMA_signal_20606 ), .Q ( new_AGEMA_signal_20607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C ( clk ), .D ( new_AGEMA_signal_20612 ), .Q ( new_AGEMA_signal_20613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C ( clk ), .D ( new_AGEMA_signal_20618 ), .Q ( new_AGEMA_signal_20619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C ( clk ), .D ( new_AGEMA_signal_20634 ), .Q ( new_AGEMA_signal_20635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C ( clk ), .D ( new_AGEMA_signal_20640 ), .Q ( new_AGEMA_signal_20641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C ( clk ), .D ( new_AGEMA_signal_20646 ), .Q ( new_AGEMA_signal_20647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C ( clk ), .D ( new_AGEMA_signal_20652 ), .Q ( new_AGEMA_signal_20653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C ( clk ), .D ( new_AGEMA_signal_20658 ), .Q ( new_AGEMA_signal_20659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C ( clk ), .D ( new_AGEMA_signal_20664 ), .Q ( new_AGEMA_signal_20665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C ( clk ), .D ( new_AGEMA_signal_20670 ), .Q ( new_AGEMA_signal_20671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C ( clk ), .D ( new_AGEMA_signal_20676 ), .Q ( new_AGEMA_signal_20677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C ( clk ), .D ( new_AGEMA_signal_20682 ), .Q ( new_AGEMA_signal_20683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C ( clk ), .D ( new_AGEMA_signal_20688 ), .Q ( new_AGEMA_signal_20689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C ( clk ), .D ( new_AGEMA_signal_20702 ), .Q ( new_AGEMA_signal_20703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C ( clk ), .D ( new_AGEMA_signal_20706 ), .Q ( new_AGEMA_signal_20707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C ( clk ), .D ( new_AGEMA_signal_20710 ), .Q ( new_AGEMA_signal_20711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C ( clk ), .D ( new_AGEMA_signal_20714 ), .Q ( new_AGEMA_signal_20715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C ( clk ), .D ( new_AGEMA_signal_20718 ), .Q ( new_AGEMA_signal_20719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C ( clk ), .D ( new_AGEMA_signal_20724 ), .Q ( new_AGEMA_signal_20725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C ( clk ), .D ( new_AGEMA_signal_20730 ), .Q ( new_AGEMA_signal_20731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C ( clk ), .D ( new_AGEMA_signal_20736 ), .Q ( new_AGEMA_signal_20737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C ( clk ), .D ( new_AGEMA_signal_20742 ), .Q ( new_AGEMA_signal_20743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C ( clk ), .D ( new_AGEMA_signal_20748 ), .Q ( new_AGEMA_signal_20749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C ( clk ), .D ( new_AGEMA_signal_20754 ), .Q ( new_AGEMA_signal_20755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C ( clk ), .D ( new_AGEMA_signal_20760 ), .Q ( new_AGEMA_signal_20761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C ( clk ), .D ( new_AGEMA_signal_20766 ), .Q ( new_AGEMA_signal_20767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C ( clk ), .D ( new_AGEMA_signal_20772 ), .Q ( new_AGEMA_signal_20773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C ( clk ), .D ( new_AGEMA_signal_20778 ), .Q ( new_AGEMA_signal_20779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C ( clk ), .D ( new_AGEMA_signal_20794 ), .Q ( new_AGEMA_signal_20795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C ( clk ), .D ( new_AGEMA_signal_20800 ), .Q ( new_AGEMA_signal_20801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C ( clk ), .D ( new_AGEMA_signal_20806 ), .Q ( new_AGEMA_signal_20807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C ( clk ), .D ( new_AGEMA_signal_20812 ), .Q ( new_AGEMA_signal_20813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C ( clk ), .D ( new_AGEMA_signal_20818 ), .Q ( new_AGEMA_signal_20819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C ( clk ), .D ( new_AGEMA_signal_20832 ), .Q ( new_AGEMA_signal_20833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C ( clk ), .D ( new_AGEMA_signal_20836 ), .Q ( new_AGEMA_signal_20837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C ( clk ), .D ( new_AGEMA_signal_20840 ), .Q ( new_AGEMA_signal_20841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C ( clk ), .D ( new_AGEMA_signal_20844 ), .Q ( new_AGEMA_signal_20845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C ( clk ), .D ( new_AGEMA_signal_20848 ), .Q ( new_AGEMA_signal_20849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C ( clk ), .D ( new_AGEMA_signal_20852 ), .Q ( new_AGEMA_signal_20853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C ( clk ), .D ( new_AGEMA_signal_20856 ), .Q ( new_AGEMA_signal_20857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C ( clk ), .D ( new_AGEMA_signal_20860 ), .Q ( new_AGEMA_signal_20861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C ( clk ), .D ( new_AGEMA_signal_20864 ), .Q ( new_AGEMA_signal_20865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C ( clk ), .D ( new_AGEMA_signal_20868 ), .Q ( new_AGEMA_signal_20869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C ( clk ), .D ( new_AGEMA_signal_20886 ), .Q ( new_AGEMA_signal_20887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C ( clk ), .D ( new_AGEMA_signal_20894 ), .Q ( new_AGEMA_signal_20895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C ( clk ), .D ( new_AGEMA_signal_20902 ), .Q ( new_AGEMA_signal_20903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C ( clk ), .D ( new_AGEMA_signal_20910 ), .Q ( new_AGEMA_signal_20911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C ( clk ), .D ( new_AGEMA_signal_20918 ), .Q ( new_AGEMA_signal_20919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C ( clk ), .D ( new_AGEMA_signal_20924 ), .Q ( new_AGEMA_signal_20925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C ( clk ), .D ( new_AGEMA_signal_20930 ), .Q ( new_AGEMA_signal_20931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C ( clk ), .D ( new_AGEMA_signal_20936 ), .Q ( new_AGEMA_signal_20937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C ( clk ), .D ( new_AGEMA_signal_20942 ), .Q ( new_AGEMA_signal_20943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C ( clk ), .D ( new_AGEMA_signal_20948 ), .Q ( new_AGEMA_signal_20949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C ( clk ), .D ( new_AGEMA_signal_20952 ), .Q ( new_AGEMA_signal_20953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C ( clk ), .D ( new_AGEMA_signal_20956 ), .Q ( new_AGEMA_signal_20957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C ( clk ), .D ( new_AGEMA_signal_20960 ), .Q ( new_AGEMA_signal_20961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C ( clk ), .D ( new_AGEMA_signal_20964 ), .Q ( new_AGEMA_signal_20965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C ( clk ), .D ( new_AGEMA_signal_20968 ), .Q ( new_AGEMA_signal_20969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C ( clk ), .D ( new_AGEMA_signal_20972 ), .Q ( new_AGEMA_signal_20973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C ( clk ), .D ( new_AGEMA_signal_20976 ), .Q ( new_AGEMA_signal_20977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C ( clk ), .D ( new_AGEMA_signal_20980 ), .Q ( new_AGEMA_signal_20981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C ( clk ), .D ( new_AGEMA_signal_20984 ), .Q ( new_AGEMA_signal_20985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C ( clk ), .D ( new_AGEMA_signal_20988 ), .Q ( new_AGEMA_signal_20989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C ( clk ), .D ( new_AGEMA_signal_21012 ), .Q ( new_AGEMA_signal_21013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C ( clk ), .D ( new_AGEMA_signal_21016 ), .Q ( new_AGEMA_signal_21017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C ( clk ), .D ( new_AGEMA_signal_21020 ), .Q ( new_AGEMA_signal_21021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C ( clk ), .D ( new_AGEMA_signal_21024 ), .Q ( new_AGEMA_signal_21025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C ( clk ), .D ( new_AGEMA_signal_21028 ), .Q ( new_AGEMA_signal_21029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C ( clk ), .D ( new_AGEMA_signal_21032 ), .Q ( new_AGEMA_signal_21033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C ( clk ), .D ( new_AGEMA_signal_21036 ), .Q ( new_AGEMA_signal_21037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C ( clk ), .D ( new_AGEMA_signal_21040 ), .Q ( new_AGEMA_signal_21041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C ( clk ), .D ( new_AGEMA_signal_21044 ), .Q ( new_AGEMA_signal_21045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C ( clk ), .D ( new_AGEMA_signal_21048 ), .Q ( new_AGEMA_signal_21049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C ( clk ), .D ( new_AGEMA_signal_21064 ), .Q ( new_AGEMA_signal_21065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C ( clk ), .D ( new_AGEMA_signal_21070 ), .Q ( new_AGEMA_signal_21071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C ( clk ), .D ( new_AGEMA_signal_21076 ), .Q ( new_AGEMA_signal_21077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C ( clk ), .D ( new_AGEMA_signal_21082 ), .Q ( new_AGEMA_signal_21083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C ( clk ), .D ( new_AGEMA_signal_21088 ), .Q ( new_AGEMA_signal_21089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C ( clk ), .D ( new_AGEMA_signal_21092 ), .Q ( new_AGEMA_signal_21093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C ( clk ), .D ( new_AGEMA_signal_21096 ), .Q ( new_AGEMA_signal_21097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C ( clk ), .D ( new_AGEMA_signal_21100 ), .Q ( new_AGEMA_signal_21101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C ( clk ), .D ( new_AGEMA_signal_21104 ), .Q ( new_AGEMA_signal_21105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C ( clk ), .D ( new_AGEMA_signal_21108 ), .Q ( new_AGEMA_signal_21109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C ( clk ), .D ( new_AGEMA_signal_21122 ), .Q ( new_AGEMA_signal_21123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C ( clk ), .D ( new_AGEMA_signal_21126 ), .Q ( new_AGEMA_signal_21127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C ( clk ), .D ( new_AGEMA_signal_21130 ), .Q ( new_AGEMA_signal_21131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C ( clk ), .D ( new_AGEMA_signal_21134 ), .Q ( new_AGEMA_signal_21135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C ( clk ), .D ( new_AGEMA_signal_21138 ), .Q ( new_AGEMA_signal_21139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C ( clk ), .D ( new_AGEMA_signal_21142 ), .Q ( new_AGEMA_signal_21143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C ( clk ), .D ( new_AGEMA_signal_21146 ), .Q ( new_AGEMA_signal_21147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C ( clk ), .D ( new_AGEMA_signal_21150 ), .Q ( new_AGEMA_signal_21151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C ( clk ), .D ( new_AGEMA_signal_21154 ), .Q ( new_AGEMA_signal_21155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C ( clk ), .D ( new_AGEMA_signal_21158 ), .Q ( new_AGEMA_signal_21159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C ( clk ), .D ( new_AGEMA_signal_21162 ), .Q ( new_AGEMA_signal_21163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C ( clk ), .D ( new_AGEMA_signal_21166 ), .Q ( new_AGEMA_signal_21167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C ( clk ), .D ( new_AGEMA_signal_21170 ), .Q ( new_AGEMA_signal_21171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C ( clk ), .D ( new_AGEMA_signal_21174 ), .Q ( new_AGEMA_signal_21175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C ( clk ), .D ( new_AGEMA_signal_21178 ), .Q ( new_AGEMA_signal_21179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C ( clk ), .D ( new_AGEMA_signal_21192 ), .Q ( new_AGEMA_signal_21193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C ( clk ), .D ( new_AGEMA_signal_21196 ), .Q ( new_AGEMA_signal_21197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C ( clk ), .D ( new_AGEMA_signal_21200 ), .Q ( new_AGEMA_signal_21201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C ( clk ), .D ( new_AGEMA_signal_21204 ), .Q ( new_AGEMA_signal_21205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C ( clk ), .D ( new_AGEMA_signal_21208 ), .Q ( new_AGEMA_signal_21209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C ( clk ), .D ( new_AGEMA_signal_21224 ), .Q ( new_AGEMA_signal_21225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C ( clk ), .D ( new_AGEMA_signal_21230 ), .Q ( new_AGEMA_signal_21231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C ( clk ), .D ( new_AGEMA_signal_21236 ), .Q ( new_AGEMA_signal_21237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C ( clk ), .D ( new_AGEMA_signal_21242 ), .Q ( new_AGEMA_signal_21243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C ( clk ), .D ( new_AGEMA_signal_21248 ), .Q ( new_AGEMA_signal_21249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C ( clk ), .D ( new_AGEMA_signal_21254 ), .Q ( new_AGEMA_signal_21255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C ( clk ), .D ( new_AGEMA_signal_21260 ), .Q ( new_AGEMA_signal_21261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C ( clk ), .D ( new_AGEMA_signal_21266 ), .Q ( new_AGEMA_signal_21267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C ( clk ), .D ( new_AGEMA_signal_21272 ), .Q ( new_AGEMA_signal_21273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C ( clk ), .D ( new_AGEMA_signal_21278 ), .Q ( new_AGEMA_signal_21279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C ( clk ), .D ( new_AGEMA_signal_21282 ), .Q ( new_AGEMA_signal_21283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C ( clk ), .D ( new_AGEMA_signal_21286 ), .Q ( new_AGEMA_signal_21287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C ( clk ), .D ( new_AGEMA_signal_21290 ), .Q ( new_AGEMA_signal_21291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C ( clk ), .D ( new_AGEMA_signal_21294 ), .Q ( new_AGEMA_signal_21295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C ( clk ), .D ( new_AGEMA_signal_21298 ), .Q ( new_AGEMA_signal_21299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C ( clk ), .D ( new_AGEMA_signal_21316 ), .Q ( new_AGEMA_signal_21317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C ( clk ), .D ( new_AGEMA_signal_21324 ), .Q ( new_AGEMA_signal_21325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C ( clk ), .D ( new_AGEMA_signal_21332 ), .Q ( new_AGEMA_signal_21333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C ( clk ), .D ( new_AGEMA_signal_21340 ), .Q ( new_AGEMA_signal_21341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C ( clk ), .D ( new_AGEMA_signal_21348 ), .Q ( new_AGEMA_signal_21349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C ( clk ), .D ( new_AGEMA_signal_21362 ), .Q ( new_AGEMA_signal_21363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C ( clk ), .D ( new_AGEMA_signal_21366 ), .Q ( new_AGEMA_signal_21367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C ( clk ), .D ( new_AGEMA_signal_21370 ), .Q ( new_AGEMA_signal_21371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C ( clk ), .D ( new_AGEMA_signal_21374 ), .Q ( new_AGEMA_signal_21375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C ( clk ), .D ( new_AGEMA_signal_21378 ), .Q ( new_AGEMA_signal_21379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C ( clk ), .D ( new_AGEMA_signal_21382 ), .Q ( new_AGEMA_signal_21383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C ( clk ), .D ( new_AGEMA_signal_21386 ), .Q ( new_AGEMA_signal_21387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C ( clk ), .D ( new_AGEMA_signal_21390 ), .Q ( new_AGEMA_signal_21391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C ( clk ), .D ( new_AGEMA_signal_21394 ), .Q ( new_AGEMA_signal_21395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C ( clk ), .D ( new_AGEMA_signal_21398 ), .Q ( new_AGEMA_signal_21399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C ( clk ), .D ( new_AGEMA_signal_21402 ), .Q ( new_AGEMA_signal_21403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C ( clk ), .D ( new_AGEMA_signal_21406 ), .Q ( new_AGEMA_signal_21407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C ( clk ), .D ( new_AGEMA_signal_21410 ), .Q ( new_AGEMA_signal_21411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C ( clk ), .D ( new_AGEMA_signal_21414 ), .Q ( new_AGEMA_signal_21415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C ( clk ), .D ( new_AGEMA_signal_21418 ), .Q ( new_AGEMA_signal_21419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C ( clk ), .D ( new_AGEMA_signal_21422 ), .Q ( new_AGEMA_signal_21423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C ( clk ), .D ( new_AGEMA_signal_21426 ), .Q ( new_AGEMA_signal_21427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C ( clk ), .D ( new_AGEMA_signal_21430 ), .Q ( new_AGEMA_signal_21431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C ( clk ), .D ( new_AGEMA_signal_21434 ), .Q ( new_AGEMA_signal_21435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C ( clk ), .D ( new_AGEMA_signal_21438 ), .Q ( new_AGEMA_signal_21439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C ( clk ), .D ( new_AGEMA_signal_21442 ), .Q ( new_AGEMA_signal_21443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C ( clk ), .D ( new_AGEMA_signal_21446 ), .Q ( new_AGEMA_signal_21447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C ( clk ), .D ( new_AGEMA_signal_21450 ), .Q ( new_AGEMA_signal_21451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C ( clk ), .D ( new_AGEMA_signal_21454 ), .Q ( new_AGEMA_signal_21455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C ( clk ), .D ( new_AGEMA_signal_21458 ), .Q ( new_AGEMA_signal_21459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C ( clk ), .D ( new_AGEMA_signal_21466 ), .Q ( new_AGEMA_signal_21467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C ( clk ), .D ( new_AGEMA_signal_21474 ), .Q ( new_AGEMA_signal_21475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C ( clk ), .D ( new_AGEMA_signal_21482 ), .Q ( new_AGEMA_signal_21483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C ( clk ), .D ( new_AGEMA_signal_21490 ), .Q ( new_AGEMA_signal_21491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C ( clk ), .D ( new_AGEMA_signal_21498 ), .Q ( new_AGEMA_signal_21499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C ( clk ), .D ( new_AGEMA_signal_21512 ), .Q ( new_AGEMA_signal_21513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C ( clk ), .D ( new_AGEMA_signal_21516 ), .Q ( new_AGEMA_signal_21517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C ( clk ), .D ( new_AGEMA_signal_21520 ), .Q ( new_AGEMA_signal_21521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C ( clk ), .D ( new_AGEMA_signal_21524 ), .Q ( new_AGEMA_signal_21525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C ( clk ), .D ( new_AGEMA_signal_21528 ), .Q ( new_AGEMA_signal_21529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C ( clk ), .D ( new_AGEMA_signal_21544 ), .Q ( new_AGEMA_signal_21545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C ( clk ), .D ( new_AGEMA_signal_21550 ), .Q ( new_AGEMA_signal_21551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C ( clk ), .D ( new_AGEMA_signal_21556 ), .Q ( new_AGEMA_signal_21557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C ( clk ), .D ( new_AGEMA_signal_21562 ), .Q ( new_AGEMA_signal_21563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C ( clk ), .D ( new_AGEMA_signal_21568 ), .Q ( new_AGEMA_signal_21569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C ( clk ), .D ( new_AGEMA_signal_21584 ), .Q ( new_AGEMA_signal_21585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C ( clk ), .D ( new_AGEMA_signal_21592 ), .Q ( new_AGEMA_signal_21593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C ( clk ), .D ( new_AGEMA_signal_21600 ), .Q ( new_AGEMA_signal_21601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C ( clk ), .D ( new_AGEMA_signal_21608 ), .Q ( new_AGEMA_signal_21609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C ( clk ), .D ( new_AGEMA_signal_21616 ), .Q ( new_AGEMA_signal_21617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C ( clk ), .D ( new_AGEMA_signal_21654 ), .Q ( new_AGEMA_signal_21655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C ( clk ), .D ( new_AGEMA_signal_21662 ), .Q ( new_AGEMA_signal_21663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C ( clk ), .D ( new_AGEMA_signal_21670 ), .Q ( new_AGEMA_signal_21671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C ( clk ), .D ( new_AGEMA_signal_21678 ), .Q ( new_AGEMA_signal_21679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C ( clk ), .D ( new_AGEMA_signal_21686 ), .Q ( new_AGEMA_signal_21687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C ( clk ), .D ( new_AGEMA_signal_21702 ), .Q ( new_AGEMA_signal_21703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C ( clk ), .D ( new_AGEMA_signal_21708 ), .Q ( new_AGEMA_signal_21709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C ( clk ), .D ( new_AGEMA_signal_21714 ), .Q ( new_AGEMA_signal_21715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C ( clk ), .D ( new_AGEMA_signal_21720 ), .Q ( new_AGEMA_signal_21721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C ( clk ), .D ( new_AGEMA_signal_21726 ), .Q ( new_AGEMA_signal_21727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C ( clk ), .D ( new_AGEMA_signal_21754 ), .Q ( new_AGEMA_signal_21755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C ( clk ), .D ( new_AGEMA_signal_21762 ), .Q ( new_AGEMA_signal_21763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C ( clk ), .D ( new_AGEMA_signal_21770 ), .Q ( new_AGEMA_signal_21771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C ( clk ), .D ( new_AGEMA_signal_21778 ), .Q ( new_AGEMA_signal_21779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C ( clk ), .D ( new_AGEMA_signal_21786 ), .Q ( new_AGEMA_signal_21787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C ( clk ), .D ( new_AGEMA_signal_21812 ), .Q ( new_AGEMA_signal_21813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C ( clk ), .D ( new_AGEMA_signal_21818 ), .Q ( new_AGEMA_signal_21819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C ( clk ), .D ( new_AGEMA_signal_21824 ), .Q ( new_AGEMA_signal_21825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C ( clk ), .D ( new_AGEMA_signal_21830 ), .Q ( new_AGEMA_signal_21831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C ( clk ), .D ( new_AGEMA_signal_21836 ), .Q ( new_AGEMA_signal_21837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C ( clk ), .D ( new_AGEMA_signal_21842 ), .Q ( new_AGEMA_signal_21843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C ( clk ), .D ( new_AGEMA_signal_21848 ), .Q ( new_AGEMA_signal_21849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C ( clk ), .D ( new_AGEMA_signal_21854 ), .Q ( new_AGEMA_signal_21855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C ( clk ), .D ( new_AGEMA_signal_21860 ), .Q ( new_AGEMA_signal_21861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C ( clk ), .D ( new_AGEMA_signal_21866 ), .Q ( new_AGEMA_signal_21867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C ( clk ), .D ( new_AGEMA_signal_21872 ), .Q ( new_AGEMA_signal_21873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C ( clk ), .D ( new_AGEMA_signal_21878 ), .Q ( new_AGEMA_signal_21879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C ( clk ), .D ( new_AGEMA_signal_21884 ), .Q ( new_AGEMA_signal_21885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C ( clk ), .D ( new_AGEMA_signal_21890 ), .Q ( new_AGEMA_signal_21891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C ( clk ), .D ( new_AGEMA_signal_21896 ), .Q ( new_AGEMA_signal_21897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C ( clk ), .D ( new_AGEMA_signal_21902 ), .Q ( new_AGEMA_signal_21903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C ( clk ), .D ( new_AGEMA_signal_21908 ), .Q ( new_AGEMA_signal_21909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C ( clk ), .D ( new_AGEMA_signal_21914 ), .Q ( new_AGEMA_signal_21915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C ( clk ), .D ( new_AGEMA_signal_21920 ), .Q ( new_AGEMA_signal_21921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C ( clk ), .D ( new_AGEMA_signal_21926 ), .Q ( new_AGEMA_signal_21927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C ( clk ), .D ( new_AGEMA_signal_21932 ), .Q ( new_AGEMA_signal_21933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C ( clk ), .D ( new_AGEMA_signal_21938 ), .Q ( new_AGEMA_signal_21939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C ( clk ), .D ( new_AGEMA_signal_21944 ), .Q ( new_AGEMA_signal_21945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C ( clk ), .D ( new_AGEMA_signal_21950 ), .Q ( new_AGEMA_signal_21951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C ( clk ), .D ( new_AGEMA_signal_21956 ), .Q ( new_AGEMA_signal_21957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C ( clk ), .D ( new_AGEMA_signal_21984 ), .Q ( new_AGEMA_signal_21985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C ( clk ), .D ( new_AGEMA_signal_21992 ), .Q ( new_AGEMA_signal_21993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C ( clk ), .D ( new_AGEMA_signal_22000 ), .Q ( new_AGEMA_signal_22001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C ( clk ), .D ( new_AGEMA_signal_22008 ), .Q ( new_AGEMA_signal_22009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C ( clk ), .D ( new_AGEMA_signal_22016 ), .Q ( new_AGEMA_signal_22017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C ( clk ), .D ( new_AGEMA_signal_22042 ), .Q ( new_AGEMA_signal_22043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C ( clk ), .D ( new_AGEMA_signal_22048 ), .Q ( new_AGEMA_signal_22049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C ( clk ), .D ( new_AGEMA_signal_22054 ), .Q ( new_AGEMA_signal_22055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C ( clk ), .D ( new_AGEMA_signal_22060 ), .Q ( new_AGEMA_signal_22061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C ( clk ), .D ( new_AGEMA_signal_22066 ), .Q ( new_AGEMA_signal_22067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C ( clk ), .D ( new_AGEMA_signal_22074 ), .Q ( new_AGEMA_signal_22075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C ( clk ), .D ( new_AGEMA_signal_22082 ), .Q ( new_AGEMA_signal_22083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C ( clk ), .D ( new_AGEMA_signal_22090 ), .Q ( new_AGEMA_signal_22091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C ( clk ), .D ( new_AGEMA_signal_22098 ), .Q ( new_AGEMA_signal_22099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C ( clk ), .D ( new_AGEMA_signal_22106 ), .Q ( new_AGEMA_signal_22107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C ( clk ), .D ( new_AGEMA_signal_22122 ), .Q ( new_AGEMA_signal_22123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C ( clk ), .D ( new_AGEMA_signal_22128 ), .Q ( new_AGEMA_signal_22129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C ( clk ), .D ( new_AGEMA_signal_22134 ), .Q ( new_AGEMA_signal_22135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C ( clk ), .D ( new_AGEMA_signal_22140 ), .Q ( new_AGEMA_signal_22141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C ( clk ), .D ( new_AGEMA_signal_22146 ), .Q ( new_AGEMA_signal_22147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C ( clk ), .D ( new_AGEMA_signal_22172 ), .Q ( new_AGEMA_signal_22173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C ( clk ), .D ( new_AGEMA_signal_22178 ), .Q ( new_AGEMA_signal_22179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C ( clk ), .D ( new_AGEMA_signal_22184 ), .Q ( new_AGEMA_signal_22185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C ( clk ), .D ( new_AGEMA_signal_22190 ), .Q ( new_AGEMA_signal_22191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C ( clk ), .D ( new_AGEMA_signal_22196 ), .Q ( new_AGEMA_signal_22197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C ( clk ), .D ( new_AGEMA_signal_22202 ), .Q ( new_AGEMA_signal_22203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C ( clk ), .D ( new_AGEMA_signal_22208 ), .Q ( new_AGEMA_signal_22209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C ( clk ), .D ( new_AGEMA_signal_22214 ), .Q ( new_AGEMA_signal_22215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C ( clk ), .D ( new_AGEMA_signal_22220 ), .Q ( new_AGEMA_signal_22221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C ( clk ), .D ( new_AGEMA_signal_22226 ), .Q ( new_AGEMA_signal_22227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C ( clk ), .D ( new_AGEMA_signal_22234 ), .Q ( new_AGEMA_signal_22235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C ( clk ), .D ( new_AGEMA_signal_22242 ), .Q ( new_AGEMA_signal_22243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C ( clk ), .D ( new_AGEMA_signal_22250 ), .Q ( new_AGEMA_signal_22251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C ( clk ), .D ( new_AGEMA_signal_22258 ), .Q ( new_AGEMA_signal_22259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C ( clk ), .D ( new_AGEMA_signal_22266 ), .Q ( new_AGEMA_signal_22267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C ( clk ), .D ( new_AGEMA_signal_22274 ), .Q ( new_AGEMA_signal_22275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C ( clk ), .D ( new_AGEMA_signal_22282 ), .Q ( new_AGEMA_signal_22283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C ( clk ), .D ( new_AGEMA_signal_22290 ), .Q ( new_AGEMA_signal_22291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C ( clk ), .D ( new_AGEMA_signal_22298 ), .Q ( new_AGEMA_signal_22299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C ( clk ), .D ( new_AGEMA_signal_22306 ), .Q ( new_AGEMA_signal_22307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C ( clk ), .D ( new_AGEMA_signal_22312 ), .Q ( new_AGEMA_signal_22313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C ( clk ), .D ( new_AGEMA_signal_22318 ), .Q ( new_AGEMA_signal_22319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C ( clk ), .D ( new_AGEMA_signal_22324 ), .Q ( new_AGEMA_signal_22325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C ( clk ), .D ( new_AGEMA_signal_22330 ), .Q ( new_AGEMA_signal_22331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C ( clk ), .D ( new_AGEMA_signal_22336 ), .Q ( new_AGEMA_signal_22337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C ( clk ), .D ( new_AGEMA_signal_22342 ), .Q ( new_AGEMA_signal_22343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C ( clk ), .D ( new_AGEMA_signal_22348 ), .Q ( new_AGEMA_signal_22349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C ( clk ), .D ( new_AGEMA_signal_22354 ), .Q ( new_AGEMA_signal_22355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C ( clk ), .D ( new_AGEMA_signal_22360 ), .Q ( new_AGEMA_signal_22361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C ( clk ), .D ( new_AGEMA_signal_22366 ), .Q ( new_AGEMA_signal_22367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C ( clk ), .D ( new_AGEMA_signal_22512 ), .Q ( new_AGEMA_signal_22513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C ( clk ), .D ( new_AGEMA_signal_22520 ), .Q ( new_AGEMA_signal_22521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C ( clk ), .D ( new_AGEMA_signal_22528 ), .Q ( new_AGEMA_signal_22529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C ( clk ), .D ( new_AGEMA_signal_22536 ), .Q ( new_AGEMA_signal_22537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C ( clk ), .D ( new_AGEMA_signal_22544 ), .Q ( new_AGEMA_signal_22545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C ( clk ), .D ( new_AGEMA_signal_22552 ), .Q ( new_AGEMA_signal_22553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C ( clk ), .D ( new_AGEMA_signal_22560 ), .Q ( new_AGEMA_signal_22561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C ( clk ), .D ( new_AGEMA_signal_22568 ), .Q ( new_AGEMA_signal_22569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C ( clk ), .D ( new_AGEMA_signal_22576 ), .Q ( new_AGEMA_signal_22577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C ( clk ), .D ( new_AGEMA_signal_22584 ), .Q ( new_AGEMA_signal_22585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C ( clk ), .D ( new_AGEMA_signal_22592 ), .Q ( new_AGEMA_signal_22593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C ( clk ), .D ( new_AGEMA_signal_22600 ), .Q ( new_AGEMA_signal_22601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C ( clk ), .D ( new_AGEMA_signal_22608 ), .Q ( new_AGEMA_signal_22609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C ( clk ), .D ( new_AGEMA_signal_22616 ), .Q ( new_AGEMA_signal_22617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C ( clk ), .D ( new_AGEMA_signal_22624 ), .Q ( new_AGEMA_signal_22625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C ( clk ), .D ( new_AGEMA_signal_22632 ), .Q ( new_AGEMA_signal_22633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C ( clk ), .D ( new_AGEMA_signal_22640 ), .Q ( new_AGEMA_signal_22641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C ( clk ), .D ( new_AGEMA_signal_22648 ), .Q ( new_AGEMA_signal_22649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C ( clk ), .D ( new_AGEMA_signal_22656 ), .Q ( new_AGEMA_signal_22657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C ( clk ), .D ( new_AGEMA_signal_22664 ), .Q ( new_AGEMA_signal_22665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C ( clk ), .D ( new_AGEMA_signal_22704 ), .Q ( new_AGEMA_signal_22705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C ( clk ), .D ( new_AGEMA_signal_22714 ), .Q ( new_AGEMA_signal_22715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C ( clk ), .D ( new_AGEMA_signal_22724 ), .Q ( new_AGEMA_signal_22725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C ( clk ), .D ( new_AGEMA_signal_22734 ), .Q ( new_AGEMA_signal_22735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C ( clk ), .D ( new_AGEMA_signal_22744 ), .Q ( new_AGEMA_signal_22745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C ( clk ), .D ( new_AGEMA_signal_22752 ), .Q ( new_AGEMA_signal_22753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C ( clk ), .D ( new_AGEMA_signal_22760 ), .Q ( new_AGEMA_signal_22761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C ( clk ), .D ( new_AGEMA_signal_22768 ), .Q ( new_AGEMA_signal_22769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C ( clk ), .D ( new_AGEMA_signal_22776 ), .Q ( new_AGEMA_signal_22777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C ( clk ), .D ( new_AGEMA_signal_22784 ), .Q ( new_AGEMA_signal_22785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C ( clk ), .D ( new_AGEMA_signal_22792 ), .Q ( new_AGEMA_signal_22793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C ( clk ), .D ( new_AGEMA_signal_22800 ), .Q ( new_AGEMA_signal_22801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C ( clk ), .D ( new_AGEMA_signal_22808 ), .Q ( new_AGEMA_signal_22809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C ( clk ), .D ( new_AGEMA_signal_22816 ), .Q ( new_AGEMA_signal_22817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C ( clk ), .D ( new_AGEMA_signal_22824 ), .Q ( new_AGEMA_signal_22825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C ( clk ), .D ( new_AGEMA_signal_22832 ), .Q ( new_AGEMA_signal_22833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C ( clk ), .D ( new_AGEMA_signal_22840 ), .Q ( new_AGEMA_signal_22841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C ( clk ), .D ( new_AGEMA_signal_22848 ), .Q ( new_AGEMA_signal_22849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C ( clk ), .D ( new_AGEMA_signal_22856 ), .Q ( new_AGEMA_signal_22857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C ( clk ), .D ( new_AGEMA_signal_22864 ), .Q ( new_AGEMA_signal_22865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C ( clk ), .D ( new_AGEMA_signal_22954 ), .Q ( new_AGEMA_signal_22955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C ( clk ), .D ( new_AGEMA_signal_22964 ), .Q ( new_AGEMA_signal_22965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C ( clk ), .D ( new_AGEMA_signal_22974 ), .Q ( new_AGEMA_signal_22975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C ( clk ), .D ( new_AGEMA_signal_22984 ), .Q ( new_AGEMA_signal_22985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C ( clk ), .D ( new_AGEMA_signal_22994 ), .Q ( new_AGEMA_signal_22995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C ( clk ), .D ( new_AGEMA_signal_23002 ), .Q ( new_AGEMA_signal_23003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C ( clk ), .D ( new_AGEMA_signal_23010 ), .Q ( new_AGEMA_signal_23011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C ( clk ), .D ( new_AGEMA_signal_23018 ), .Q ( new_AGEMA_signal_23019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C ( clk ), .D ( new_AGEMA_signal_23026 ), .Q ( new_AGEMA_signal_23027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C ( clk ), .D ( new_AGEMA_signal_23034 ), .Q ( new_AGEMA_signal_23035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C ( clk ), .D ( new_AGEMA_signal_23072 ), .Q ( new_AGEMA_signal_23073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C ( clk ), .D ( new_AGEMA_signal_23080 ), .Q ( new_AGEMA_signal_23081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C ( clk ), .D ( new_AGEMA_signal_23088 ), .Q ( new_AGEMA_signal_23089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C ( clk ), .D ( new_AGEMA_signal_23096 ), .Q ( new_AGEMA_signal_23097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C ( clk ), .D ( new_AGEMA_signal_23104 ), .Q ( new_AGEMA_signal_23105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C ( clk ), .D ( new_AGEMA_signal_23112 ), .Q ( new_AGEMA_signal_23113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C ( clk ), .D ( new_AGEMA_signal_23120 ), .Q ( new_AGEMA_signal_23121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C ( clk ), .D ( new_AGEMA_signal_23128 ), .Q ( new_AGEMA_signal_23129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C ( clk ), .D ( new_AGEMA_signal_23136 ), .Q ( new_AGEMA_signal_23137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C ( clk ), .D ( new_AGEMA_signal_23144 ), .Q ( new_AGEMA_signal_23145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C ( clk ), .D ( new_AGEMA_signal_23202 ), .Q ( new_AGEMA_signal_23203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C ( clk ), .D ( new_AGEMA_signal_23210 ), .Q ( new_AGEMA_signal_23211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C ( clk ), .D ( new_AGEMA_signal_23218 ), .Q ( new_AGEMA_signal_23219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C ( clk ), .D ( new_AGEMA_signal_23226 ), .Q ( new_AGEMA_signal_23227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C ( clk ), .D ( new_AGEMA_signal_23234 ), .Q ( new_AGEMA_signal_23235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C ( clk ), .D ( new_AGEMA_signal_23532 ), .Q ( new_AGEMA_signal_23533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C ( clk ), .D ( new_AGEMA_signal_23542 ), .Q ( new_AGEMA_signal_23543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C ( clk ), .D ( new_AGEMA_signal_23552 ), .Q ( new_AGEMA_signal_23553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C ( clk ), .D ( new_AGEMA_signal_23562 ), .Q ( new_AGEMA_signal_23563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C ( clk ), .D ( new_AGEMA_signal_23572 ), .Q ( new_AGEMA_signal_23573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7738 ( .C ( clk ), .D ( new_AGEMA_signal_24512 ), .Q ( new_AGEMA_signal_24513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7752 ( .C ( clk ), .D ( new_AGEMA_signal_24526 ), .Q ( new_AGEMA_signal_24527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7766 ( .C ( clk ), .D ( new_AGEMA_signal_24540 ), .Q ( new_AGEMA_signal_24541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7780 ( .C ( clk ), .D ( new_AGEMA_signal_24554 ), .Q ( new_AGEMA_signal_24555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7794 ( .C ( clk ), .D ( new_AGEMA_signal_24568 ), .Q ( new_AGEMA_signal_24569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7848 ( .C ( clk ), .D ( new_AGEMA_signal_24622 ), .Q ( new_AGEMA_signal_24623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7862 ( .C ( clk ), .D ( new_AGEMA_signal_24636 ), .Q ( new_AGEMA_signal_24637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7876 ( .C ( clk ), .D ( new_AGEMA_signal_24650 ), .Q ( new_AGEMA_signal_24651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7890 ( .C ( clk ), .D ( new_AGEMA_signal_24664 ), .Q ( new_AGEMA_signal_24665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7904 ( .C ( clk ), .D ( new_AGEMA_signal_24678 ), .Q ( new_AGEMA_signal_24679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8028 ( .C ( clk ), .D ( new_AGEMA_signal_24802 ), .Q ( new_AGEMA_signal_24803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8044 ( .C ( clk ), .D ( new_AGEMA_signal_24818 ), .Q ( new_AGEMA_signal_24819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8060 ( .C ( clk ), .D ( new_AGEMA_signal_24834 ), .Q ( new_AGEMA_signal_24835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8076 ( .C ( clk ), .D ( new_AGEMA_signal_24850 ), .Q ( new_AGEMA_signal_24851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8092 ( .C ( clk ), .D ( new_AGEMA_signal_24866 ), .Q ( new_AGEMA_signal_24867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8138 ( .C ( clk ), .D ( new_AGEMA_signal_24912 ), .Q ( new_AGEMA_signal_24913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8154 ( .C ( clk ), .D ( new_AGEMA_signal_24928 ), .Q ( new_AGEMA_signal_24929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8170 ( .C ( clk ), .D ( new_AGEMA_signal_24944 ), .Q ( new_AGEMA_signal_24945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8186 ( .C ( clk ), .D ( new_AGEMA_signal_24960 ), .Q ( new_AGEMA_signal_24961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8202 ( .C ( clk ), .D ( new_AGEMA_signal_24976 ), .Q ( new_AGEMA_signal_24977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8518 ( .C ( clk ), .D ( new_AGEMA_signal_25292 ), .Q ( new_AGEMA_signal_25293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8536 ( .C ( clk ), .D ( new_AGEMA_signal_25310 ), .Q ( new_AGEMA_signal_25311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8554 ( .C ( clk ), .D ( new_AGEMA_signal_25328 ), .Q ( new_AGEMA_signal_25329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8572 ( .C ( clk ), .D ( new_AGEMA_signal_25346 ), .Q ( new_AGEMA_signal_25347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8590 ( .C ( clk ), .D ( new_AGEMA_signal_25364 ), .Q ( new_AGEMA_signal_25365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8768 ( .C ( clk ), .D ( new_AGEMA_signal_25542 ), .Q ( new_AGEMA_signal_25543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8788 ( .C ( clk ), .D ( new_AGEMA_signal_25562 ), .Q ( new_AGEMA_signal_25563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8808 ( .C ( clk ), .D ( new_AGEMA_signal_25582 ), .Q ( new_AGEMA_signal_25583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8828 ( .C ( clk ), .D ( new_AGEMA_signal_25602 ), .Q ( new_AGEMA_signal_25603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8848 ( .C ( clk ), .D ( new_AGEMA_signal_25622 ), .Q ( new_AGEMA_signal_25623 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_3639 ( .C ( clk ), .D ( new_AGEMA_signal_20413 ), .Q ( new_AGEMA_signal_20414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C ( clk ), .D ( new_AGEMA_signal_20417 ), .Q ( new_AGEMA_signal_20418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C ( clk ), .D ( new_AGEMA_signal_20421 ), .Q ( new_AGEMA_signal_20422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C ( clk ), .D ( new_AGEMA_signal_20425 ), .Q ( new_AGEMA_signal_20426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C ( clk ), .D ( new_AGEMA_signal_20429 ), .Q ( new_AGEMA_signal_20430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C ( clk ), .D ( new_AGEMA_signal_20433 ), .Q ( new_AGEMA_signal_20434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C ( clk ), .D ( new_AGEMA_signal_20437 ), .Q ( new_AGEMA_signal_20438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C ( clk ), .D ( new_AGEMA_signal_20441 ), .Q ( new_AGEMA_signal_20442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C ( clk ), .D ( new_AGEMA_signal_20445 ), .Q ( new_AGEMA_signal_20446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C ( clk ), .D ( new_AGEMA_signal_20449 ), .Q ( new_AGEMA_signal_20450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C ( clk ), .D ( new_AGEMA_signal_20457 ), .Q ( new_AGEMA_signal_20458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C ( clk ), .D ( new_AGEMA_signal_20465 ), .Q ( new_AGEMA_signal_20466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C ( clk ), .D ( new_AGEMA_signal_20473 ), .Q ( new_AGEMA_signal_20474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C ( clk ), .D ( new_AGEMA_signal_20481 ), .Q ( new_AGEMA_signal_20482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C ( clk ), .D ( new_AGEMA_signal_20489 ), .Q ( new_AGEMA_signal_20490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_20492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C ( clk ), .D ( new_AGEMA_signal_3102 ), .Q ( new_AGEMA_signal_20494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C ( clk ), .D ( new_AGEMA_signal_3103 ), .Q ( new_AGEMA_signal_20496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C ( clk ), .D ( new_AGEMA_signal_3104 ), .Q ( new_AGEMA_signal_20498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C ( clk ), .D ( new_AGEMA_signal_3105 ), .Q ( new_AGEMA_signal_20500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C ( clk ), .D ( new_AGEMA_signal_20507 ), .Q ( new_AGEMA_signal_20508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C ( clk ), .D ( new_AGEMA_signal_20515 ), .Q ( new_AGEMA_signal_20516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C ( clk ), .D ( new_AGEMA_signal_20523 ), .Q ( new_AGEMA_signal_20524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C ( clk ), .D ( new_AGEMA_signal_20531 ), .Q ( new_AGEMA_signal_20532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C ( clk ), .D ( new_AGEMA_signal_20539 ), .Q ( new_AGEMA_signal_20540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C ( clk ), .D ( new_AGEMA_signal_20545 ), .Q ( new_AGEMA_signal_20546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C ( clk ), .D ( new_AGEMA_signal_20551 ), .Q ( new_AGEMA_signal_20552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C ( clk ), .D ( new_AGEMA_signal_20557 ), .Q ( new_AGEMA_signal_20558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C ( clk ), .D ( new_AGEMA_signal_20563 ), .Q ( new_AGEMA_signal_20564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C ( clk ), .D ( new_AGEMA_signal_20569 ), .Q ( new_AGEMA_signal_20570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C ( clk ), .D ( new_AGEMA_signal_20573 ), .Q ( new_AGEMA_signal_20574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C ( clk ), .D ( new_AGEMA_signal_20577 ), .Q ( new_AGEMA_signal_20578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C ( clk ), .D ( new_AGEMA_signal_20581 ), .Q ( new_AGEMA_signal_20582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C ( clk ), .D ( new_AGEMA_signal_20585 ), .Q ( new_AGEMA_signal_20586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C ( clk ), .D ( new_AGEMA_signal_20589 ), .Q ( new_AGEMA_signal_20590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C ( clk ), .D ( new_AGEMA_signal_20595 ), .Q ( new_AGEMA_signal_20596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C ( clk ), .D ( new_AGEMA_signal_20601 ), .Q ( new_AGEMA_signal_20602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C ( clk ), .D ( new_AGEMA_signal_20607 ), .Q ( new_AGEMA_signal_20608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C ( clk ), .D ( new_AGEMA_signal_20613 ), .Q ( new_AGEMA_signal_20614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C ( clk ), .D ( new_AGEMA_signal_20619 ), .Q ( new_AGEMA_signal_20620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C ( clk ), .D ( new_AGEMA_signal_20135 ), .Q ( new_AGEMA_signal_20622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C ( clk ), .D ( new_AGEMA_signal_20139 ), .Q ( new_AGEMA_signal_20624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C ( clk ), .D ( new_AGEMA_signal_20143 ), .Q ( new_AGEMA_signal_20626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C ( clk ), .D ( new_AGEMA_signal_20147 ), .Q ( new_AGEMA_signal_20628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C ( clk ), .D ( new_AGEMA_signal_20151 ), .Q ( new_AGEMA_signal_20630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C ( clk ), .D ( new_AGEMA_signal_20635 ), .Q ( new_AGEMA_signal_20636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C ( clk ), .D ( new_AGEMA_signal_20641 ), .Q ( new_AGEMA_signal_20642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C ( clk ), .D ( new_AGEMA_signal_20647 ), .Q ( new_AGEMA_signal_20648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C ( clk ), .D ( new_AGEMA_signal_20653 ), .Q ( new_AGEMA_signal_20654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C ( clk ), .D ( new_AGEMA_signal_20659 ), .Q ( new_AGEMA_signal_20660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C ( clk ), .D ( new_AGEMA_signal_20665 ), .Q ( new_AGEMA_signal_20666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C ( clk ), .D ( new_AGEMA_signal_20671 ), .Q ( new_AGEMA_signal_20672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C ( clk ), .D ( new_AGEMA_signal_20677 ), .Q ( new_AGEMA_signal_20678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C ( clk ), .D ( new_AGEMA_signal_20683 ), .Q ( new_AGEMA_signal_20684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C ( clk ), .D ( new_AGEMA_signal_20689 ), .Q ( new_AGEMA_signal_20690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_20692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C ( clk ), .D ( new_AGEMA_signal_3174 ), .Q ( new_AGEMA_signal_20694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C ( clk ), .D ( new_AGEMA_signal_3175 ), .Q ( new_AGEMA_signal_20696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C ( clk ), .D ( new_AGEMA_signal_3176 ), .Q ( new_AGEMA_signal_20698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C ( clk ), .D ( new_AGEMA_signal_3177 ), .Q ( new_AGEMA_signal_20700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C ( clk ), .D ( new_AGEMA_signal_20703 ), .Q ( new_AGEMA_signal_20704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C ( clk ), .D ( new_AGEMA_signal_20707 ), .Q ( new_AGEMA_signal_20708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C ( clk ), .D ( new_AGEMA_signal_20711 ), .Q ( new_AGEMA_signal_20712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C ( clk ), .D ( new_AGEMA_signal_20715 ), .Q ( new_AGEMA_signal_20716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C ( clk ), .D ( new_AGEMA_signal_20719 ), .Q ( new_AGEMA_signal_20720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C ( clk ), .D ( new_AGEMA_signal_20725 ), .Q ( new_AGEMA_signal_20726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C ( clk ), .D ( new_AGEMA_signal_20731 ), .Q ( new_AGEMA_signal_20732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C ( clk ), .D ( new_AGEMA_signal_20737 ), .Q ( new_AGEMA_signal_20738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C ( clk ), .D ( new_AGEMA_signal_20743 ), .Q ( new_AGEMA_signal_20744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C ( clk ), .D ( new_AGEMA_signal_20749 ), .Q ( new_AGEMA_signal_20750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C ( clk ), .D ( new_AGEMA_signal_20755 ), .Q ( new_AGEMA_signal_20756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C ( clk ), .D ( new_AGEMA_signal_20761 ), .Q ( new_AGEMA_signal_20762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C ( clk ), .D ( new_AGEMA_signal_20767 ), .Q ( new_AGEMA_signal_20768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C ( clk ), .D ( new_AGEMA_signal_20773 ), .Q ( new_AGEMA_signal_20774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C ( clk ), .D ( new_AGEMA_signal_20779 ), .Q ( new_AGEMA_signal_20780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_20782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C ( clk ), .D ( new_AGEMA_signal_3198 ), .Q ( new_AGEMA_signal_20784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C ( clk ), .D ( new_AGEMA_signal_3199 ), .Q ( new_AGEMA_signal_20786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C ( clk ), .D ( new_AGEMA_signal_3200 ), .Q ( new_AGEMA_signal_20788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C ( clk ), .D ( new_AGEMA_signal_3201 ), .Q ( new_AGEMA_signal_20790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C ( clk ), .D ( new_AGEMA_signal_20795 ), .Q ( new_AGEMA_signal_20796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C ( clk ), .D ( new_AGEMA_signal_20801 ), .Q ( new_AGEMA_signal_20802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C ( clk ), .D ( new_AGEMA_signal_20807 ), .Q ( new_AGEMA_signal_20808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C ( clk ), .D ( new_AGEMA_signal_20813 ), .Q ( new_AGEMA_signal_20814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C ( clk ), .D ( new_AGEMA_signal_20819 ), .Q ( new_AGEMA_signal_20820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_20822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C ( clk ), .D ( new_AGEMA_signal_3214 ), .Q ( new_AGEMA_signal_20824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C ( clk ), .D ( new_AGEMA_signal_3215 ), .Q ( new_AGEMA_signal_20826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C ( clk ), .D ( new_AGEMA_signal_3216 ), .Q ( new_AGEMA_signal_20828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C ( clk ), .D ( new_AGEMA_signal_3217 ), .Q ( new_AGEMA_signal_20830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C ( clk ), .D ( new_AGEMA_signal_20833 ), .Q ( new_AGEMA_signal_20834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C ( clk ), .D ( new_AGEMA_signal_20837 ), .Q ( new_AGEMA_signal_20838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C ( clk ), .D ( new_AGEMA_signal_20841 ), .Q ( new_AGEMA_signal_20842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C ( clk ), .D ( new_AGEMA_signal_20845 ), .Q ( new_AGEMA_signal_20846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C ( clk ), .D ( new_AGEMA_signal_20849 ), .Q ( new_AGEMA_signal_20850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C ( clk ), .D ( new_AGEMA_signal_20853 ), .Q ( new_AGEMA_signal_20854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C ( clk ), .D ( new_AGEMA_signal_20857 ), .Q ( new_AGEMA_signal_20858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C ( clk ), .D ( new_AGEMA_signal_20861 ), .Q ( new_AGEMA_signal_20862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C ( clk ), .D ( new_AGEMA_signal_20865 ), .Q ( new_AGEMA_signal_20866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C ( clk ), .D ( new_AGEMA_signal_20869 ), .Q ( new_AGEMA_signal_20870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C ( clk ), .D ( new_AGEMA_signal_20103 ), .Q ( new_AGEMA_signal_20872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C ( clk ), .D ( new_AGEMA_signal_20105 ), .Q ( new_AGEMA_signal_20874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C ( clk ), .D ( new_AGEMA_signal_20107 ), .Q ( new_AGEMA_signal_20876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C ( clk ), .D ( new_AGEMA_signal_20109 ), .Q ( new_AGEMA_signal_20878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C ( clk ), .D ( new_AGEMA_signal_20111 ), .Q ( new_AGEMA_signal_20880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C ( clk ), .D ( new_AGEMA_signal_20887 ), .Q ( new_AGEMA_signal_20888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C ( clk ), .D ( new_AGEMA_signal_20895 ), .Q ( new_AGEMA_signal_20896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C ( clk ), .D ( new_AGEMA_signal_20903 ), .Q ( new_AGEMA_signal_20904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C ( clk ), .D ( new_AGEMA_signal_20911 ), .Q ( new_AGEMA_signal_20912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C ( clk ), .D ( new_AGEMA_signal_20919 ), .Q ( new_AGEMA_signal_20920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C ( clk ), .D ( new_AGEMA_signal_20925 ), .Q ( new_AGEMA_signal_20926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C ( clk ), .D ( new_AGEMA_signal_20931 ), .Q ( new_AGEMA_signal_20932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C ( clk ), .D ( new_AGEMA_signal_20937 ), .Q ( new_AGEMA_signal_20938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C ( clk ), .D ( new_AGEMA_signal_20943 ), .Q ( new_AGEMA_signal_20944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C ( clk ), .D ( new_AGEMA_signal_20949 ), .Q ( new_AGEMA_signal_20950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C ( clk ), .D ( new_AGEMA_signal_20953 ), .Q ( new_AGEMA_signal_20954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C ( clk ), .D ( new_AGEMA_signal_20957 ), .Q ( new_AGEMA_signal_20958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C ( clk ), .D ( new_AGEMA_signal_20961 ), .Q ( new_AGEMA_signal_20962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C ( clk ), .D ( new_AGEMA_signal_20965 ), .Q ( new_AGEMA_signal_20966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C ( clk ), .D ( new_AGEMA_signal_20969 ), .Q ( new_AGEMA_signal_20970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C ( clk ), .D ( new_AGEMA_signal_20973 ), .Q ( new_AGEMA_signal_20974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C ( clk ), .D ( new_AGEMA_signal_20977 ), .Q ( new_AGEMA_signal_20978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C ( clk ), .D ( new_AGEMA_signal_20981 ), .Q ( new_AGEMA_signal_20982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C ( clk ), .D ( new_AGEMA_signal_20985 ), .Q ( new_AGEMA_signal_20986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C ( clk ), .D ( new_AGEMA_signal_20989 ), .Q ( new_AGEMA_signal_20990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_20992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C ( clk ), .D ( new_AGEMA_signal_2718 ), .Q ( new_AGEMA_signal_20994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C ( clk ), .D ( new_AGEMA_signal_2719 ), .Q ( new_AGEMA_signal_20996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C ( clk ), .D ( new_AGEMA_signal_2720 ), .Q ( new_AGEMA_signal_20998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C ( clk ), .D ( new_AGEMA_signal_2721 ), .Q ( new_AGEMA_signal_21000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_21002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C ( clk ), .D ( new_AGEMA_signal_3286 ), .Q ( new_AGEMA_signal_21004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C ( clk ), .D ( new_AGEMA_signal_3287 ), .Q ( new_AGEMA_signal_21006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C ( clk ), .D ( new_AGEMA_signal_3288 ), .Q ( new_AGEMA_signal_21008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C ( clk ), .D ( new_AGEMA_signal_3289 ), .Q ( new_AGEMA_signal_21010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C ( clk ), .D ( new_AGEMA_signal_21013 ), .Q ( new_AGEMA_signal_21014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C ( clk ), .D ( new_AGEMA_signal_21017 ), .Q ( new_AGEMA_signal_21018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C ( clk ), .D ( new_AGEMA_signal_21021 ), .Q ( new_AGEMA_signal_21022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C ( clk ), .D ( new_AGEMA_signal_21025 ), .Q ( new_AGEMA_signal_21026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C ( clk ), .D ( new_AGEMA_signal_21029 ), .Q ( new_AGEMA_signal_21030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C ( clk ), .D ( new_AGEMA_signal_21033 ), .Q ( new_AGEMA_signal_21034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C ( clk ), .D ( new_AGEMA_signal_21037 ), .Q ( new_AGEMA_signal_21038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C ( clk ), .D ( new_AGEMA_signal_21041 ), .Q ( new_AGEMA_signal_21042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C ( clk ), .D ( new_AGEMA_signal_21045 ), .Q ( new_AGEMA_signal_21046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C ( clk ), .D ( new_AGEMA_signal_21049 ), .Q ( new_AGEMA_signal_21050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_21052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C ( clk ), .D ( new_AGEMA_signal_2762 ), .Q ( new_AGEMA_signal_21054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C ( clk ), .D ( new_AGEMA_signal_2763 ), .Q ( new_AGEMA_signal_21056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C ( clk ), .D ( new_AGEMA_signal_2764 ), .Q ( new_AGEMA_signal_21058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C ( clk ), .D ( new_AGEMA_signal_2765 ), .Q ( new_AGEMA_signal_21060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C ( clk ), .D ( new_AGEMA_signal_21065 ), .Q ( new_AGEMA_signal_21066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C ( clk ), .D ( new_AGEMA_signal_21071 ), .Q ( new_AGEMA_signal_21072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C ( clk ), .D ( new_AGEMA_signal_21077 ), .Q ( new_AGEMA_signal_21078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C ( clk ), .D ( new_AGEMA_signal_21083 ), .Q ( new_AGEMA_signal_21084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C ( clk ), .D ( new_AGEMA_signal_21089 ), .Q ( new_AGEMA_signal_21090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C ( clk ), .D ( new_AGEMA_signal_21093 ), .Q ( new_AGEMA_signal_21094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C ( clk ), .D ( new_AGEMA_signal_21097 ), .Q ( new_AGEMA_signal_21098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C ( clk ), .D ( new_AGEMA_signal_21101 ), .Q ( new_AGEMA_signal_21102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C ( clk ), .D ( new_AGEMA_signal_21105 ), .Q ( new_AGEMA_signal_21106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C ( clk ), .D ( new_AGEMA_signal_21109 ), .Q ( new_AGEMA_signal_21110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C ( clk ), .D ( new_AGEMA_signal_20123 ), .Q ( new_AGEMA_signal_21112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C ( clk ), .D ( new_AGEMA_signal_20125 ), .Q ( new_AGEMA_signal_21114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C ( clk ), .D ( new_AGEMA_signal_20127 ), .Q ( new_AGEMA_signal_21116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C ( clk ), .D ( new_AGEMA_signal_20129 ), .Q ( new_AGEMA_signal_21118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C ( clk ), .D ( new_AGEMA_signal_20131 ), .Q ( new_AGEMA_signal_21120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C ( clk ), .D ( new_AGEMA_signal_21123 ), .Q ( new_AGEMA_signal_21124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C ( clk ), .D ( new_AGEMA_signal_21127 ), .Q ( new_AGEMA_signal_21128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C ( clk ), .D ( new_AGEMA_signal_21131 ), .Q ( new_AGEMA_signal_21132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C ( clk ), .D ( new_AGEMA_signal_21135 ), .Q ( new_AGEMA_signal_21136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C ( clk ), .D ( new_AGEMA_signal_21139 ), .Q ( new_AGEMA_signal_21140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C ( clk ), .D ( new_AGEMA_signal_21143 ), .Q ( new_AGEMA_signal_21144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C ( clk ), .D ( new_AGEMA_signal_21147 ), .Q ( new_AGEMA_signal_21148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C ( clk ), .D ( new_AGEMA_signal_21151 ), .Q ( new_AGEMA_signal_21152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C ( clk ), .D ( new_AGEMA_signal_21155 ), .Q ( new_AGEMA_signal_21156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C ( clk ), .D ( new_AGEMA_signal_21159 ), .Q ( new_AGEMA_signal_21160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C ( clk ), .D ( new_AGEMA_signal_21163 ), .Q ( new_AGEMA_signal_21164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C ( clk ), .D ( new_AGEMA_signal_21167 ), .Q ( new_AGEMA_signal_21168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C ( clk ), .D ( new_AGEMA_signal_21171 ), .Q ( new_AGEMA_signal_21172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C ( clk ), .D ( new_AGEMA_signal_21175 ), .Q ( new_AGEMA_signal_21176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C ( clk ), .D ( new_AGEMA_signal_21179 ), .Q ( new_AGEMA_signal_21180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_21182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C ( clk ), .D ( new_AGEMA_signal_2838 ), .Q ( new_AGEMA_signal_21184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C ( clk ), .D ( new_AGEMA_signal_2839 ), .Q ( new_AGEMA_signal_21186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C ( clk ), .D ( new_AGEMA_signal_2840 ), .Q ( new_AGEMA_signal_21188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C ( clk ), .D ( new_AGEMA_signal_2841 ), .Q ( new_AGEMA_signal_21190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C ( clk ), .D ( new_AGEMA_signal_21193 ), .Q ( new_AGEMA_signal_21194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C ( clk ), .D ( new_AGEMA_signal_21197 ), .Q ( new_AGEMA_signal_21198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C ( clk ), .D ( new_AGEMA_signal_21201 ), .Q ( new_AGEMA_signal_21202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C ( clk ), .D ( new_AGEMA_signal_21205 ), .Q ( new_AGEMA_signal_21206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C ( clk ), .D ( new_AGEMA_signal_21209 ), .Q ( new_AGEMA_signal_21210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C ( clk ), .D ( new_AGEMA_signal_19933 ), .Q ( new_AGEMA_signal_21212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C ( clk ), .D ( new_AGEMA_signal_19935 ), .Q ( new_AGEMA_signal_21214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C ( clk ), .D ( new_AGEMA_signal_19937 ), .Q ( new_AGEMA_signal_21216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C ( clk ), .D ( new_AGEMA_signal_19939 ), .Q ( new_AGEMA_signal_21218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C ( clk ), .D ( new_AGEMA_signal_19941 ), .Q ( new_AGEMA_signal_21220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C ( clk ), .D ( new_AGEMA_signal_21225 ), .Q ( new_AGEMA_signal_21226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C ( clk ), .D ( new_AGEMA_signal_21231 ), .Q ( new_AGEMA_signal_21232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C ( clk ), .D ( new_AGEMA_signal_21237 ), .Q ( new_AGEMA_signal_21238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C ( clk ), .D ( new_AGEMA_signal_21243 ), .Q ( new_AGEMA_signal_21244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C ( clk ), .D ( new_AGEMA_signal_21249 ), .Q ( new_AGEMA_signal_21250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C ( clk ), .D ( new_AGEMA_signal_21255 ), .Q ( new_AGEMA_signal_21256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C ( clk ), .D ( new_AGEMA_signal_21261 ), .Q ( new_AGEMA_signal_21262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C ( clk ), .D ( new_AGEMA_signal_21267 ), .Q ( new_AGEMA_signal_21268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C ( clk ), .D ( new_AGEMA_signal_21273 ), .Q ( new_AGEMA_signal_21274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C ( clk ), .D ( new_AGEMA_signal_21279 ), .Q ( new_AGEMA_signal_21280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C ( clk ), .D ( new_AGEMA_signal_21283 ), .Q ( new_AGEMA_signal_21284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C ( clk ), .D ( new_AGEMA_signal_21287 ), .Q ( new_AGEMA_signal_21288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C ( clk ), .D ( new_AGEMA_signal_21291 ), .Q ( new_AGEMA_signal_21292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C ( clk ), .D ( new_AGEMA_signal_21295 ), .Q ( new_AGEMA_signal_21296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C ( clk ), .D ( new_AGEMA_signal_21299 ), .Q ( new_AGEMA_signal_21300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C ( clk ), .D ( new_AGEMA_signal_19877 ), .Q ( new_AGEMA_signal_21302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C ( clk ), .D ( new_AGEMA_signal_19883 ), .Q ( new_AGEMA_signal_21304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C ( clk ), .D ( new_AGEMA_signal_19889 ), .Q ( new_AGEMA_signal_21306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C ( clk ), .D ( new_AGEMA_signal_19895 ), .Q ( new_AGEMA_signal_21308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C ( clk ), .D ( new_AGEMA_signal_19901 ), .Q ( new_AGEMA_signal_21310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C ( clk ), .D ( new_AGEMA_signal_21317 ), .Q ( new_AGEMA_signal_21318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C ( clk ), .D ( new_AGEMA_signal_21325 ), .Q ( new_AGEMA_signal_21326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C ( clk ), .D ( new_AGEMA_signal_21333 ), .Q ( new_AGEMA_signal_21334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C ( clk ), .D ( new_AGEMA_signal_21341 ), .Q ( new_AGEMA_signal_21342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C ( clk ), .D ( new_AGEMA_signal_21349 ), .Q ( new_AGEMA_signal_21350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_21352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C ( clk ), .D ( new_AGEMA_signal_2910 ), .Q ( new_AGEMA_signal_21354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C ( clk ), .D ( new_AGEMA_signal_2911 ), .Q ( new_AGEMA_signal_21356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C ( clk ), .D ( new_AGEMA_signal_2912 ), .Q ( new_AGEMA_signal_21358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C ( clk ), .D ( new_AGEMA_signal_2913 ), .Q ( new_AGEMA_signal_21360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C ( clk ), .D ( new_AGEMA_signal_21363 ), .Q ( new_AGEMA_signal_21364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C ( clk ), .D ( new_AGEMA_signal_21367 ), .Q ( new_AGEMA_signal_21368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C ( clk ), .D ( new_AGEMA_signal_21371 ), .Q ( new_AGEMA_signal_21372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C ( clk ), .D ( new_AGEMA_signal_21375 ), .Q ( new_AGEMA_signal_21376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C ( clk ), .D ( new_AGEMA_signal_21379 ), .Q ( new_AGEMA_signal_21380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C ( clk ), .D ( new_AGEMA_signal_21383 ), .Q ( new_AGEMA_signal_21384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C ( clk ), .D ( new_AGEMA_signal_21387 ), .Q ( new_AGEMA_signal_21388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C ( clk ), .D ( new_AGEMA_signal_21391 ), .Q ( new_AGEMA_signal_21392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C ( clk ), .D ( new_AGEMA_signal_21395 ), .Q ( new_AGEMA_signal_21396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C ( clk ), .D ( new_AGEMA_signal_21399 ), .Q ( new_AGEMA_signal_21400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C ( clk ), .D ( new_AGEMA_signal_21403 ), .Q ( new_AGEMA_signal_21404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C ( clk ), .D ( new_AGEMA_signal_21407 ), .Q ( new_AGEMA_signal_21408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C ( clk ), .D ( new_AGEMA_signal_21411 ), .Q ( new_AGEMA_signal_21412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C ( clk ), .D ( new_AGEMA_signal_21415 ), .Q ( new_AGEMA_signal_21416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C ( clk ), .D ( new_AGEMA_signal_21419 ), .Q ( new_AGEMA_signal_21420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C ( clk ), .D ( new_AGEMA_signal_21423 ), .Q ( new_AGEMA_signal_21424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C ( clk ), .D ( new_AGEMA_signal_21427 ), .Q ( new_AGEMA_signal_21428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C ( clk ), .D ( new_AGEMA_signal_21431 ), .Q ( new_AGEMA_signal_21432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C ( clk ), .D ( new_AGEMA_signal_21435 ), .Q ( new_AGEMA_signal_21436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C ( clk ), .D ( new_AGEMA_signal_21439 ), .Q ( new_AGEMA_signal_21440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C ( clk ), .D ( new_AGEMA_signal_21443 ), .Q ( new_AGEMA_signal_21444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C ( clk ), .D ( new_AGEMA_signal_21447 ), .Q ( new_AGEMA_signal_21448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C ( clk ), .D ( new_AGEMA_signal_21451 ), .Q ( new_AGEMA_signal_21452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C ( clk ), .D ( new_AGEMA_signal_21455 ), .Q ( new_AGEMA_signal_21456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C ( clk ), .D ( new_AGEMA_signal_21459 ), .Q ( new_AGEMA_signal_21460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C ( clk ), .D ( new_AGEMA_signal_21467 ), .Q ( new_AGEMA_signal_21468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C ( clk ), .D ( new_AGEMA_signal_21475 ), .Q ( new_AGEMA_signal_21476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C ( clk ), .D ( new_AGEMA_signal_21483 ), .Q ( new_AGEMA_signal_21484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C ( clk ), .D ( new_AGEMA_signal_21491 ), .Q ( new_AGEMA_signal_21492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C ( clk ), .D ( new_AGEMA_signal_21499 ), .Q ( new_AGEMA_signal_21500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_21502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C ( clk ), .D ( new_AGEMA_signal_3490 ), .Q ( new_AGEMA_signal_21504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C ( clk ), .D ( new_AGEMA_signal_3491 ), .Q ( new_AGEMA_signal_21506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C ( clk ), .D ( new_AGEMA_signal_3492 ), .Q ( new_AGEMA_signal_21508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C ( clk ), .D ( new_AGEMA_signal_3493 ), .Q ( new_AGEMA_signal_21510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C ( clk ), .D ( new_AGEMA_signal_21513 ), .Q ( new_AGEMA_signal_21514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C ( clk ), .D ( new_AGEMA_signal_21517 ), .Q ( new_AGEMA_signal_21518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C ( clk ), .D ( new_AGEMA_signal_21521 ), .Q ( new_AGEMA_signal_21522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C ( clk ), .D ( new_AGEMA_signal_21525 ), .Q ( new_AGEMA_signal_21526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C ( clk ), .D ( new_AGEMA_signal_21529 ), .Q ( new_AGEMA_signal_21530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_21532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C ( clk ), .D ( new_AGEMA_signal_3506 ), .Q ( new_AGEMA_signal_21534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C ( clk ), .D ( new_AGEMA_signal_3507 ), .Q ( new_AGEMA_signal_21536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C ( clk ), .D ( new_AGEMA_signal_3508 ), .Q ( new_AGEMA_signal_21538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C ( clk ), .D ( new_AGEMA_signal_3509 ), .Q ( new_AGEMA_signal_21540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C ( clk ), .D ( new_AGEMA_signal_21545 ), .Q ( new_AGEMA_signal_21546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C ( clk ), .D ( new_AGEMA_signal_21551 ), .Q ( new_AGEMA_signal_21552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C ( clk ), .D ( new_AGEMA_signal_21557 ), .Q ( new_AGEMA_signal_21558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C ( clk ), .D ( new_AGEMA_signal_21563 ), .Q ( new_AGEMA_signal_21564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C ( clk ), .D ( new_AGEMA_signal_21569 ), .Q ( new_AGEMA_signal_21570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C ( clk ), .D ( new_AGEMA_signal_21585 ), .Q ( new_AGEMA_signal_21586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C ( clk ), .D ( new_AGEMA_signal_21593 ), .Q ( new_AGEMA_signal_21594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C ( clk ), .D ( new_AGEMA_signal_21601 ), .Q ( new_AGEMA_signal_21602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C ( clk ), .D ( new_AGEMA_signal_21609 ), .Q ( new_AGEMA_signal_21610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C ( clk ), .D ( new_AGEMA_signal_21617 ), .Q ( new_AGEMA_signal_21618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_21632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C ( clk ), .D ( new_AGEMA_signal_3122 ), .Q ( new_AGEMA_signal_21636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C ( clk ), .D ( new_AGEMA_signal_3123 ), .Q ( new_AGEMA_signal_21640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C ( clk ), .D ( new_AGEMA_signal_3124 ), .Q ( new_AGEMA_signal_21644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C ( clk ), .D ( new_AGEMA_signal_3125 ), .Q ( new_AGEMA_signal_21648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C ( clk ), .D ( new_AGEMA_signal_21655 ), .Q ( new_AGEMA_signal_21656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C ( clk ), .D ( new_AGEMA_signal_21663 ), .Q ( new_AGEMA_signal_21664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C ( clk ), .D ( new_AGEMA_signal_21671 ), .Q ( new_AGEMA_signal_21672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C ( clk ), .D ( new_AGEMA_signal_21679 ), .Q ( new_AGEMA_signal_21680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C ( clk ), .D ( new_AGEMA_signal_21687 ), .Q ( new_AGEMA_signal_21688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C ( clk ), .D ( new_AGEMA_signal_21703 ), .Q ( new_AGEMA_signal_21704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C ( clk ), .D ( new_AGEMA_signal_21709 ), .Q ( new_AGEMA_signal_21710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C ( clk ), .D ( new_AGEMA_signal_21715 ), .Q ( new_AGEMA_signal_21716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C ( clk ), .D ( new_AGEMA_signal_21721 ), .Q ( new_AGEMA_signal_21722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C ( clk ), .D ( new_AGEMA_signal_21727 ), .Q ( new_AGEMA_signal_21728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_21732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C ( clk ), .D ( new_AGEMA_signal_3158 ), .Q ( new_AGEMA_signal_21736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C ( clk ), .D ( new_AGEMA_signal_3159 ), .Q ( new_AGEMA_signal_21740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C ( clk ), .D ( new_AGEMA_signal_3160 ), .Q ( new_AGEMA_signal_21744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C ( clk ), .D ( new_AGEMA_signal_3161 ), .Q ( new_AGEMA_signal_21748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C ( clk ), .D ( new_AGEMA_signal_21755 ), .Q ( new_AGEMA_signal_21756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C ( clk ), .D ( new_AGEMA_signal_21763 ), .Q ( new_AGEMA_signal_21764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C ( clk ), .D ( new_AGEMA_signal_21771 ), .Q ( new_AGEMA_signal_21772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C ( clk ), .D ( new_AGEMA_signal_21779 ), .Q ( new_AGEMA_signal_21780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C ( clk ), .D ( new_AGEMA_signal_21787 ), .Q ( new_AGEMA_signal_21788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_21792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C ( clk ), .D ( new_AGEMA_signal_3206 ), .Q ( new_AGEMA_signal_21796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C ( clk ), .D ( new_AGEMA_signal_3207 ), .Q ( new_AGEMA_signal_21800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C ( clk ), .D ( new_AGEMA_signal_3208 ), .Q ( new_AGEMA_signal_21804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C ( clk ), .D ( new_AGEMA_signal_3209 ), .Q ( new_AGEMA_signal_21808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C ( clk ), .D ( new_AGEMA_signal_21813 ), .Q ( new_AGEMA_signal_21814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C ( clk ), .D ( new_AGEMA_signal_21819 ), .Q ( new_AGEMA_signal_21820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C ( clk ), .D ( new_AGEMA_signal_21825 ), .Q ( new_AGEMA_signal_21826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C ( clk ), .D ( new_AGEMA_signal_21831 ), .Q ( new_AGEMA_signal_21832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C ( clk ), .D ( new_AGEMA_signal_21837 ), .Q ( new_AGEMA_signal_21838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C ( clk ), .D ( new_AGEMA_signal_21843 ), .Q ( new_AGEMA_signal_21844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C ( clk ), .D ( new_AGEMA_signal_21849 ), .Q ( new_AGEMA_signal_21850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C ( clk ), .D ( new_AGEMA_signal_21855 ), .Q ( new_AGEMA_signal_21856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C ( clk ), .D ( new_AGEMA_signal_21861 ), .Q ( new_AGEMA_signal_21862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C ( clk ), .D ( new_AGEMA_signal_21867 ), .Q ( new_AGEMA_signal_21868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C ( clk ), .D ( new_AGEMA_signal_21873 ), .Q ( new_AGEMA_signal_21874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C ( clk ), .D ( new_AGEMA_signal_21879 ), .Q ( new_AGEMA_signal_21880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C ( clk ), .D ( new_AGEMA_signal_21885 ), .Q ( new_AGEMA_signal_21886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C ( clk ), .D ( new_AGEMA_signal_21891 ), .Q ( new_AGEMA_signal_21892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C ( clk ), .D ( new_AGEMA_signal_21897 ), .Q ( new_AGEMA_signal_21898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C ( clk ), .D ( new_AGEMA_signal_21903 ), .Q ( new_AGEMA_signal_21904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C ( clk ), .D ( new_AGEMA_signal_21909 ), .Q ( new_AGEMA_signal_21910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C ( clk ), .D ( new_AGEMA_signal_21915 ), .Q ( new_AGEMA_signal_21916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C ( clk ), .D ( new_AGEMA_signal_21921 ), .Q ( new_AGEMA_signal_21922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C ( clk ), .D ( new_AGEMA_signal_21927 ), .Q ( new_AGEMA_signal_21928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C ( clk ), .D ( new_AGEMA_signal_21933 ), .Q ( new_AGEMA_signal_21934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C ( clk ), .D ( new_AGEMA_signal_21939 ), .Q ( new_AGEMA_signal_21940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C ( clk ), .D ( new_AGEMA_signal_21945 ), .Q ( new_AGEMA_signal_21946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C ( clk ), .D ( new_AGEMA_signal_21951 ), .Q ( new_AGEMA_signal_21952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C ( clk ), .D ( new_AGEMA_signal_21957 ), .Q ( new_AGEMA_signal_21958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_21962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C ( clk ), .D ( new_AGEMA_signal_3298 ), .Q ( new_AGEMA_signal_21966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C ( clk ), .D ( new_AGEMA_signal_3299 ), .Q ( new_AGEMA_signal_21970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C ( clk ), .D ( new_AGEMA_signal_3300 ), .Q ( new_AGEMA_signal_21974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C ( clk ), .D ( new_AGEMA_signal_3301 ), .Q ( new_AGEMA_signal_21978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C ( clk ), .D ( new_AGEMA_signal_21985 ), .Q ( new_AGEMA_signal_21986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C ( clk ), .D ( new_AGEMA_signal_21993 ), .Q ( new_AGEMA_signal_21994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C ( clk ), .D ( new_AGEMA_signal_22001 ), .Q ( new_AGEMA_signal_22002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C ( clk ), .D ( new_AGEMA_signal_22009 ), .Q ( new_AGEMA_signal_22010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C ( clk ), .D ( new_AGEMA_signal_22017 ), .Q ( new_AGEMA_signal_22018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_22022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C ( clk ), .D ( new_AGEMA_signal_3678 ), .Q ( new_AGEMA_signal_22026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C ( clk ), .D ( new_AGEMA_signal_3679 ), .Q ( new_AGEMA_signal_22030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C ( clk ), .D ( new_AGEMA_signal_3680 ), .Q ( new_AGEMA_signal_22034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C ( clk ), .D ( new_AGEMA_signal_3681 ), .Q ( new_AGEMA_signal_22038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C ( clk ), .D ( new_AGEMA_signal_22043 ), .Q ( new_AGEMA_signal_22044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C ( clk ), .D ( new_AGEMA_signal_22049 ), .Q ( new_AGEMA_signal_22050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C ( clk ), .D ( new_AGEMA_signal_22055 ), .Q ( new_AGEMA_signal_22056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C ( clk ), .D ( new_AGEMA_signal_22061 ), .Q ( new_AGEMA_signal_22062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C ( clk ), .D ( new_AGEMA_signal_22067 ), .Q ( new_AGEMA_signal_22068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C ( clk ), .D ( new_AGEMA_signal_22075 ), .Q ( new_AGEMA_signal_22076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C ( clk ), .D ( new_AGEMA_signal_22083 ), .Q ( new_AGEMA_signal_22084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C ( clk ), .D ( new_AGEMA_signal_22091 ), .Q ( new_AGEMA_signal_22092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C ( clk ), .D ( new_AGEMA_signal_22099 ), .Q ( new_AGEMA_signal_22100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C ( clk ), .D ( new_AGEMA_signal_22107 ), .Q ( new_AGEMA_signal_22108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C ( clk ), .D ( new_AGEMA_signal_22123 ), .Q ( new_AGEMA_signal_22124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C ( clk ), .D ( new_AGEMA_signal_22129 ), .Q ( new_AGEMA_signal_22130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C ( clk ), .D ( new_AGEMA_signal_22135 ), .Q ( new_AGEMA_signal_22136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C ( clk ), .D ( new_AGEMA_signal_22141 ), .Q ( new_AGEMA_signal_22142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C ( clk ), .D ( new_AGEMA_signal_22147 ), .Q ( new_AGEMA_signal_22148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C ( clk ), .D ( new_AGEMA_signal_22173 ), .Q ( new_AGEMA_signal_22174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C ( clk ), .D ( new_AGEMA_signal_22179 ), .Q ( new_AGEMA_signal_22180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C ( clk ), .D ( new_AGEMA_signal_22185 ), .Q ( new_AGEMA_signal_22186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C ( clk ), .D ( new_AGEMA_signal_22191 ), .Q ( new_AGEMA_signal_22192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C ( clk ), .D ( new_AGEMA_signal_22197 ), .Q ( new_AGEMA_signal_22198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C ( clk ), .D ( new_AGEMA_signal_22203 ), .Q ( new_AGEMA_signal_22204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C ( clk ), .D ( new_AGEMA_signal_22209 ), .Q ( new_AGEMA_signal_22210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C ( clk ), .D ( new_AGEMA_signal_22215 ), .Q ( new_AGEMA_signal_22216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C ( clk ), .D ( new_AGEMA_signal_22221 ), .Q ( new_AGEMA_signal_22222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C ( clk ), .D ( new_AGEMA_signal_22227 ), .Q ( new_AGEMA_signal_22228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C ( clk ), .D ( new_AGEMA_signal_22235 ), .Q ( new_AGEMA_signal_22236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C ( clk ), .D ( new_AGEMA_signal_22243 ), .Q ( new_AGEMA_signal_22244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C ( clk ), .D ( new_AGEMA_signal_22251 ), .Q ( new_AGEMA_signal_22252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C ( clk ), .D ( new_AGEMA_signal_22259 ), .Q ( new_AGEMA_signal_22260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C ( clk ), .D ( new_AGEMA_signal_22267 ), .Q ( new_AGEMA_signal_22268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C ( clk ), .D ( new_AGEMA_signal_22275 ), .Q ( new_AGEMA_signal_22276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C ( clk ), .D ( new_AGEMA_signal_22283 ), .Q ( new_AGEMA_signal_22284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C ( clk ), .D ( new_AGEMA_signal_22291 ), .Q ( new_AGEMA_signal_22292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C ( clk ), .D ( new_AGEMA_signal_22299 ), .Q ( new_AGEMA_signal_22300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C ( clk ), .D ( new_AGEMA_signal_22307 ), .Q ( new_AGEMA_signal_22308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C ( clk ), .D ( new_AGEMA_signal_22313 ), .Q ( new_AGEMA_signal_22314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C ( clk ), .D ( new_AGEMA_signal_22319 ), .Q ( new_AGEMA_signal_22320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C ( clk ), .D ( new_AGEMA_signal_22325 ), .Q ( new_AGEMA_signal_22326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C ( clk ), .D ( new_AGEMA_signal_22331 ), .Q ( new_AGEMA_signal_22332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C ( clk ), .D ( new_AGEMA_signal_22337 ), .Q ( new_AGEMA_signal_22338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C ( clk ), .D ( new_AGEMA_signal_22343 ), .Q ( new_AGEMA_signal_22344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C ( clk ), .D ( new_AGEMA_signal_22349 ), .Q ( new_AGEMA_signal_22350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C ( clk ), .D ( new_AGEMA_signal_22355 ), .Q ( new_AGEMA_signal_22356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C ( clk ), .D ( new_AGEMA_signal_22361 ), .Q ( new_AGEMA_signal_22362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C ( clk ), .D ( new_AGEMA_signal_22367 ), .Q ( new_AGEMA_signal_22368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_22382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C ( clk ), .D ( new_AGEMA_signal_3086 ), .Q ( new_AGEMA_signal_22386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C ( clk ), .D ( new_AGEMA_signal_3087 ), .Q ( new_AGEMA_signal_22390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C ( clk ), .D ( new_AGEMA_signal_3088 ), .Q ( new_AGEMA_signal_22394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C ( clk ), .D ( new_AGEMA_signal_3089 ), .Q ( new_AGEMA_signal_22398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_22402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C ( clk ), .D ( new_AGEMA_signal_3466 ), .Q ( new_AGEMA_signal_22406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C ( clk ), .D ( new_AGEMA_signal_3467 ), .Q ( new_AGEMA_signal_22410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C ( clk ), .D ( new_AGEMA_signal_3468 ), .Q ( new_AGEMA_signal_22414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C ( clk ), .D ( new_AGEMA_signal_3469 ), .Q ( new_AGEMA_signal_22418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_22422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C ( clk ), .D ( new_AGEMA_signal_3498 ), .Q ( new_AGEMA_signal_22426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C ( clk ), .D ( new_AGEMA_signal_3499 ), .Q ( new_AGEMA_signal_22430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C ( clk ), .D ( new_AGEMA_signal_3500 ), .Q ( new_AGEMA_signal_22434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C ( clk ), .D ( new_AGEMA_signal_3501 ), .Q ( new_AGEMA_signal_22438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_22452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C ( clk ), .D ( new_AGEMA_signal_3054 ), .Q ( new_AGEMA_signal_22458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C ( clk ), .D ( new_AGEMA_signal_3055 ), .Q ( new_AGEMA_signal_22464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C ( clk ), .D ( new_AGEMA_signal_3056 ), .Q ( new_AGEMA_signal_22470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C ( clk ), .D ( new_AGEMA_signal_3057 ), .Q ( new_AGEMA_signal_22476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C ( clk ), .D ( new_AGEMA_signal_22513 ), .Q ( new_AGEMA_signal_22514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C ( clk ), .D ( new_AGEMA_signal_22521 ), .Q ( new_AGEMA_signal_22522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C ( clk ), .D ( new_AGEMA_signal_22529 ), .Q ( new_AGEMA_signal_22530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C ( clk ), .D ( new_AGEMA_signal_22537 ), .Q ( new_AGEMA_signal_22538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C ( clk ), .D ( new_AGEMA_signal_22545 ), .Q ( new_AGEMA_signal_22546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C ( clk ), .D ( new_AGEMA_signal_22553 ), .Q ( new_AGEMA_signal_22554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C ( clk ), .D ( new_AGEMA_signal_22561 ), .Q ( new_AGEMA_signal_22562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C ( clk ), .D ( new_AGEMA_signal_22569 ), .Q ( new_AGEMA_signal_22570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C ( clk ), .D ( new_AGEMA_signal_22577 ), .Q ( new_AGEMA_signal_22578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C ( clk ), .D ( new_AGEMA_signal_22585 ), .Q ( new_AGEMA_signal_22586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C ( clk ), .D ( new_AGEMA_signal_22593 ), .Q ( new_AGEMA_signal_22594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C ( clk ), .D ( new_AGEMA_signal_22601 ), .Q ( new_AGEMA_signal_22602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C ( clk ), .D ( new_AGEMA_signal_22609 ), .Q ( new_AGEMA_signal_22610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C ( clk ), .D ( new_AGEMA_signal_22617 ), .Q ( new_AGEMA_signal_22618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C ( clk ), .D ( new_AGEMA_signal_22625 ), .Q ( new_AGEMA_signal_22626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C ( clk ), .D ( new_AGEMA_signal_22633 ), .Q ( new_AGEMA_signal_22634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C ( clk ), .D ( new_AGEMA_signal_22641 ), .Q ( new_AGEMA_signal_22642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C ( clk ), .D ( new_AGEMA_signal_22649 ), .Q ( new_AGEMA_signal_22650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C ( clk ), .D ( new_AGEMA_signal_22657 ), .Q ( new_AGEMA_signal_22658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C ( clk ), .D ( new_AGEMA_signal_22665 ), .Q ( new_AGEMA_signal_22666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_22672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C ( clk ), .D ( new_AGEMA_signal_3170 ), .Q ( new_AGEMA_signal_22678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C ( clk ), .D ( new_AGEMA_signal_3171 ), .Q ( new_AGEMA_signal_22684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C ( clk ), .D ( new_AGEMA_signal_3172 ), .Q ( new_AGEMA_signal_22690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C ( clk ), .D ( new_AGEMA_signal_3173 ), .Q ( new_AGEMA_signal_22696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C ( clk ), .D ( new_AGEMA_signal_22705 ), .Q ( new_AGEMA_signal_22706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C ( clk ), .D ( new_AGEMA_signal_22715 ), .Q ( new_AGEMA_signal_22716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C ( clk ), .D ( new_AGEMA_signal_22725 ), .Q ( new_AGEMA_signal_22726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C ( clk ), .D ( new_AGEMA_signal_22735 ), .Q ( new_AGEMA_signal_22736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C ( clk ), .D ( new_AGEMA_signal_22745 ), .Q ( new_AGEMA_signal_22746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C ( clk ), .D ( new_AGEMA_signal_22753 ), .Q ( new_AGEMA_signal_22754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C ( clk ), .D ( new_AGEMA_signal_22761 ), .Q ( new_AGEMA_signal_22762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C ( clk ), .D ( new_AGEMA_signal_22769 ), .Q ( new_AGEMA_signal_22770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C ( clk ), .D ( new_AGEMA_signal_22777 ), .Q ( new_AGEMA_signal_22778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C ( clk ), .D ( new_AGEMA_signal_22785 ), .Q ( new_AGEMA_signal_22786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C ( clk ), .D ( new_AGEMA_signal_22793 ), .Q ( new_AGEMA_signal_22794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C ( clk ), .D ( new_AGEMA_signal_22801 ), .Q ( new_AGEMA_signal_22802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C ( clk ), .D ( new_AGEMA_signal_22809 ), .Q ( new_AGEMA_signal_22810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C ( clk ), .D ( new_AGEMA_signal_22817 ), .Q ( new_AGEMA_signal_22818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C ( clk ), .D ( new_AGEMA_signal_22825 ), .Q ( new_AGEMA_signal_22826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C ( clk ), .D ( new_AGEMA_signal_22833 ), .Q ( new_AGEMA_signal_22834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C ( clk ), .D ( new_AGEMA_signal_22841 ), .Q ( new_AGEMA_signal_22842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C ( clk ), .D ( new_AGEMA_signal_22849 ), .Q ( new_AGEMA_signal_22850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C ( clk ), .D ( new_AGEMA_signal_22857 ), .Q ( new_AGEMA_signal_22858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C ( clk ), .D ( new_AGEMA_signal_22865 ), .Q ( new_AGEMA_signal_22866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_22902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C ( clk ), .D ( new_AGEMA_signal_3306 ), .Q ( new_AGEMA_signal_22908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C ( clk ), .D ( new_AGEMA_signal_3307 ), .Q ( new_AGEMA_signal_22914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C ( clk ), .D ( new_AGEMA_signal_3308 ), .Q ( new_AGEMA_signal_22920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C ( clk ), .D ( new_AGEMA_signal_3309 ), .Q ( new_AGEMA_signal_22926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C ( clk ), .D ( new_AGEMA_signal_22955 ), .Q ( new_AGEMA_signal_22956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C ( clk ), .D ( new_AGEMA_signal_22965 ), .Q ( new_AGEMA_signal_22966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C ( clk ), .D ( new_AGEMA_signal_22975 ), .Q ( new_AGEMA_signal_22976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C ( clk ), .D ( new_AGEMA_signal_22985 ), .Q ( new_AGEMA_signal_22986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C ( clk ), .D ( new_AGEMA_signal_22995 ), .Q ( new_AGEMA_signal_22996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C ( clk ), .D ( new_AGEMA_signal_23003 ), .Q ( new_AGEMA_signal_23004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C ( clk ), .D ( new_AGEMA_signal_23011 ), .Q ( new_AGEMA_signal_23012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C ( clk ), .D ( new_AGEMA_signal_23019 ), .Q ( new_AGEMA_signal_23020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C ( clk ), .D ( new_AGEMA_signal_23027 ), .Q ( new_AGEMA_signal_23028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C ( clk ), .D ( new_AGEMA_signal_23035 ), .Q ( new_AGEMA_signal_23036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C ( clk ), .D ( new_AGEMA_signal_23073 ), .Q ( new_AGEMA_signal_23074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C ( clk ), .D ( new_AGEMA_signal_23081 ), .Q ( new_AGEMA_signal_23082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C ( clk ), .D ( new_AGEMA_signal_23089 ), .Q ( new_AGEMA_signal_23090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C ( clk ), .D ( new_AGEMA_signal_23097 ), .Q ( new_AGEMA_signal_23098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C ( clk ), .D ( new_AGEMA_signal_23105 ), .Q ( new_AGEMA_signal_23106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C ( clk ), .D ( new_AGEMA_signal_23113 ), .Q ( new_AGEMA_signal_23114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C ( clk ), .D ( new_AGEMA_signal_23121 ), .Q ( new_AGEMA_signal_23122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C ( clk ), .D ( new_AGEMA_signal_23129 ), .Q ( new_AGEMA_signal_23130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C ( clk ), .D ( new_AGEMA_signal_23137 ), .Q ( new_AGEMA_signal_23138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C ( clk ), .D ( new_AGEMA_signal_23145 ), .Q ( new_AGEMA_signal_23146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C ( clk ), .D ( new_AGEMA_signal_19795 ), .Q ( new_AGEMA_signal_23152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C ( clk ), .D ( new_AGEMA_signal_19799 ), .Q ( new_AGEMA_signal_23158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C ( clk ), .D ( new_AGEMA_signal_19803 ), .Q ( new_AGEMA_signal_23164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C ( clk ), .D ( new_AGEMA_signal_19807 ), .Q ( new_AGEMA_signal_23170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C ( clk ), .D ( new_AGEMA_signal_19811 ), .Q ( new_AGEMA_signal_23176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C ( clk ), .D ( new_AGEMA_signal_23203 ), .Q ( new_AGEMA_signal_23204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C ( clk ), .D ( new_AGEMA_signal_23211 ), .Q ( new_AGEMA_signal_23212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C ( clk ), .D ( new_AGEMA_signal_23219 ), .Q ( new_AGEMA_signal_23220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C ( clk ), .D ( new_AGEMA_signal_23227 ), .Q ( new_AGEMA_signal_23228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C ( clk ), .D ( new_AGEMA_signal_23235 ), .Q ( new_AGEMA_signal_23236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C ( clk ), .D ( new_AGEMA_signal_20355 ), .Q ( new_AGEMA_signal_23362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C ( clk ), .D ( new_AGEMA_signal_20359 ), .Q ( new_AGEMA_signal_23370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C ( clk ), .D ( new_AGEMA_signal_20363 ), .Q ( new_AGEMA_signal_23378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C ( clk ), .D ( new_AGEMA_signal_20367 ), .Q ( new_AGEMA_signal_23386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C ( clk ), .D ( new_AGEMA_signal_20371 ), .Q ( new_AGEMA_signal_23394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_23452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C ( clk ), .D ( new_AGEMA_signal_3186 ), .Q ( new_AGEMA_signal_23460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C ( clk ), .D ( new_AGEMA_signal_3187 ), .Q ( new_AGEMA_signal_23468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C ( clk ), .D ( new_AGEMA_signal_3188 ), .Q ( new_AGEMA_signal_23476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C ( clk ), .D ( new_AGEMA_signal_3189 ), .Q ( new_AGEMA_signal_23484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C ( clk ), .D ( new_AGEMA_signal_19593 ), .Q ( new_AGEMA_signal_23492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C ( clk ), .D ( new_AGEMA_signal_19595 ), .Q ( new_AGEMA_signal_23500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C ( clk ), .D ( new_AGEMA_signal_19597 ), .Q ( new_AGEMA_signal_23508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C ( clk ), .D ( new_AGEMA_signal_19599 ), .Q ( new_AGEMA_signal_23516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C ( clk ), .D ( new_AGEMA_signal_19601 ), .Q ( new_AGEMA_signal_23524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C ( clk ), .D ( new_AGEMA_signal_23533 ), .Q ( new_AGEMA_signal_23534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C ( clk ), .D ( new_AGEMA_signal_23543 ), .Q ( new_AGEMA_signal_23544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C ( clk ), .D ( new_AGEMA_signal_23553 ), .Q ( new_AGEMA_signal_23554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C ( clk ), .D ( new_AGEMA_signal_23563 ), .Q ( new_AGEMA_signal_23564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C ( clk ), .D ( new_AGEMA_signal_23573 ), .Q ( new_AGEMA_signal_23574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C ( clk ), .D ( new_AGEMA_signal_20055 ), .Q ( new_AGEMA_signal_23582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C ( clk ), .D ( new_AGEMA_signal_20059 ), .Q ( new_AGEMA_signal_23590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C ( clk ), .D ( new_AGEMA_signal_20063 ), .Q ( new_AGEMA_signal_23598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C ( clk ), .D ( new_AGEMA_signal_20067 ), .Q ( new_AGEMA_signal_23606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C ( clk ), .D ( new_AGEMA_signal_20071 ), .Q ( new_AGEMA_signal_23614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_23702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C ( clk ), .D ( new_AGEMA_signal_2774 ), .Q ( new_AGEMA_signal_23710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C ( clk ), .D ( new_AGEMA_signal_2775 ), .Q ( new_AGEMA_signal_23718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C ( clk ), .D ( new_AGEMA_signal_2776 ), .Q ( new_AGEMA_signal_23726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C ( clk ), .D ( new_AGEMA_signal_2777 ), .Q ( new_AGEMA_signal_23734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_23782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C ( clk ), .D ( new_AGEMA_signal_3430 ), .Q ( new_AGEMA_signal_23790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C ( clk ), .D ( new_AGEMA_signal_3431 ), .Q ( new_AGEMA_signal_23798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C ( clk ), .D ( new_AGEMA_signal_3432 ), .Q ( new_AGEMA_signal_23806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C ( clk ), .D ( new_AGEMA_signal_3433 ), .Q ( new_AGEMA_signal_23814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_24002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C ( clk ), .D ( new_AGEMA_signal_3166 ), .Q ( new_AGEMA_signal_24012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C ( clk ), .D ( new_AGEMA_signal_3167 ), .Q ( new_AGEMA_signal_24022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C ( clk ), .D ( new_AGEMA_signal_3168 ), .Q ( new_AGEMA_signal_24032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C ( clk ), .D ( new_AGEMA_signal_3169 ), .Q ( new_AGEMA_signal_24042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7677 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_24452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7689 ( .C ( clk ), .D ( new_AGEMA_signal_2602 ), .Q ( new_AGEMA_signal_24464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7701 ( .C ( clk ), .D ( new_AGEMA_signal_2603 ), .Q ( new_AGEMA_signal_24476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7713 ( .C ( clk ), .D ( new_AGEMA_signal_2604 ), .Q ( new_AGEMA_signal_24488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7725 ( .C ( clk ), .D ( new_AGEMA_signal_2605 ), .Q ( new_AGEMA_signal_24500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7739 ( .C ( clk ), .D ( new_AGEMA_signal_24513 ), .Q ( new_AGEMA_signal_24514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7753 ( .C ( clk ), .D ( new_AGEMA_signal_24527 ), .Q ( new_AGEMA_signal_24528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7767 ( .C ( clk ), .D ( new_AGEMA_signal_24541 ), .Q ( new_AGEMA_signal_24542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7781 ( .C ( clk ), .D ( new_AGEMA_signal_24555 ), .Q ( new_AGEMA_signal_24556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7795 ( .C ( clk ), .D ( new_AGEMA_signal_24569 ), .Q ( new_AGEMA_signal_24570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7849 ( .C ( clk ), .D ( new_AGEMA_signal_24623 ), .Q ( new_AGEMA_signal_24624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7863 ( .C ( clk ), .D ( new_AGEMA_signal_24637 ), .Q ( new_AGEMA_signal_24638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7877 ( .C ( clk ), .D ( new_AGEMA_signal_24651 ), .Q ( new_AGEMA_signal_24652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7891 ( .C ( clk ), .D ( new_AGEMA_signal_24665 ), .Q ( new_AGEMA_signal_24666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7905 ( .C ( clk ), .D ( new_AGEMA_signal_24679 ), .Q ( new_AGEMA_signal_24680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8029 ( .C ( clk ), .D ( new_AGEMA_signal_24803 ), .Q ( new_AGEMA_signal_24804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8045 ( .C ( clk ), .D ( new_AGEMA_signal_24819 ), .Q ( new_AGEMA_signal_24820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8061 ( .C ( clk ), .D ( new_AGEMA_signal_24835 ), .Q ( new_AGEMA_signal_24836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8077 ( .C ( clk ), .D ( new_AGEMA_signal_24851 ), .Q ( new_AGEMA_signal_24852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8093 ( .C ( clk ), .D ( new_AGEMA_signal_24867 ), .Q ( new_AGEMA_signal_24868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8139 ( .C ( clk ), .D ( new_AGEMA_signal_24913 ), .Q ( new_AGEMA_signal_24914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8155 ( .C ( clk ), .D ( new_AGEMA_signal_24929 ), .Q ( new_AGEMA_signal_24930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8171 ( .C ( clk ), .D ( new_AGEMA_signal_24945 ), .Q ( new_AGEMA_signal_24946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8187 ( .C ( clk ), .D ( new_AGEMA_signal_24961 ), .Q ( new_AGEMA_signal_24962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8203 ( .C ( clk ), .D ( new_AGEMA_signal_24977 ), .Q ( new_AGEMA_signal_24978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8387 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_25162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8403 ( .C ( clk ), .D ( new_AGEMA_signal_2610 ), .Q ( new_AGEMA_signal_25178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8419 ( .C ( clk ), .D ( new_AGEMA_signal_2611 ), .Q ( new_AGEMA_signal_25194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8435 ( .C ( clk ), .D ( new_AGEMA_signal_2612 ), .Q ( new_AGEMA_signal_25210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8451 ( .C ( clk ), .D ( new_AGEMA_signal_2613 ), .Q ( new_AGEMA_signal_25226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8519 ( .C ( clk ), .D ( new_AGEMA_signal_25293 ), .Q ( new_AGEMA_signal_25294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8537 ( .C ( clk ), .D ( new_AGEMA_signal_25311 ), .Q ( new_AGEMA_signal_25312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8555 ( .C ( clk ), .D ( new_AGEMA_signal_25329 ), .Q ( new_AGEMA_signal_25330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8573 ( .C ( clk ), .D ( new_AGEMA_signal_25347 ), .Q ( new_AGEMA_signal_25348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8591 ( .C ( clk ), .D ( new_AGEMA_signal_25365 ), .Q ( new_AGEMA_signal_25366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8769 ( .C ( clk ), .D ( new_AGEMA_signal_25543 ), .Q ( new_AGEMA_signal_25544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8789 ( .C ( clk ), .D ( new_AGEMA_signal_25563 ), .Q ( new_AGEMA_signal_25564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8809 ( .C ( clk ), .D ( new_AGEMA_signal_25583 ), .Q ( new_AGEMA_signal_25584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8829 ( .C ( clk ), .D ( new_AGEMA_signal_25603 ), .Q ( new_AGEMA_signal_25604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8849 ( .C ( clk ), .D ( new_AGEMA_signal_25623 ), .Q ( new_AGEMA_signal_25624 ) ) ;

    /* cells in depth 10 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1983 ( .ina ({new_AGEMA_signal_19421, new_AGEMA_signal_19417, new_AGEMA_signal_19413, new_AGEMA_signal_19409, new_AGEMA_signal_19405}), .inb ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, n1928}), .clk ( clk ), .rnd ({Fresh[8639], Fresh[8638], Fresh[8637], Fresh[8636], Fresh[8635], Fresh[8634], Fresh[8633], Fresh[8632], Fresh[8631], Fresh[8630], Fresh[8629], Fresh[8628], Fresh[8627], Fresh[8626], Fresh[8625]}), .outt ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, n1934}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U1998 ( .ina ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, n1931}), .inb ({new_AGEMA_signal_19441, new_AGEMA_signal_19437, new_AGEMA_signal_19433, new_AGEMA_signal_19429, new_AGEMA_signal_19425}), .clk ( clk ), .rnd ({Fresh[8654], Fresh[8653], Fresh[8652], Fresh[8651], Fresh[8650], Fresh[8649], Fresh[8648], Fresh[8647], Fresh[8646], Fresh[8645], Fresh[8644], Fresh[8643], Fresh[8642], Fresh[8641], Fresh[8640]}), .outt ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, n1932}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2015 ( .ina ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n1939}), .inb ({new_AGEMA_signal_19451, new_AGEMA_signal_19449, new_AGEMA_signal_19447, new_AGEMA_signal_19445, new_AGEMA_signal_19443}), .clk ( clk ), .rnd ({Fresh[8669], Fresh[8668], Fresh[8667], Fresh[8666], Fresh[8665], Fresh[8664], Fresh[8663], Fresh[8662], Fresh[8661], Fresh[8660], Fresh[8659], Fresh[8658], Fresh[8657], Fresh[8656], Fresh[8655]}), .outt ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, n1940}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2033 ( .ina ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, n1948}), .inb ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, n1947}), .clk ( clk ), .rnd ({Fresh[8684], Fresh[8683], Fresh[8682], Fresh[8681], Fresh[8680], Fresh[8679], Fresh[8678], Fresh[8677], Fresh[8676], Fresh[8675], Fresh[8674], Fresh[8673], Fresh[8672], Fresh[8671], Fresh[8670]}), .outt ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, n1961}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2050 ( .ina ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n1954}), .inb ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, n1953}), .clk ( clk ), .rnd ({Fresh[8699], Fresh[8698], Fresh[8697], Fresh[8696], Fresh[8695], Fresh[8694], Fresh[8693], Fresh[8692], Fresh[8691], Fresh[8690], Fresh[8689], Fresh[8688], Fresh[8687], Fresh[8686], Fresh[8685]}), .outt ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, n1955}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2066 ( .ina ({new_AGEMA_signal_19461, new_AGEMA_signal_19459, new_AGEMA_signal_19457, new_AGEMA_signal_19455, new_AGEMA_signal_19453}), .inb ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, n1965}), .clk ( clk ), .rnd ({Fresh[8714], Fresh[8713], Fresh[8712], Fresh[8711], Fresh[8710], Fresh[8709], Fresh[8708], Fresh[8707], Fresh[8706], Fresh[8705], Fresh[8704], Fresh[8703], Fresh[8702], Fresh[8701], Fresh[8700]}), .outt ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n1967}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2085 ( .ina ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, n1970}), .inb ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, n1969}), .clk ( clk ), .rnd ({Fresh[8729], Fresh[8728], Fresh[8727], Fresh[8726], Fresh[8725], Fresh[8724], Fresh[8723], Fresh[8722], Fresh[8721], Fresh[8720], Fresh[8719], Fresh[8718], Fresh[8717], Fresh[8716], Fresh[8715]}), .outt ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, new_AGEMA_signal_3851, new_AGEMA_signal_3850, n1984}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2103 ( .ina ({new_AGEMA_signal_19481, new_AGEMA_signal_19477, new_AGEMA_signal_19473, new_AGEMA_signal_19469, new_AGEMA_signal_19465}), .inb ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, n1975}), .clk ( clk ), .rnd ({Fresh[8744], Fresh[8743], Fresh[8742], Fresh[8741], Fresh[8740], Fresh[8739], Fresh[8738], Fresh[8737], Fresh[8736], Fresh[8735], Fresh[8734], Fresh[8733], Fresh[8732], Fresh[8731], Fresh[8730]}), .outt ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, new_AGEMA_signal_3542, n1977}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2108 ( .ina ({new_AGEMA_signal_19491, new_AGEMA_signal_19489, new_AGEMA_signal_19487, new_AGEMA_signal_19485, new_AGEMA_signal_19483}), .inb ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, n1980}), .clk ( clk ), .rnd ({Fresh[8759], Fresh[8758], Fresh[8757], Fresh[8756], Fresh[8755], Fresh[8754], Fresh[8753], Fresh[8752], Fresh[8751], Fresh[8750], Fresh[8749], Fresh[8748], Fresh[8747], Fresh[8746], Fresh[8745]}), .outt ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n1981}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2115 ( .ina ({new_AGEMA_signal_19511, new_AGEMA_signal_19507, new_AGEMA_signal_19503, new_AGEMA_signal_19499, new_AGEMA_signal_19495}), .inb ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n1986}), .clk ( clk ), .rnd ({Fresh[8774], Fresh[8773], Fresh[8772], Fresh[8771], Fresh[8770], Fresh[8769], Fresh[8768], Fresh[8767], Fresh[8766], Fresh[8765], Fresh[8764], Fresh[8763], Fresh[8762], Fresh[8761], Fresh[8760]}), .outt ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n1987}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2127 ( .ina ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, n1997}), .inb ({new_AGEMA_signal_19521, new_AGEMA_signal_19519, new_AGEMA_signal_19517, new_AGEMA_signal_19515, new_AGEMA_signal_19513}), .clk ( clk ), .rnd ({Fresh[8789], Fresh[8788], Fresh[8787], Fresh[8786], Fresh[8785], Fresh[8784], Fresh[8783], Fresh[8782], Fresh[8781], Fresh[8780], Fresh[8779], Fresh[8778], Fresh[8777], Fresh[8776], Fresh[8775]}), .outt ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, n1998}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2146 ( .ina ({new_AGEMA_signal_19541, new_AGEMA_signal_19537, new_AGEMA_signal_19533, new_AGEMA_signal_19529, new_AGEMA_signal_19525}), .inb ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n2007}), .clk ( clk ), .rnd ({Fresh[8804], Fresh[8803], Fresh[8802], Fresh[8801], Fresh[8800], Fresh[8799], Fresh[8798], Fresh[8797], Fresh[8796], Fresh[8795], Fresh[8794], Fresh[8793], Fresh[8792], Fresh[8791], Fresh[8790]}), .outt ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, n2010}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2162 ( .ina ({new_AGEMA_signal_19561, new_AGEMA_signal_19557, new_AGEMA_signal_19553, new_AGEMA_signal_19549, new_AGEMA_signal_19545}), .inb ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, n2021}), .clk ( clk ), .rnd ({Fresh[8819], Fresh[8818], Fresh[8817], Fresh[8816], Fresh[8815], Fresh[8814], Fresh[8813], Fresh[8812], Fresh[8811], Fresh[8810], Fresh[8809], Fresh[8808], Fresh[8807], Fresh[8806], Fresh[8805]}), .outt ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, n2024}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2177 ( .ina ({new_AGEMA_signal_19571, new_AGEMA_signal_19569, new_AGEMA_signal_19567, new_AGEMA_signal_19565, new_AGEMA_signal_19563}), .inb ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, n2032}), .clk ( clk ), .rnd ({Fresh[8834], Fresh[8833], Fresh[8832], Fresh[8831], Fresh[8830], Fresh[8829], Fresh[8828], Fresh[8827], Fresh[8826], Fresh[8825], Fresh[8824], Fresh[8823], Fresh[8822], Fresh[8821], Fresh[8820]}), .outt ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, n2035}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2186 ( .ina ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2041}), .inb ({new_AGEMA_signal_19581, new_AGEMA_signal_19579, new_AGEMA_signal_19577, new_AGEMA_signal_19575, new_AGEMA_signal_19573}), .clk ( clk ), .rnd ({Fresh[8849], Fresh[8848], Fresh[8847], Fresh[8846], Fresh[8845], Fresh[8844], Fresh[8843], Fresh[8842], Fresh[8841], Fresh[8840], Fresh[8839], Fresh[8838], Fresh[8837], Fresh[8836], Fresh[8835]}), .outt ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, new_AGEMA_signal_3566, n2054}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2190 ( .ina ({new_AGEMA_signal_19591, new_AGEMA_signal_19589, new_AGEMA_signal_19587, new_AGEMA_signal_19585, new_AGEMA_signal_19583}), .inb ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, n2043}), .clk ( clk ), .rnd ({Fresh[8864], Fresh[8863], Fresh[8862], Fresh[8861], Fresh[8860], Fresh[8859], Fresh[8858], Fresh[8857], Fresh[8856], Fresh[8855], Fresh[8854], Fresh[8853], Fresh[8852], Fresh[8851], Fresh[8850]}), .outt ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2048}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2195 ( .ina ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, new_AGEMA_signal_3146, n2046}), .inb ({new_AGEMA_signal_19601, new_AGEMA_signal_19599, new_AGEMA_signal_19597, new_AGEMA_signal_19595, new_AGEMA_signal_19593}), .clk ( clk ), .rnd ({Fresh[8879], Fresh[8878], Fresh[8877], Fresh[8876], Fresh[8875], Fresh[8874], Fresh[8873], Fresh[8872], Fresh[8871], Fresh[8870], Fresh[8869], Fresh[8868], Fresh[8867], Fresh[8866], Fresh[8865]}), .outt ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, n2047}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2206 ( .ina ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2058}), .inb ({new_AGEMA_signal_19621, new_AGEMA_signal_19617, new_AGEMA_signal_19613, new_AGEMA_signal_19609, new_AGEMA_signal_19605}), .clk ( clk ), .rnd ({Fresh[8894], Fresh[8893], Fresh[8892], Fresh[8891], Fresh[8890], Fresh[8889], Fresh[8888], Fresh[8887], Fresh[8886], Fresh[8885], Fresh[8884], Fresh[8883], Fresh[8882], Fresh[8881], Fresh[8880]}), .outt ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, new_AGEMA_signal_3578, n2059}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2213 ( .ina ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, n2063}), .inb ({new_AGEMA_signal_19641, new_AGEMA_signal_19637, new_AGEMA_signal_19633, new_AGEMA_signal_19629, new_AGEMA_signal_19625}), .clk ( clk ), .rnd ({Fresh[8909], Fresh[8908], Fresh[8907], Fresh[8906], Fresh[8905], Fresh[8904], Fresh[8903], Fresh[8902], Fresh[8901], Fresh[8900], Fresh[8899], Fresh[8898], Fresh[8897], Fresh[8896], Fresh[8895]}), .outt ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2064}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2229 ( .ina ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2076}), .inb ({new_AGEMA_signal_19661, new_AGEMA_signal_19657, new_AGEMA_signal_19653, new_AGEMA_signal_19649, new_AGEMA_signal_19645}), .clk ( clk ), .rnd ({Fresh[8924], Fresh[8923], Fresh[8922], Fresh[8921], Fresh[8920], Fresh[8919], Fresh[8918], Fresh[8917], Fresh[8916], Fresh[8915], Fresh[8914], Fresh[8913], Fresh[8912], Fresh[8911], Fresh[8910]}), .outt ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, n2077}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2249 ( .ina ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, n2090}), .inb ({new_AGEMA_signal_19671, new_AGEMA_signal_19669, new_AGEMA_signal_19667, new_AGEMA_signal_19665, new_AGEMA_signal_19663}), .clk ( clk ), .rnd ({Fresh[8939], Fresh[8938], Fresh[8937], Fresh[8936], Fresh[8935], Fresh[8934], Fresh[8933], Fresh[8932], Fresh[8931], Fresh[8930], Fresh[8929], Fresh[8928], Fresh[8927], Fresh[8926], Fresh[8925]}), .outt ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, n2158}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2255 ( .ina ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, n2093}), .inb ({new_AGEMA_signal_19681, new_AGEMA_signal_19679, new_AGEMA_signal_19677, new_AGEMA_signal_19675, new_AGEMA_signal_19673}), .clk ( clk ), .rnd ({Fresh[8954], Fresh[8953], Fresh[8952], Fresh[8951], Fresh[8950], Fresh[8949], Fresh[8948], Fresh[8947], Fresh[8946], Fresh[8945], Fresh[8944], Fresh[8943], Fresh[8942], Fresh[8941], Fresh[8940]}), .outt ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2095}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2274 ( .ina ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, n2116}), .inb ({new_AGEMA_signal_19691, new_AGEMA_signal_19689, new_AGEMA_signal_19687, new_AGEMA_signal_19685, new_AGEMA_signal_19683}), .clk ( clk ), .rnd ({Fresh[8969], Fresh[8968], Fresh[8967], Fresh[8966], Fresh[8965], Fresh[8964], Fresh[8963], Fresh[8962], Fresh[8961], Fresh[8960], Fresh[8959], Fresh[8958], Fresh[8957], Fresh[8956], Fresh[8955]}), .outt ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, new_AGEMA_signal_3899, new_AGEMA_signal_3898, n2117}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2283 ( .ina ({new_AGEMA_signal_19711, new_AGEMA_signal_19707, new_AGEMA_signal_19703, new_AGEMA_signal_19699, new_AGEMA_signal_19695}), .inb ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, n2120}), .clk ( clk ), .rnd ({Fresh[8984], Fresh[8983], Fresh[8982], Fresh[8981], Fresh[8980], Fresh[8979], Fresh[8978], Fresh[8977], Fresh[8976], Fresh[8975], Fresh[8974], Fresh[8973], Fresh[8972], Fresh[8971], Fresh[8970]}), .outt ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, n2123}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2300 ( .ina ({new_AGEMA_signal_19721, new_AGEMA_signal_19719, new_AGEMA_signal_19717, new_AGEMA_signal_19715, new_AGEMA_signal_19713}), .inb ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, n2134}), .clk ( clk ), .rnd ({Fresh[8999], Fresh[8998], Fresh[8997], Fresh[8996], Fresh[8995], Fresh[8994], Fresh[8993], Fresh[8992], Fresh[8991], Fresh[8990], Fresh[8989], Fresh[8988], Fresh[8987], Fresh[8986], Fresh[8985]}), .outt ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, n2135}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2309 ( .ina ({new_AGEMA_signal_19741, new_AGEMA_signal_19737, new_AGEMA_signal_19733, new_AGEMA_signal_19729, new_AGEMA_signal_19725}), .inb ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2140}), .clk ( clk ), .rnd ({Fresh[9014], Fresh[9013], Fresh[9012], Fresh[9011], Fresh[9010], Fresh[9009], Fresh[9008], Fresh[9007], Fresh[9006], Fresh[9005], Fresh[9004], Fresh[9003], Fresh[9002], Fresh[9001], Fresh[9000]}), .outt ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, n2141}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2327 ( .ina ({new_AGEMA_signal_19771, new_AGEMA_signal_19765, new_AGEMA_signal_19759, new_AGEMA_signal_19753, new_AGEMA_signal_19747}), .inb ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, n2161}), .clk ( clk ), .rnd ({Fresh[9029], Fresh[9028], Fresh[9027], Fresh[9026], Fresh[9025], Fresh[9024], Fresh[9023], Fresh[9022], Fresh[9021], Fresh[9020], Fresh[9019], Fresh[9018], Fresh[9017], Fresh[9016], Fresh[9015]}), .outt ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, n2166}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2331 ( .ina ({new_AGEMA_signal_19791, new_AGEMA_signal_19787, new_AGEMA_signal_19783, new_AGEMA_signal_19779, new_AGEMA_signal_19775}), .inb ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, n2164}), .clk ( clk ), .rnd ({Fresh[9044], Fresh[9043], Fresh[9042], Fresh[9041], Fresh[9040], Fresh[9039], Fresh[9038], Fresh[9037], Fresh[9036], Fresh[9035], Fresh[9034], Fresh[9033], Fresh[9032], Fresh[9031], Fresh[9030]}), .outt ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2165}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2346 ( .ina ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, n2179}), .inb ({new_AGEMA_signal_19811, new_AGEMA_signal_19807, new_AGEMA_signal_19803, new_AGEMA_signal_19799, new_AGEMA_signal_19795}), .clk ( clk ), .rnd ({Fresh[9059], Fresh[9058], Fresh[9057], Fresh[9056], Fresh[9055], Fresh[9054], Fresh[9053], Fresh[9052], Fresh[9051], Fresh[9050], Fresh[9049], Fresh[9048], Fresh[9047], Fresh[9046], Fresh[9045]}), .outt ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2180}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2360 ( .ina ({new_AGEMA_signal_19821, new_AGEMA_signal_19819, new_AGEMA_signal_19817, new_AGEMA_signal_19815, new_AGEMA_signal_19813}), .inb ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, n2192}), .clk ( clk ), .rnd ({Fresh[9074], Fresh[9073], Fresh[9072], Fresh[9071], Fresh[9070], Fresh[9069], Fresh[9068], Fresh[9067], Fresh[9066], Fresh[9065], Fresh[9064], Fresh[9063], Fresh[9062], Fresh[9061], Fresh[9060]}), .outt ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, n2194}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2372 ( .ina ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, n2203}), .inb ({new_AGEMA_signal_19831, new_AGEMA_signal_19829, new_AGEMA_signal_19827, new_AGEMA_signal_19825, new_AGEMA_signal_19823}), .clk ( clk ), .rnd ({Fresh[9089], Fresh[9088], Fresh[9087], Fresh[9086], Fresh[9085], Fresh[9084], Fresh[9083], Fresh[9082], Fresh[9081], Fresh[9080], Fresh[9079], Fresh[9078], Fresh[9077], Fresh[9076], Fresh[9075]}), .outt ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, new_AGEMA_signal_3927, new_AGEMA_signal_3926, n2204}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2389 ( .ina ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, n2224}), .inb ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2223}), .clk ( clk ), .rnd ({Fresh[9104], Fresh[9103], Fresh[9102], Fresh[9101], Fresh[9100], Fresh[9099], Fresh[9098], Fresh[9097], Fresh[9096], Fresh[9095], Fresh[9094], Fresh[9093], Fresh[9092], Fresh[9091], Fresh[9090]}), .outt ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2225}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2394 ( .ina ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, n2229}), .inb ({new_AGEMA_signal_19841, new_AGEMA_signal_19839, new_AGEMA_signal_19837, new_AGEMA_signal_19835, new_AGEMA_signal_19833}), .clk ( clk ), .rnd ({Fresh[9119], Fresh[9118], Fresh[9117], Fresh[9116], Fresh[9115], Fresh[9114], Fresh[9113], Fresh[9112], Fresh[9111], Fresh[9110], Fresh[9109], Fresh[9108], Fresh[9107], Fresh[9106], Fresh[9105]}), .outt ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, n2230}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2400 ( .ina ({new_AGEMA_signal_19851, new_AGEMA_signal_19849, new_AGEMA_signal_19847, new_AGEMA_signal_19845, new_AGEMA_signal_19843}), .inb ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, n2234}), .clk ( clk ), .rnd ({Fresh[9134], Fresh[9133], Fresh[9132], Fresh[9131], Fresh[9130], Fresh[9129], Fresh[9128], Fresh[9127], Fresh[9126], Fresh[9125], Fresh[9124], Fresh[9123], Fresh[9122], Fresh[9121], Fresh[9120]}), .outt ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, n2236}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2412 ( .ina ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2246}), .inb ({new_AGEMA_signal_19871, new_AGEMA_signal_19867, new_AGEMA_signal_19863, new_AGEMA_signal_19859, new_AGEMA_signal_19855}), .clk ( clk ), .rnd ({Fresh[9149], Fresh[9148], Fresh[9147], Fresh[9146], Fresh[9145], Fresh[9144], Fresh[9143], Fresh[9142], Fresh[9141], Fresh[9140], Fresh[9139], Fresh[9138], Fresh[9137], Fresh[9136], Fresh[9135]}), .outt ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2247}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2419 ( .ina ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, n2254}), .inb ({new_AGEMA_signal_19901, new_AGEMA_signal_19895, new_AGEMA_signal_19889, new_AGEMA_signal_19883, new_AGEMA_signal_19877}), .clk ( clk ), .rnd ({Fresh[9164], Fresh[9163], Fresh[9162], Fresh[9161], Fresh[9160], Fresh[9159], Fresh[9158], Fresh[9157], Fresh[9156], Fresh[9155], Fresh[9154], Fresh[9153], Fresh[9152], Fresh[9151], Fresh[9150]}), .outt ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, n2255}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2427 ( .ina ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, new_AGEMA_signal_3266, n2263}), .inb ({new_AGEMA_signal_19921, new_AGEMA_signal_19917, new_AGEMA_signal_19913, new_AGEMA_signal_19909, new_AGEMA_signal_19905}), .clk ( clk ), .rnd ({Fresh[9179], Fresh[9178], Fresh[9177], Fresh[9176], Fresh[9175], Fresh[9174], Fresh[9173], Fresh[9172], Fresh[9171], Fresh[9170], Fresh[9169], Fresh[9168], Fresh[9167], Fresh[9166], Fresh[9165]}), .outt ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, n2264}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2435 ( .ina ({new_AGEMA_signal_19931, new_AGEMA_signal_19929, new_AGEMA_signal_19927, new_AGEMA_signal_19925, new_AGEMA_signal_19923}), .inb ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, n2267}), .clk ( clk ), .rnd ({Fresh[9194], Fresh[9193], Fresh[9192], Fresh[9191], Fresh[9190], Fresh[9189], Fresh[9188], Fresh[9187], Fresh[9186], Fresh[9185], Fresh[9184], Fresh[9183], Fresh[9182], Fresh[9181], Fresh[9180]}), .outt ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2271}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2446 ( .ina ({new_AGEMA_signal_19511, new_AGEMA_signal_19507, new_AGEMA_signal_19503, new_AGEMA_signal_19499, new_AGEMA_signal_19495}), .inb ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, n2279}), .clk ( clk ), .rnd ({Fresh[9209], Fresh[9208], Fresh[9207], Fresh[9206], Fresh[9205], Fresh[9204], Fresh[9203], Fresh[9202], Fresh[9201], Fresh[9200], Fresh[9199], Fresh[9198], Fresh[9197], Fresh[9196], Fresh[9195]}), .outt ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, new_AGEMA_signal_3278, n2280}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2451 ( .ina ({new_AGEMA_signal_19941, new_AGEMA_signal_19939, new_AGEMA_signal_19937, new_AGEMA_signal_19935, new_AGEMA_signal_19933}), .inb ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, n2283}), .clk ( clk ), .rnd ({Fresh[9224], Fresh[9223], Fresh[9222], Fresh[9221], Fresh[9220], Fresh[9219], Fresh[9218], Fresh[9217], Fresh[9216], Fresh[9215], Fresh[9214], Fresh[9213], Fresh[9212], Fresh[9211], Fresh[9210]}), .outt ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2286}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2461 ( .ina ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, n2686}), .inb ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n2289}), .clk ( clk ), .rnd ({Fresh[9239], Fresh[9238], Fresh[9237], Fresh[9236], Fresh[9235], Fresh[9234], Fresh[9233], Fresh[9232], Fresh[9231], Fresh[9230], Fresh[9229], Fresh[9228], Fresh[9227], Fresh[9226], Fresh[9225]}), .outt ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, n2304}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2466 ( .ina ({new_AGEMA_signal_19951, new_AGEMA_signal_19949, new_AGEMA_signal_19947, new_AGEMA_signal_19945, new_AGEMA_signal_19943}), .inb ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, n2292}), .clk ( clk ), .rnd ({Fresh[9254], Fresh[9253], Fresh[9252], Fresh[9251], Fresh[9250], Fresh[9249], Fresh[9248], Fresh[9247], Fresh[9246], Fresh[9245], Fresh[9244], Fresh[9243], Fresh[9242], Fresh[9241], Fresh[9240]}), .outt ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2295}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2488 ( .ina ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, n2321}), .inb ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n2320}), .clk ( clk ), .rnd ({Fresh[9269], Fresh[9268], Fresh[9267], Fresh[9266], Fresh[9265], Fresh[9264], Fresh[9263], Fresh[9262], Fresh[9261], Fresh[9260], Fresh[9259], Fresh[9258], Fresh[9257], Fresh[9256], Fresh[9255]}), .outt ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, n2322}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2499 ( .ina ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, n2332}), .inb ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2331}), .clk ( clk ), .rnd ({Fresh[9284], Fresh[9283], Fresh[9282], Fresh[9281], Fresh[9280], Fresh[9279], Fresh[9278], Fresh[9277], Fresh[9276], Fresh[9275], Fresh[9274], Fresh[9273], Fresh[9272], Fresh[9271], Fresh[9270]}), .outt ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, n2333}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2509 ( .ina ({new_AGEMA_signal_19971, new_AGEMA_signal_19967, new_AGEMA_signal_19963, new_AGEMA_signal_19959, new_AGEMA_signal_19955}), .inb ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, n2342}), .clk ( clk ), .rnd ({Fresh[9299], Fresh[9298], Fresh[9297], Fresh[9296], Fresh[9295], Fresh[9294], Fresh[9293], Fresh[9292], Fresh[9291], Fresh[9290], Fresh[9289], Fresh[9288], Fresh[9287], Fresh[9286], Fresh[9285]}), .outt ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, n2345}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2526 ( .ina ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2358}), .inb ({new_AGEMA_signal_19981, new_AGEMA_signal_19979, new_AGEMA_signal_19977, new_AGEMA_signal_19975, new_AGEMA_signal_19973}), .clk ( clk ), .rnd ({Fresh[9314], Fresh[9313], Fresh[9312], Fresh[9311], Fresh[9310], Fresh[9309], Fresh[9308], Fresh[9307], Fresh[9306], Fresh[9305], Fresh[9304], Fresh[9303], Fresh[9302], Fresh[9301], Fresh[9300]}), .outt ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, new_AGEMA_signal_3686, n2361}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2549 ( .ina ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, n2387}), .inb ({new_AGEMA_signal_19991, new_AGEMA_signal_19989, new_AGEMA_signal_19987, new_AGEMA_signal_19985, new_AGEMA_signal_19983}), .clk ( clk ), .rnd ({Fresh[9329], Fresh[9328], Fresh[9327], Fresh[9326], Fresh[9325], Fresh[9324], Fresh[9323], Fresh[9322], Fresh[9321], Fresh[9320], Fresh[9319], Fresh[9318], Fresh[9317], Fresh[9316], Fresh[9315]}), .outt ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, new_AGEMA_signal_3338, n2388}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2556 ( .ina ({new_AGEMA_signal_20011, new_AGEMA_signal_20007, new_AGEMA_signal_20003, new_AGEMA_signal_19999, new_AGEMA_signal_19995}), .inb ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2392}), .clk ( clk ), .rnd ({Fresh[9344], Fresh[9343], Fresh[9342], Fresh[9341], Fresh[9340], Fresh[9339], Fresh[9338], Fresh[9337], Fresh[9336], Fresh[9335], Fresh[9334], Fresh[9333], Fresh[9332], Fresh[9331], Fresh[9330]}), .outt ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, n2393}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2567 ( .ina ({new_AGEMA_signal_20031, new_AGEMA_signal_20027, new_AGEMA_signal_20023, new_AGEMA_signal_20019, new_AGEMA_signal_20015}), .inb ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2404}), .clk ( clk ), .rnd ({Fresh[9359], Fresh[9358], Fresh[9357], Fresh[9356], Fresh[9355], Fresh[9354], Fresh[9353], Fresh[9352], Fresh[9351], Fresh[9350], Fresh[9349], Fresh[9348], Fresh[9347], Fresh[9346], Fresh[9345]}), .outt ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, n2405}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2571 ( .ina ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, n2409}), .inb ({new_AGEMA_signal_20051, new_AGEMA_signal_20047, new_AGEMA_signal_20043, new_AGEMA_signal_20039, new_AGEMA_signal_20035}), .clk ( clk ), .rnd ({Fresh[9374], Fresh[9373], Fresh[9372], Fresh[9371], Fresh[9370], Fresh[9369], Fresh[9368], Fresh[9367], Fresh[9366], Fresh[9365], Fresh[9364], Fresh[9363], Fresh[9362], Fresh[9361], Fresh[9360]}), .outt ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, n2410}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2576 ( .ina ({new_AGEMA_signal_20071, new_AGEMA_signal_20067, new_AGEMA_signal_20063, new_AGEMA_signal_20059, new_AGEMA_signal_20055}), .inb ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2414}), .clk ( clk ), .rnd ({Fresh[9389], Fresh[9388], Fresh[9387], Fresh[9386], Fresh[9385], Fresh[9384], Fresh[9383], Fresh[9382], Fresh[9381], Fresh[9380], Fresh[9379], Fresh[9378], Fresh[9377], Fresh[9376], Fresh[9375]}), .outt ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, n2421}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2579 ( .ina ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2418}), .inb ({new_AGEMA_signal_20091, new_AGEMA_signal_20087, new_AGEMA_signal_20083, new_AGEMA_signal_20079, new_AGEMA_signal_20075}), .clk ( clk ), .rnd ({Fresh[9404], Fresh[9403], Fresh[9402], Fresh[9401], Fresh[9400], Fresh[9399], Fresh[9398], Fresh[9397], Fresh[9396], Fresh[9395], Fresh[9394], Fresh[9393], Fresh[9392], Fresh[9391], Fresh[9390]}), .outt ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, n2419}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2590 ( .ina ({new_AGEMA_signal_20101, new_AGEMA_signal_20099, new_AGEMA_signal_20097, new_AGEMA_signal_20095, new_AGEMA_signal_20093}), .inb ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, new_AGEMA_signal_3362, n2432}), .clk ( clk ), .rnd ({Fresh[9419], Fresh[9418], Fresh[9417], Fresh[9416], Fresh[9415], Fresh[9414], Fresh[9413], Fresh[9412], Fresh[9411], Fresh[9410], Fresh[9409], Fresh[9408], Fresh[9407], Fresh[9406], Fresh[9405]}), .outt ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2436}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2604 ( .ina ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2449}), .inb ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, n2448}), .clk ( clk ), .rnd ({Fresh[9434], Fresh[9433], Fresh[9432], Fresh[9431], Fresh[9430], Fresh[9429], Fresh[9428], Fresh[9427], Fresh[9426], Fresh[9425], Fresh[9424], Fresh[9423], Fresh[9422], Fresh[9421], Fresh[9420]}), .outt ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, new_AGEMA_signal_3719, new_AGEMA_signal_3718, n2450}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2610 ( .ina ({new_AGEMA_signal_20111, new_AGEMA_signal_20109, new_AGEMA_signal_20107, new_AGEMA_signal_20105, new_AGEMA_signal_20103}), .inb ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, n2455}), .clk ( clk ), .rnd ({Fresh[9449], Fresh[9448], Fresh[9447], Fresh[9446], Fresh[9445], Fresh[9444], Fresh[9443], Fresh[9442], Fresh[9441], Fresh[9440], Fresh[9439], Fresh[9438], Fresh[9437], Fresh[9436], Fresh[9435]}), .outt ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723, new_AGEMA_signal_3722, n2456}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2613 ( .ina ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2460}), .inb ({new_AGEMA_signal_20121, new_AGEMA_signal_20119, new_AGEMA_signal_20117, new_AGEMA_signal_20115, new_AGEMA_signal_20113}), .clk ( clk ), .rnd ({Fresh[9464], Fresh[9463], Fresh[9462], Fresh[9461], Fresh[9460], Fresh[9459], Fresh[9458], Fresh[9457], Fresh[9456], Fresh[9455], Fresh[9454], Fresh[9453], Fresh[9452], Fresh[9451], Fresh[9450]}), .outt ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, n2461}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2619 ( .ina ({new_AGEMA_signal_20131, new_AGEMA_signal_20129, new_AGEMA_signal_20127, new_AGEMA_signal_20125, new_AGEMA_signal_20123}), .inb ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2466}), .clk ( clk ), .rnd ({Fresh[9479], Fresh[9478], Fresh[9477], Fresh[9476], Fresh[9475], Fresh[9474], Fresh[9473], Fresh[9472], Fresh[9471], Fresh[9470], Fresh[9469], Fresh[9468], Fresh[9467], Fresh[9466], Fresh[9465]}), .outt ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, n2469}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2630 ( .ina ({new_AGEMA_signal_20151, new_AGEMA_signal_20147, new_AGEMA_signal_20143, new_AGEMA_signal_20139, new_AGEMA_signal_20135}), .inb ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, n2477}), .clk ( clk ), .rnd ({Fresh[9494], Fresh[9493], Fresh[9492], Fresh[9491], Fresh[9490], Fresh[9489], Fresh[9488], Fresh[9487], Fresh[9486], Fresh[9485], Fresh[9484], Fresh[9483], Fresh[9482], Fresh[9481], Fresh[9480]}), .outt ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, n2478}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2635 ( .ina ({new_AGEMA_signal_20171, new_AGEMA_signal_20167, new_AGEMA_signal_20163, new_AGEMA_signal_20159, new_AGEMA_signal_20155}), .inb ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2482}), .clk ( clk ), .rnd ({Fresh[9509], Fresh[9508], Fresh[9507], Fresh[9506], Fresh[9505], Fresh[9504], Fresh[9503], Fresh[9502], Fresh[9501], Fresh[9500], Fresh[9499], Fresh[9498], Fresh[9497], Fresh[9496], Fresh[9495]}), .outt ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, n2484}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2643 ( .ina ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n2490}), .inb ({new_AGEMA_signal_20181, new_AGEMA_signal_20179, new_AGEMA_signal_20177, new_AGEMA_signal_20175, new_AGEMA_signal_20173}), .clk ( clk ), .rnd ({Fresh[9524], Fresh[9523], Fresh[9522], Fresh[9521], Fresh[9520], Fresh[9519], Fresh[9518], Fresh[9517], Fresh[9516], Fresh[9515], Fresh[9514], Fresh[9513], Fresh[9512], Fresh[9511], Fresh[9510]}), .outt ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, n2491}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2649 ( .ina ({new_AGEMA_signal_20191, new_AGEMA_signal_20189, new_AGEMA_signal_20187, new_AGEMA_signal_20185, new_AGEMA_signal_20183}), .inb ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, n2496}), .clk ( clk ), .rnd ({Fresh[9539], Fresh[9538], Fresh[9537], Fresh[9536], Fresh[9535], Fresh[9534], Fresh[9533], Fresh[9532], Fresh[9531], Fresh[9530], Fresh[9529], Fresh[9528], Fresh[9527], Fresh[9526], Fresh[9525]}), .outt ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, new_AGEMA_signal_3742, n2500}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2656 ( .ina ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, new_AGEMA_signal_3746, n2507}), .inb ({new_AGEMA_signal_20201, new_AGEMA_signal_20199, new_AGEMA_signal_20197, new_AGEMA_signal_20195, new_AGEMA_signal_20193}), .clk ( clk ), .rnd ({Fresh[9554], Fresh[9553], Fresh[9552], Fresh[9551], Fresh[9550], Fresh[9549], Fresh[9548], Fresh[9547], Fresh[9546], Fresh[9545], Fresh[9544], Fresh[9543], Fresh[9542], Fresh[9541], Fresh[9540]}), .outt ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, new_AGEMA_signal_4007, new_AGEMA_signal_4006, n2508}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2670 ( .ina ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, n2525}), .inb ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, n2524}), .clk ( clk ), .rnd ({Fresh[9569], Fresh[9568], Fresh[9567], Fresh[9566], Fresh[9565], Fresh[9564], Fresh[9563], Fresh[9562], Fresh[9561], Fresh[9560], Fresh[9559], Fresh[9558], Fresh[9557], Fresh[9556], Fresh[9555]}), .outt ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, new_AGEMA_signal_4010, n2526}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2679 ( .ina ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2537}), .inb ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, n2536}), .clk ( clk ), .rnd ({Fresh[9584], Fresh[9583], Fresh[9582], Fresh[9581], Fresh[9580], Fresh[9579], Fresh[9578], Fresh[9577], Fresh[9576], Fresh[9575], Fresh[9574], Fresh[9573], Fresh[9572], Fresh[9571], Fresh[9570]}), .outt ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, new_AGEMA_signal_3755, new_AGEMA_signal_3754, n2539}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2682 ( .ina ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2543}), .inb ({new_AGEMA_signal_20211, new_AGEMA_signal_20209, new_AGEMA_signal_20207, new_AGEMA_signal_20205, new_AGEMA_signal_20203}), .clk ( clk ), .rnd ({Fresh[9599], Fresh[9598], Fresh[9597], Fresh[9596], Fresh[9595], Fresh[9594], Fresh[9593], Fresh[9592], Fresh[9591], Fresh[9590], Fresh[9589], Fresh[9588], Fresh[9587], Fresh[9586], Fresh[9585]}), .outt ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, new_AGEMA_signal_3758, n2548}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2694 ( .ina ({new_AGEMA_signal_20221, new_AGEMA_signal_20219, new_AGEMA_signal_20217, new_AGEMA_signal_20215, new_AGEMA_signal_20213}), .inb ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, n2557}), .clk ( clk ), .rnd ({Fresh[9614], Fresh[9613], Fresh[9612], Fresh[9611], Fresh[9610], Fresh[9609], Fresh[9608], Fresh[9607], Fresh[9606], Fresh[9605], Fresh[9604], Fresh[9603], Fresh[9602], Fresh[9601], Fresh[9600]}), .outt ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, n2568}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2700 ( .ina ({new_AGEMA_signal_20231, new_AGEMA_signal_20229, new_AGEMA_signal_20227, new_AGEMA_signal_20225, new_AGEMA_signal_20223}), .inb ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n2565}), .clk ( clk ), .rnd ({Fresh[9629], Fresh[9628], Fresh[9627], Fresh[9626], Fresh[9625], Fresh[9624], Fresh[9623], Fresh[9622], Fresh[9621], Fresh[9620], Fresh[9619], Fresh[9618], Fresh[9617], Fresh[9616], Fresh[9615]}), .outt ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, new_AGEMA_signal_3767, new_AGEMA_signal_3766, n2567}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2710 ( .ina ({new_AGEMA_signal_20241, new_AGEMA_signal_20239, new_AGEMA_signal_20237, new_AGEMA_signal_20235, new_AGEMA_signal_20233}), .inb ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, n2580}), .clk ( clk ), .rnd ({Fresh[9644], Fresh[9643], Fresh[9642], Fresh[9641], Fresh[9640], Fresh[9639], Fresh[9638], Fresh[9637], Fresh[9636], Fresh[9635], Fresh[9634], Fresh[9633], Fresh[9632], Fresh[9631], Fresh[9630]}), .outt ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, n2583}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2728 ( .ina ({new_AGEMA_signal_20251, new_AGEMA_signal_20249, new_AGEMA_signal_20247, new_AGEMA_signal_20245, new_AGEMA_signal_20243}), .inb ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, n2602}), .clk ( clk ), .rnd ({Fresh[9659], Fresh[9658], Fresh[9657], Fresh[9656], Fresh[9655], Fresh[9654], Fresh[9653], Fresh[9652], Fresh[9651], Fresh[9650], Fresh[9649], Fresh[9648], Fresh[9647], Fresh[9646], Fresh[9645]}), .outt ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2604}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2739 ( .ina ({new_AGEMA_signal_20261, new_AGEMA_signal_20259, new_AGEMA_signal_20257, new_AGEMA_signal_20255, new_AGEMA_signal_20253}), .inb ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, n2619}), .clk ( clk ), .rnd ({Fresh[9674], Fresh[9673], Fresh[9672], Fresh[9671], Fresh[9670], Fresh[9669], Fresh[9668], Fresh[9667], Fresh[9666], Fresh[9665], Fresh[9664], Fresh[9663], Fresh[9662], Fresh[9661], Fresh[9660]}), .outt ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, new_AGEMA_signal_3778, n2621}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2745 ( .ina ({new_AGEMA_signal_20281, new_AGEMA_signal_20277, new_AGEMA_signal_20273, new_AGEMA_signal_20269, new_AGEMA_signal_20265}), .inb ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, n2628}), .clk ( clk ), .rnd ({Fresh[9689], Fresh[9688], Fresh[9687], Fresh[9686], Fresh[9685], Fresh[9684], Fresh[9683], Fresh[9682], Fresh[9681], Fresh[9680], Fresh[9679], Fresh[9678], Fresh[9677], Fresh[9676], Fresh[9675]}), .outt ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, new_AGEMA_signal_3783, new_AGEMA_signal_3782, n2633}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2756 ( .ina ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2649}), .inb ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, n2648}), .clk ( clk ), .rnd ({Fresh[9704], Fresh[9703], Fresh[9702], Fresh[9701], Fresh[9700], Fresh[9699], Fresh[9698], Fresh[9697], Fresh[9696], Fresh[9695], Fresh[9694], Fresh[9693], Fresh[9692], Fresh[9691], Fresh[9690]}), .outt ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786, n2660}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2759 ( .ina ({new_AGEMA_signal_20291, new_AGEMA_signal_20289, new_AGEMA_signal_20287, new_AGEMA_signal_20285, new_AGEMA_signal_20283}), .inb ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, new_AGEMA_signal_3158, n2652}), .clk ( clk ), .rnd ({Fresh[9719], Fresh[9718], Fresh[9717], Fresh[9716], Fresh[9715], Fresh[9714], Fresh[9713], Fresh[9712], Fresh[9711], Fresh[9710], Fresh[9709], Fresh[9708], Fresh[9707], Fresh[9706], Fresh[9705]}), .outt ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_3791, new_AGEMA_signal_3790, n2656}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2766 ( .ina ({new_AGEMA_signal_20301, new_AGEMA_signal_20299, new_AGEMA_signal_20297, new_AGEMA_signal_20295, new_AGEMA_signal_20293}), .inb ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, n2664}), .clk ( clk ), .rnd ({Fresh[9734], Fresh[9733], Fresh[9732], Fresh[9731], Fresh[9730], Fresh[9729], Fresh[9728], Fresh[9727], Fresh[9726], Fresh[9725], Fresh[9724], Fresh[9723], Fresh[9722], Fresh[9721], Fresh[9720]}), .outt ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, new_AGEMA_signal_3795, new_AGEMA_signal_3794, n2666}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2774 ( .ina ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, n2681}), .inb ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, n2680}), .clk ( clk ), .rnd ({Fresh[9749], Fresh[9748], Fresh[9747], Fresh[9746], Fresh[9745], Fresh[9744], Fresh[9743], Fresh[9742], Fresh[9741], Fresh[9740], Fresh[9739], Fresh[9738], Fresh[9737], Fresh[9736], Fresh[9735]}), .outt ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, new_AGEMA_signal_3799, new_AGEMA_signal_3798, n2706}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2777 ( .ina ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, n2686}), .inb ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2685}), .clk ( clk ), .rnd ({Fresh[9764], Fresh[9763], Fresh[9762], Fresh[9761], Fresh[9760], Fresh[9759], Fresh[9758], Fresh[9757], Fresh[9756], Fresh[9755], Fresh[9754], Fresh[9753], Fresh[9752], Fresh[9751], Fresh[9750]}), .outt ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, new_AGEMA_signal_3803, new_AGEMA_signal_3802, n2704}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2781 ( .ina ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, n2692}), .inb ({new_AGEMA_signal_20311, new_AGEMA_signal_20309, new_AGEMA_signal_20307, new_AGEMA_signal_20305, new_AGEMA_signal_20303}), .clk ( clk ), .rnd ({Fresh[9779], Fresh[9778], Fresh[9777], Fresh[9776], Fresh[9775], Fresh[9774], Fresh[9773], Fresh[9772], Fresh[9771], Fresh[9770], Fresh[9769], Fresh[9768], Fresh[9767], Fresh[9766], Fresh[9765]}), .outt ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, n2696}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2794 ( .ina ({new_AGEMA_signal_20321, new_AGEMA_signal_20319, new_AGEMA_signal_20317, new_AGEMA_signal_20315, new_AGEMA_signal_20313}), .inb ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2716}), .clk ( clk ), .rnd ({Fresh[9794], Fresh[9793], Fresh[9792], Fresh[9791], Fresh[9790], Fresh[9789], Fresh[9788], Fresh[9787], Fresh[9786], Fresh[9785], Fresh[9784], Fresh[9783], Fresh[9782], Fresh[9781], Fresh[9780]}), .outt ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, n2718}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2801 ( .ina ({new_AGEMA_signal_20331, new_AGEMA_signal_20329, new_AGEMA_signal_20327, new_AGEMA_signal_20325, new_AGEMA_signal_20323}), .inb ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, n2728}), .clk ( clk ), .rnd ({Fresh[9809], Fresh[9808], Fresh[9807], Fresh[9806], Fresh[9805], Fresh[9804], Fresh[9803], Fresh[9802], Fresh[9801], Fresh[9800], Fresh[9799], Fresh[9798], Fresh[9797], Fresh[9796], Fresh[9795]}), .outt ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, new_AGEMA_signal_3814, n2730}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2805 ( .ina ({new_AGEMA_signal_20351, new_AGEMA_signal_20347, new_AGEMA_signal_20343, new_AGEMA_signal_20339, new_AGEMA_signal_20335}), .inb ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, n2735}), .clk ( clk ), .rnd ({Fresh[9824], Fresh[9823], Fresh[9822], Fresh[9821], Fresh[9820], Fresh[9819], Fresh[9818], Fresh[9817], Fresh[9816], Fresh[9815], Fresh[9814], Fresh[9813], Fresh[9812], Fresh[9811], Fresh[9810]}), .outt ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, new_AGEMA_signal_3819, new_AGEMA_signal_3818, n2745}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2809 ( .ina ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2743}), .inb ({new_AGEMA_signal_20371, new_AGEMA_signal_20367, new_AGEMA_signal_20363, new_AGEMA_signal_20359, new_AGEMA_signal_20355}), .clk ( clk ), .rnd ({Fresh[9839], Fresh[9838], Fresh[9837], Fresh[9836], Fresh[9835], Fresh[9834], Fresh[9833], Fresh[9832], Fresh[9831], Fresh[9830], Fresh[9829], Fresh[9828], Fresh[9827], Fresh[9826], Fresh[9825]}), .outt ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, n2744}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2814 ( .ina ({new_AGEMA_signal_19931, new_AGEMA_signal_19929, new_AGEMA_signal_19927, new_AGEMA_signal_19925, new_AGEMA_signal_19923}), .inb ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, n2751}), .clk ( clk ), .rnd ({Fresh[9854], Fresh[9853], Fresh[9852], Fresh[9851], Fresh[9850], Fresh[9849], Fresh[9848], Fresh[9847], Fresh[9846], Fresh[9845], Fresh[9844], Fresh[9843], Fresh[9842], Fresh[9841], Fresh[9840]}), .outt ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, new_AGEMA_signal_3827, new_AGEMA_signal_3826, n2759}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2821 ( .ina ({new_AGEMA_signal_20391, new_AGEMA_signal_20387, new_AGEMA_signal_20383, new_AGEMA_signal_20379, new_AGEMA_signal_20375}), .inb ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, n2764}), .clk ( clk ), .rnd ({Fresh[9869], Fresh[9868], Fresh[9867], Fresh[9866], Fresh[9865], Fresh[9864], Fresh[9863], Fresh[9862], Fresh[9861], Fresh[9860], Fresh[9859], Fresh[9858], Fresh[9857], Fresh[9856], Fresh[9855]}), .outt ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, new_AGEMA_signal_3831, new_AGEMA_signal_3830, n2771}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2833 ( .ina ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, new_AGEMA_signal_3038, n2788}), .inb ({new_AGEMA_signal_20411, new_AGEMA_signal_20407, new_AGEMA_signal_20403, new_AGEMA_signal_20399, new_AGEMA_signal_20395}), .clk ( clk ), .rnd ({Fresh[9884], Fresh[9883], Fresh[9882], Fresh[9881], Fresh[9880], Fresh[9879], Fresh[9878], Fresh[9877], Fresh[9876], Fresh[9875], Fresh[9874], Fresh[9873], Fresh[9872], Fresh[9871], Fresh[9870]}), .outt ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, n2798}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2850 ( .ina ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2822}), .inb ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, n2821}), .clk ( clk ), .rnd ({Fresh[9899], Fresh[9898], Fresh[9897], Fresh[9896], Fresh[9895], Fresh[9894], Fresh[9893], Fresh[9892], Fresh[9891], Fresh[9890], Fresh[9889], Fresh[9888], Fresh[9887], Fresh[9886], Fresh[9885]}), .outt ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, new_AGEMA_signal_3839, new_AGEMA_signal_3838, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C ( clk ), .D ( new_AGEMA_signal_20414 ), .Q ( new_AGEMA_signal_20415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C ( clk ), .D ( new_AGEMA_signal_20418 ), .Q ( new_AGEMA_signal_20419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C ( clk ), .D ( new_AGEMA_signal_20422 ), .Q ( new_AGEMA_signal_20423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C ( clk ), .D ( new_AGEMA_signal_20426 ), .Q ( new_AGEMA_signal_20427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C ( clk ), .D ( new_AGEMA_signal_20430 ), .Q ( new_AGEMA_signal_20431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C ( clk ), .D ( new_AGEMA_signal_20434 ), .Q ( new_AGEMA_signal_20435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C ( clk ), .D ( new_AGEMA_signal_20438 ), .Q ( new_AGEMA_signal_20439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C ( clk ), .D ( new_AGEMA_signal_20442 ), .Q ( new_AGEMA_signal_20443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C ( clk ), .D ( new_AGEMA_signal_20446 ), .Q ( new_AGEMA_signal_20447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C ( clk ), .D ( new_AGEMA_signal_20450 ), .Q ( new_AGEMA_signal_20451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C ( clk ), .D ( new_AGEMA_signal_20458 ), .Q ( new_AGEMA_signal_20459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C ( clk ), .D ( new_AGEMA_signal_20466 ), .Q ( new_AGEMA_signal_20467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C ( clk ), .D ( new_AGEMA_signal_20474 ), .Q ( new_AGEMA_signal_20475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C ( clk ), .D ( new_AGEMA_signal_20482 ), .Q ( new_AGEMA_signal_20483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C ( clk ), .D ( new_AGEMA_signal_20490 ), .Q ( new_AGEMA_signal_20491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C ( clk ), .D ( new_AGEMA_signal_20492 ), .Q ( new_AGEMA_signal_20493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C ( clk ), .D ( new_AGEMA_signal_20494 ), .Q ( new_AGEMA_signal_20495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C ( clk ), .D ( new_AGEMA_signal_20496 ), .Q ( new_AGEMA_signal_20497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C ( clk ), .D ( new_AGEMA_signal_20498 ), .Q ( new_AGEMA_signal_20499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C ( clk ), .D ( new_AGEMA_signal_20500 ), .Q ( new_AGEMA_signal_20501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C ( clk ), .D ( new_AGEMA_signal_20508 ), .Q ( new_AGEMA_signal_20509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C ( clk ), .D ( new_AGEMA_signal_20516 ), .Q ( new_AGEMA_signal_20517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C ( clk ), .D ( new_AGEMA_signal_20524 ), .Q ( new_AGEMA_signal_20525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C ( clk ), .D ( new_AGEMA_signal_20532 ), .Q ( new_AGEMA_signal_20533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C ( clk ), .D ( new_AGEMA_signal_20540 ), .Q ( new_AGEMA_signal_20541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C ( clk ), .D ( new_AGEMA_signal_20546 ), .Q ( new_AGEMA_signal_20547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C ( clk ), .D ( new_AGEMA_signal_20552 ), .Q ( new_AGEMA_signal_20553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C ( clk ), .D ( new_AGEMA_signal_20558 ), .Q ( new_AGEMA_signal_20559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C ( clk ), .D ( new_AGEMA_signal_20564 ), .Q ( new_AGEMA_signal_20565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C ( clk ), .D ( new_AGEMA_signal_20570 ), .Q ( new_AGEMA_signal_20571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C ( clk ), .D ( new_AGEMA_signal_20574 ), .Q ( new_AGEMA_signal_20575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C ( clk ), .D ( new_AGEMA_signal_20578 ), .Q ( new_AGEMA_signal_20579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C ( clk ), .D ( new_AGEMA_signal_20582 ), .Q ( new_AGEMA_signal_20583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C ( clk ), .D ( new_AGEMA_signal_20586 ), .Q ( new_AGEMA_signal_20587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C ( clk ), .D ( new_AGEMA_signal_20590 ), .Q ( new_AGEMA_signal_20591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C ( clk ), .D ( new_AGEMA_signal_20596 ), .Q ( new_AGEMA_signal_20597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C ( clk ), .D ( new_AGEMA_signal_20602 ), .Q ( new_AGEMA_signal_20603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C ( clk ), .D ( new_AGEMA_signal_20608 ), .Q ( new_AGEMA_signal_20609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C ( clk ), .D ( new_AGEMA_signal_20614 ), .Q ( new_AGEMA_signal_20615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C ( clk ), .D ( new_AGEMA_signal_20620 ), .Q ( new_AGEMA_signal_20621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C ( clk ), .D ( new_AGEMA_signal_20622 ), .Q ( new_AGEMA_signal_20623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C ( clk ), .D ( new_AGEMA_signal_20624 ), .Q ( new_AGEMA_signal_20625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C ( clk ), .D ( new_AGEMA_signal_20626 ), .Q ( new_AGEMA_signal_20627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C ( clk ), .D ( new_AGEMA_signal_20628 ), .Q ( new_AGEMA_signal_20629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C ( clk ), .D ( new_AGEMA_signal_20630 ), .Q ( new_AGEMA_signal_20631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C ( clk ), .D ( new_AGEMA_signal_20636 ), .Q ( new_AGEMA_signal_20637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C ( clk ), .D ( new_AGEMA_signal_20642 ), .Q ( new_AGEMA_signal_20643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C ( clk ), .D ( new_AGEMA_signal_20648 ), .Q ( new_AGEMA_signal_20649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C ( clk ), .D ( new_AGEMA_signal_20654 ), .Q ( new_AGEMA_signal_20655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C ( clk ), .D ( new_AGEMA_signal_20660 ), .Q ( new_AGEMA_signal_20661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C ( clk ), .D ( new_AGEMA_signal_20666 ), .Q ( new_AGEMA_signal_20667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C ( clk ), .D ( new_AGEMA_signal_20672 ), .Q ( new_AGEMA_signal_20673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C ( clk ), .D ( new_AGEMA_signal_20678 ), .Q ( new_AGEMA_signal_20679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C ( clk ), .D ( new_AGEMA_signal_20684 ), .Q ( new_AGEMA_signal_20685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C ( clk ), .D ( new_AGEMA_signal_20690 ), .Q ( new_AGEMA_signal_20691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C ( clk ), .D ( new_AGEMA_signal_20692 ), .Q ( new_AGEMA_signal_20693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C ( clk ), .D ( new_AGEMA_signal_20694 ), .Q ( new_AGEMA_signal_20695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C ( clk ), .D ( new_AGEMA_signal_20696 ), .Q ( new_AGEMA_signal_20697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C ( clk ), .D ( new_AGEMA_signal_20698 ), .Q ( new_AGEMA_signal_20699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C ( clk ), .D ( new_AGEMA_signal_20700 ), .Q ( new_AGEMA_signal_20701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C ( clk ), .D ( new_AGEMA_signal_20704 ), .Q ( new_AGEMA_signal_20705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C ( clk ), .D ( new_AGEMA_signal_20708 ), .Q ( new_AGEMA_signal_20709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C ( clk ), .D ( new_AGEMA_signal_20712 ), .Q ( new_AGEMA_signal_20713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C ( clk ), .D ( new_AGEMA_signal_20716 ), .Q ( new_AGEMA_signal_20717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C ( clk ), .D ( new_AGEMA_signal_20720 ), .Q ( new_AGEMA_signal_20721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C ( clk ), .D ( new_AGEMA_signal_20726 ), .Q ( new_AGEMA_signal_20727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C ( clk ), .D ( new_AGEMA_signal_20732 ), .Q ( new_AGEMA_signal_20733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C ( clk ), .D ( new_AGEMA_signal_20738 ), .Q ( new_AGEMA_signal_20739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C ( clk ), .D ( new_AGEMA_signal_20744 ), .Q ( new_AGEMA_signal_20745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C ( clk ), .D ( new_AGEMA_signal_20750 ), .Q ( new_AGEMA_signal_20751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C ( clk ), .D ( new_AGEMA_signal_20756 ), .Q ( new_AGEMA_signal_20757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C ( clk ), .D ( new_AGEMA_signal_20762 ), .Q ( new_AGEMA_signal_20763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C ( clk ), .D ( new_AGEMA_signal_20768 ), .Q ( new_AGEMA_signal_20769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C ( clk ), .D ( new_AGEMA_signal_20774 ), .Q ( new_AGEMA_signal_20775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C ( clk ), .D ( new_AGEMA_signal_20780 ), .Q ( new_AGEMA_signal_20781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C ( clk ), .D ( new_AGEMA_signal_20782 ), .Q ( new_AGEMA_signal_20783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C ( clk ), .D ( new_AGEMA_signal_20784 ), .Q ( new_AGEMA_signal_20785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C ( clk ), .D ( new_AGEMA_signal_20786 ), .Q ( new_AGEMA_signal_20787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C ( clk ), .D ( new_AGEMA_signal_20788 ), .Q ( new_AGEMA_signal_20789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C ( clk ), .D ( new_AGEMA_signal_20790 ), .Q ( new_AGEMA_signal_20791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C ( clk ), .D ( new_AGEMA_signal_20796 ), .Q ( new_AGEMA_signal_20797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C ( clk ), .D ( new_AGEMA_signal_20802 ), .Q ( new_AGEMA_signal_20803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C ( clk ), .D ( new_AGEMA_signal_20808 ), .Q ( new_AGEMA_signal_20809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C ( clk ), .D ( new_AGEMA_signal_20814 ), .Q ( new_AGEMA_signal_20815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C ( clk ), .D ( new_AGEMA_signal_20820 ), .Q ( new_AGEMA_signal_20821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C ( clk ), .D ( new_AGEMA_signal_20822 ), .Q ( new_AGEMA_signal_20823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C ( clk ), .D ( new_AGEMA_signal_20824 ), .Q ( new_AGEMA_signal_20825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C ( clk ), .D ( new_AGEMA_signal_20826 ), .Q ( new_AGEMA_signal_20827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C ( clk ), .D ( new_AGEMA_signal_20828 ), .Q ( new_AGEMA_signal_20829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C ( clk ), .D ( new_AGEMA_signal_20830 ), .Q ( new_AGEMA_signal_20831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C ( clk ), .D ( new_AGEMA_signal_20834 ), .Q ( new_AGEMA_signal_20835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C ( clk ), .D ( new_AGEMA_signal_20838 ), .Q ( new_AGEMA_signal_20839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C ( clk ), .D ( new_AGEMA_signal_20842 ), .Q ( new_AGEMA_signal_20843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C ( clk ), .D ( new_AGEMA_signal_20846 ), .Q ( new_AGEMA_signal_20847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C ( clk ), .D ( new_AGEMA_signal_20850 ), .Q ( new_AGEMA_signal_20851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C ( clk ), .D ( new_AGEMA_signal_20854 ), .Q ( new_AGEMA_signal_20855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C ( clk ), .D ( new_AGEMA_signal_20858 ), .Q ( new_AGEMA_signal_20859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C ( clk ), .D ( new_AGEMA_signal_20862 ), .Q ( new_AGEMA_signal_20863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C ( clk ), .D ( new_AGEMA_signal_20866 ), .Q ( new_AGEMA_signal_20867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C ( clk ), .D ( new_AGEMA_signal_20870 ), .Q ( new_AGEMA_signal_20871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C ( clk ), .D ( new_AGEMA_signal_20872 ), .Q ( new_AGEMA_signal_20873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C ( clk ), .D ( new_AGEMA_signal_20874 ), .Q ( new_AGEMA_signal_20875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C ( clk ), .D ( new_AGEMA_signal_20876 ), .Q ( new_AGEMA_signal_20877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C ( clk ), .D ( new_AGEMA_signal_20878 ), .Q ( new_AGEMA_signal_20879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C ( clk ), .D ( new_AGEMA_signal_20880 ), .Q ( new_AGEMA_signal_20881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C ( clk ), .D ( new_AGEMA_signal_20888 ), .Q ( new_AGEMA_signal_20889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C ( clk ), .D ( new_AGEMA_signal_20896 ), .Q ( new_AGEMA_signal_20897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C ( clk ), .D ( new_AGEMA_signal_20904 ), .Q ( new_AGEMA_signal_20905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C ( clk ), .D ( new_AGEMA_signal_20912 ), .Q ( new_AGEMA_signal_20913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C ( clk ), .D ( new_AGEMA_signal_20920 ), .Q ( new_AGEMA_signal_20921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C ( clk ), .D ( new_AGEMA_signal_20926 ), .Q ( new_AGEMA_signal_20927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C ( clk ), .D ( new_AGEMA_signal_20932 ), .Q ( new_AGEMA_signal_20933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C ( clk ), .D ( new_AGEMA_signal_20938 ), .Q ( new_AGEMA_signal_20939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C ( clk ), .D ( new_AGEMA_signal_20944 ), .Q ( new_AGEMA_signal_20945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C ( clk ), .D ( new_AGEMA_signal_20950 ), .Q ( new_AGEMA_signal_20951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C ( clk ), .D ( new_AGEMA_signal_20954 ), .Q ( new_AGEMA_signal_20955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C ( clk ), .D ( new_AGEMA_signal_20958 ), .Q ( new_AGEMA_signal_20959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C ( clk ), .D ( new_AGEMA_signal_20962 ), .Q ( new_AGEMA_signal_20963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C ( clk ), .D ( new_AGEMA_signal_20966 ), .Q ( new_AGEMA_signal_20967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C ( clk ), .D ( new_AGEMA_signal_20970 ), .Q ( new_AGEMA_signal_20971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C ( clk ), .D ( new_AGEMA_signal_20974 ), .Q ( new_AGEMA_signal_20975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C ( clk ), .D ( new_AGEMA_signal_20978 ), .Q ( new_AGEMA_signal_20979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C ( clk ), .D ( new_AGEMA_signal_20982 ), .Q ( new_AGEMA_signal_20983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C ( clk ), .D ( new_AGEMA_signal_20986 ), .Q ( new_AGEMA_signal_20987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C ( clk ), .D ( new_AGEMA_signal_20990 ), .Q ( new_AGEMA_signal_20991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C ( clk ), .D ( new_AGEMA_signal_20992 ), .Q ( new_AGEMA_signal_20993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C ( clk ), .D ( new_AGEMA_signal_20994 ), .Q ( new_AGEMA_signal_20995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C ( clk ), .D ( new_AGEMA_signal_20996 ), .Q ( new_AGEMA_signal_20997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C ( clk ), .D ( new_AGEMA_signal_20998 ), .Q ( new_AGEMA_signal_20999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C ( clk ), .D ( new_AGEMA_signal_21000 ), .Q ( new_AGEMA_signal_21001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C ( clk ), .D ( new_AGEMA_signal_21002 ), .Q ( new_AGEMA_signal_21003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C ( clk ), .D ( new_AGEMA_signal_21004 ), .Q ( new_AGEMA_signal_21005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C ( clk ), .D ( new_AGEMA_signal_21006 ), .Q ( new_AGEMA_signal_21007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C ( clk ), .D ( new_AGEMA_signal_21008 ), .Q ( new_AGEMA_signal_21009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C ( clk ), .D ( new_AGEMA_signal_21010 ), .Q ( new_AGEMA_signal_21011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C ( clk ), .D ( new_AGEMA_signal_21014 ), .Q ( new_AGEMA_signal_21015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C ( clk ), .D ( new_AGEMA_signal_21018 ), .Q ( new_AGEMA_signal_21019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C ( clk ), .D ( new_AGEMA_signal_21022 ), .Q ( new_AGEMA_signal_21023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C ( clk ), .D ( new_AGEMA_signal_21026 ), .Q ( new_AGEMA_signal_21027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C ( clk ), .D ( new_AGEMA_signal_21030 ), .Q ( new_AGEMA_signal_21031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C ( clk ), .D ( new_AGEMA_signal_21034 ), .Q ( new_AGEMA_signal_21035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C ( clk ), .D ( new_AGEMA_signal_21038 ), .Q ( new_AGEMA_signal_21039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C ( clk ), .D ( new_AGEMA_signal_21042 ), .Q ( new_AGEMA_signal_21043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C ( clk ), .D ( new_AGEMA_signal_21046 ), .Q ( new_AGEMA_signal_21047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C ( clk ), .D ( new_AGEMA_signal_21050 ), .Q ( new_AGEMA_signal_21051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C ( clk ), .D ( new_AGEMA_signal_21052 ), .Q ( new_AGEMA_signal_21053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C ( clk ), .D ( new_AGEMA_signal_21054 ), .Q ( new_AGEMA_signal_21055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C ( clk ), .D ( new_AGEMA_signal_21056 ), .Q ( new_AGEMA_signal_21057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C ( clk ), .D ( new_AGEMA_signal_21058 ), .Q ( new_AGEMA_signal_21059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C ( clk ), .D ( new_AGEMA_signal_21060 ), .Q ( new_AGEMA_signal_21061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C ( clk ), .D ( new_AGEMA_signal_21066 ), .Q ( new_AGEMA_signal_21067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C ( clk ), .D ( new_AGEMA_signal_21072 ), .Q ( new_AGEMA_signal_21073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C ( clk ), .D ( new_AGEMA_signal_21078 ), .Q ( new_AGEMA_signal_21079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C ( clk ), .D ( new_AGEMA_signal_21084 ), .Q ( new_AGEMA_signal_21085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C ( clk ), .D ( new_AGEMA_signal_21090 ), .Q ( new_AGEMA_signal_21091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C ( clk ), .D ( new_AGEMA_signal_21094 ), .Q ( new_AGEMA_signal_21095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C ( clk ), .D ( new_AGEMA_signal_21098 ), .Q ( new_AGEMA_signal_21099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C ( clk ), .D ( new_AGEMA_signal_21102 ), .Q ( new_AGEMA_signal_21103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C ( clk ), .D ( new_AGEMA_signal_21106 ), .Q ( new_AGEMA_signal_21107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C ( clk ), .D ( new_AGEMA_signal_21110 ), .Q ( new_AGEMA_signal_21111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C ( clk ), .D ( new_AGEMA_signal_21112 ), .Q ( new_AGEMA_signal_21113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C ( clk ), .D ( new_AGEMA_signal_21114 ), .Q ( new_AGEMA_signal_21115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C ( clk ), .D ( new_AGEMA_signal_21116 ), .Q ( new_AGEMA_signal_21117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C ( clk ), .D ( new_AGEMA_signal_21118 ), .Q ( new_AGEMA_signal_21119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C ( clk ), .D ( new_AGEMA_signal_21120 ), .Q ( new_AGEMA_signal_21121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C ( clk ), .D ( new_AGEMA_signal_21124 ), .Q ( new_AGEMA_signal_21125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C ( clk ), .D ( new_AGEMA_signal_21128 ), .Q ( new_AGEMA_signal_21129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C ( clk ), .D ( new_AGEMA_signal_21132 ), .Q ( new_AGEMA_signal_21133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C ( clk ), .D ( new_AGEMA_signal_21136 ), .Q ( new_AGEMA_signal_21137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C ( clk ), .D ( new_AGEMA_signal_21140 ), .Q ( new_AGEMA_signal_21141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C ( clk ), .D ( new_AGEMA_signal_21144 ), .Q ( new_AGEMA_signal_21145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C ( clk ), .D ( new_AGEMA_signal_21148 ), .Q ( new_AGEMA_signal_21149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C ( clk ), .D ( new_AGEMA_signal_21152 ), .Q ( new_AGEMA_signal_21153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C ( clk ), .D ( new_AGEMA_signal_21156 ), .Q ( new_AGEMA_signal_21157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C ( clk ), .D ( new_AGEMA_signal_21160 ), .Q ( new_AGEMA_signal_21161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C ( clk ), .D ( new_AGEMA_signal_21164 ), .Q ( new_AGEMA_signal_21165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C ( clk ), .D ( new_AGEMA_signal_21168 ), .Q ( new_AGEMA_signal_21169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C ( clk ), .D ( new_AGEMA_signal_21172 ), .Q ( new_AGEMA_signal_21173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C ( clk ), .D ( new_AGEMA_signal_21176 ), .Q ( new_AGEMA_signal_21177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C ( clk ), .D ( new_AGEMA_signal_21180 ), .Q ( new_AGEMA_signal_21181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C ( clk ), .D ( new_AGEMA_signal_21182 ), .Q ( new_AGEMA_signal_21183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C ( clk ), .D ( new_AGEMA_signal_21184 ), .Q ( new_AGEMA_signal_21185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C ( clk ), .D ( new_AGEMA_signal_21186 ), .Q ( new_AGEMA_signal_21187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C ( clk ), .D ( new_AGEMA_signal_21188 ), .Q ( new_AGEMA_signal_21189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C ( clk ), .D ( new_AGEMA_signal_21190 ), .Q ( new_AGEMA_signal_21191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C ( clk ), .D ( new_AGEMA_signal_21194 ), .Q ( new_AGEMA_signal_21195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C ( clk ), .D ( new_AGEMA_signal_21198 ), .Q ( new_AGEMA_signal_21199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C ( clk ), .D ( new_AGEMA_signal_21202 ), .Q ( new_AGEMA_signal_21203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C ( clk ), .D ( new_AGEMA_signal_21206 ), .Q ( new_AGEMA_signal_21207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C ( clk ), .D ( new_AGEMA_signal_21210 ), .Q ( new_AGEMA_signal_21211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C ( clk ), .D ( new_AGEMA_signal_21212 ), .Q ( new_AGEMA_signal_21213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C ( clk ), .D ( new_AGEMA_signal_21214 ), .Q ( new_AGEMA_signal_21215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C ( clk ), .D ( new_AGEMA_signal_21216 ), .Q ( new_AGEMA_signal_21217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C ( clk ), .D ( new_AGEMA_signal_21218 ), .Q ( new_AGEMA_signal_21219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C ( clk ), .D ( new_AGEMA_signal_21220 ), .Q ( new_AGEMA_signal_21221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C ( clk ), .D ( new_AGEMA_signal_21226 ), .Q ( new_AGEMA_signal_21227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C ( clk ), .D ( new_AGEMA_signal_21232 ), .Q ( new_AGEMA_signal_21233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C ( clk ), .D ( new_AGEMA_signal_21238 ), .Q ( new_AGEMA_signal_21239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C ( clk ), .D ( new_AGEMA_signal_21244 ), .Q ( new_AGEMA_signal_21245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C ( clk ), .D ( new_AGEMA_signal_21250 ), .Q ( new_AGEMA_signal_21251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C ( clk ), .D ( new_AGEMA_signal_21256 ), .Q ( new_AGEMA_signal_21257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C ( clk ), .D ( new_AGEMA_signal_21262 ), .Q ( new_AGEMA_signal_21263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C ( clk ), .D ( new_AGEMA_signal_21268 ), .Q ( new_AGEMA_signal_21269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C ( clk ), .D ( new_AGEMA_signal_21274 ), .Q ( new_AGEMA_signal_21275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C ( clk ), .D ( new_AGEMA_signal_21280 ), .Q ( new_AGEMA_signal_21281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C ( clk ), .D ( new_AGEMA_signal_21284 ), .Q ( new_AGEMA_signal_21285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C ( clk ), .D ( new_AGEMA_signal_21288 ), .Q ( new_AGEMA_signal_21289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C ( clk ), .D ( new_AGEMA_signal_21292 ), .Q ( new_AGEMA_signal_21293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C ( clk ), .D ( new_AGEMA_signal_21296 ), .Q ( new_AGEMA_signal_21297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C ( clk ), .D ( new_AGEMA_signal_21300 ), .Q ( new_AGEMA_signal_21301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C ( clk ), .D ( new_AGEMA_signal_21302 ), .Q ( new_AGEMA_signal_21303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C ( clk ), .D ( new_AGEMA_signal_21304 ), .Q ( new_AGEMA_signal_21305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C ( clk ), .D ( new_AGEMA_signal_21306 ), .Q ( new_AGEMA_signal_21307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C ( clk ), .D ( new_AGEMA_signal_21308 ), .Q ( new_AGEMA_signal_21309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C ( clk ), .D ( new_AGEMA_signal_21310 ), .Q ( new_AGEMA_signal_21311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C ( clk ), .D ( new_AGEMA_signal_21318 ), .Q ( new_AGEMA_signal_21319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C ( clk ), .D ( new_AGEMA_signal_21326 ), .Q ( new_AGEMA_signal_21327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C ( clk ), .D ( new_AGEMA_signal_21334 ), .Q ( new_AGEMA_signal_21335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C ( clk ), .D ( new_AGEMA_signal_21342 ), .Q ( new_AGEMA_signal_21343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C ( clk ), .D ( new_AGEMA_signal_21350 ), .Q ( new_AGEMA_signal_21351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C ( clk ), .D ( new_AGEMA_signal_21352 ), .Q ( new_AGEMA_signal_21353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C ( clk ), .D ( new_AGEMA_signal_21354 ), .Q ( new_AGEMA_signal_21355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C ( clk ), .D ( new_AGEMA_signal_21356 ), .Q ( new_AGEMA_signal_21357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C ( clk ), .D ( new_AGEMA_signal_21358 ), .Q ( new_AGEMA_signal_21359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C ( clk ), .D ( new_AGEMA_signal_21360 ), .Q ( new_AGEMA_signal_21361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C ( clk ), .D ( new_AGEMA_signal_21364 ), .Q ( new_AGEMA_signal_21365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C ( clk ), .D ( new_AGEMA_signal_21368 ), .Q ( new_AGEMA_signal_21369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C ( clk ), .D ( new_AGEMA_signal_21372 ), .Q ( new_AGEMA_signal_21373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C ( clk ), .D ( new_AGEMA_signal_21376 ), .Q ( new_AGEMA_signal_21377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C ( clk ), .D ( new_AGEMA_signal_21380 ), .Q ( new_AGEMA_signal_21381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C ( clk ), .D ( new_AGEMA_signal_21384 ), .Q ( new_AGEMA_signal_21385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C ( clk ), .D ( new_AGEMA_signal_21388 ), .Q ( new_AGEMA_signal_21389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C ( clk ), .D ( new_AGEMA_signal_21392 ), .Q ( new_AGEMA_signal_21393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C ( clk ), .D ( new_AGEMA_signal_21396 ), .Q ( new_AGEMA_signal_21397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C ( clk ), .D ( new_AGEMA_signal_21400 ), .Q ( new_AGEMA_signal_21401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C ( clk ), .D ( new_AGEMA_signal_21404 ), .Q ( new_AGEMA_signal_21405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C ( clk ), .D ( new_AGEMA_signal_21408 ), .Q ( new_AGEMA_signal_21409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C ( clk ), .D ( new_AGEMA_signal_21412 ), .Q ( new_AGEMA_signal_21413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C ( clk ), .D ( new_AGEMA_signal_21416 ), .Q ( new_AGEMA_signal_21417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C ( clk ), .D ( new_AGEMA_signal_21420 ), .Q ( new_AGEMA_signal_21421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C ( clk ), .D ( new_AGEMA_signal_21424 ), .Q ( new_AGEMA_signal_21425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C ( clk ), .D ( new_AGEMA_signal_21428 ), .Q ( new_AGEMA_signal_21429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C ( clk ), .D ( new_AGEMA_signal_21432 ), .Q ( new_AGEMA_signal_21433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C ( clk ), .D ( new_AGEMA_signal_21436 ), .Q ( new_AGEMA_signal_21437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C ( clk ), .D ( new_AGEMA_signal_21440 ), .Q ( new_AGEMA_signal_21441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C ( clk ), .D ( new_AGEMA_signal_21444 ), .Q ( new_AGEMA_signal_21445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C ( clk ), .D ( new_AGEMA_signal_21448 ), .Q ( new_AGEMA_signal_21449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C ( clk ), .D ( new_AGEMA_signal_21452 ), .Q ( new_AGEMA_signal_21453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C ( clk ), .D ( new_AGEMA_signal_21456 ), .Q ( new_AGEMA_signal_21457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C ( clk ), .D ( new_AGEMA_signal_21460 ), .Q ( new_AGEMA_signal_21461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C ( clk ), .D ( new_AGEMA_signal_21468 ), .Q ( new_AGEMA_signal_21469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C ( clk ), .D ( new_AGEMA_signal_21476 ), .Q ( new_AGEMA_signal_21477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C ( clk ), .D ( new_AGEMA_signal_21484 ), .Q ( new_AGEMA_signal_21485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C ( clk ), .D ( new_AGEMA_signal_21492 ), .Q ( new_AGEMA_signal_21493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C ( clk ), .D ( new_AGEMA_signal_21500 ), .Q ( new_AGEMA_signal_21501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C ( clk ), .D ( new_AGEMA_signal_21502 ), .Q ( new_AGEMA_signal_21503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C ( clk ), .D ( new_AGEMA_signal_21504 ), .Q ( new_AGEMA_signal_21505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C ( clk ), .D ( new_AGEMA_signal_21506 ), .Q ( new_AGEMA_signal_21507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C ( clk ), .D ( new_AGEMA_signal_21508 ), .Q ( new_AGEMA_signal_21509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C ( clk ), .D ( new_AGEMA_signal_21510 ), .Q ( new_AGEMA_signal_21511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C ( clk ), .D ( new_AGEMA_signal_21514 ), .Q ( new_AGEMA_signal_21515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C ( clk ), .D ( new_AGEMA_signal_21518 ), .Q ( new_AGEMA_signal_21519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C ( clk ), .D ( new_AGEMA_signal_21522 ), .Q ( new_AGEMA_signal_21523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C ( clk ), .D ( new_AGEMA_signal_21526 ), .Q ( new_AGEMA_signal_21527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C ( clk ), .D ( new_AGEMA_signal_21530 ), .Q ( new_AGEMA_signal_21531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C ( clk ), .D ( new_AGEMA_signal_21532 ), .Q ( new_AGEMA_signal_21533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C ( clk ), .D ( new_AGEMA_signal_21534 ), .Q ( new_AGEMA_signal_21535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C ( clk ), .D ( new_AGEMA_signal_21536 ), .Q ( new_AGEMA_signal_21537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C ( clk ), .D ( new_AGEMA_signal_21538 ), .Q ( new_AGEMA_signal_21539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C ( clk ), .D ( new_AGEMA_signal_21540 ), .Q ( new_AGEMA_signal_21541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C ( clk ), .D ( new_AGEMA_signal_21546 ), .Q ( new_AGEMA_signal_21547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C ( clk ), .D ( new_AGEMA_signal_21552 ), .Q ( new_AGEMA_signal_21553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C ( clk ), .D ( new_AGEMA_signal_21558 ), .Q ( new_AGEMA_signal_21559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C ( clk ), .D ( new_AGEMA_signal_21564 ), .Q ( new_AGEMA_signal_21565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C ( clk ), .D ( new_AGEMA_signal_21570 ), .Q ( new_AGEMA_signal_21571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C ( clk ), .D ( new_AGEMA_signal_21586 ), .Q ( new_AGEMA_signal_21587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C ( clk ), .D ( new_AGEMA_signal_21594 ), .Q ( new_AGEMA_signal_21595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C ( clk ), .D ( new_AGEMA_signal_21602 ), .Q ( new_AGEMA_signal_21603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C ( clk ), .D ( new_AGEMA_signal_21610 ), .Q ( new_AGEMA_signal_21611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C ( clk ), .D ( new_AGEMA_signal_21618 ), .Q ( new_AGEMA_signal_21619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C ( clk ), .D ( new_AGEMA_signal_21632 ), .Q ( new_AGEMA_signal_21633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C ( clk ), .D ( new_AGEMA_signal_21636 ), .Q ( new_AGEMA_signal_21637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C ( clk ), .D ( new_AGEMA_signal_21640 ), .Q ( new_AGEMA_signal_21641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C ( clk ), .D ( new_AGEMA_signal_21644 ), .Q ( new_AGEMA_signal_21645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C ( clk ), .D ( new_AGEMA_signal_21648 ), .Q ( new_AGEMA_signal_21649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C ( clk ), .D ( new_AGEMA_signal_21656 ), .Q ( new_AGEMA_signal_21657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C ( clk ), .D ( new_AGEMA_signal_21664 ), .Q ( new_AGEMA_signal_21665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C ( clk ), .D ( new_AGEMA_signal_21672 ), .Q ( new_AGEMA_signal_21673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C ( clk ), .D ( new_AGEMA_signal_21680 ), .Q ( new_AGEMA_signal_21681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C ( clk ), .D ( new_AGEMA_signal_21688 ), .Q ( new_AGEMA_signal_21689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C ( clk ), .D ( new_AGEMA_signal_21704 ), .Q ( new_AGEMA_signal_21705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C ( clk ), .D ( new_AGEMA_signal_21710 ), .Q ( new_AGEMA_signal_21711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C ( clk ), .D ( new_AGEMA_signal_21716 ), .Q ( new_AGEMA_signal_21717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C ( clk ), .D ( new_AGEMA_signal_21722 ), .Q ( new_AGEMA_signal_21723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C ( clk ), .D ( new_AGEMA_signal_21728 ), .Q ( new_AGEMA_signal_21729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C ( clk ), .D ( new_AGEMA_signal_21732 ), .Q ( new_AGEMA_signal_21733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C ( clk ), .D ( new_AGEMA_signal_21736 ), .Q ( new_AGEMA_signal_21737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C ( clk ), .D ( new_AGEMA_signal_21740 ), .Q ( new_AGEMA_signal_21741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C ( clk ), .D ( new_AGEMA_signal_21744 ), .Q ( new_AGEMA_signal_21745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C ( clk ), .D ( new_AGEMA_signal_21748 ), .Q ( new_AGEMA_signal_21749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C ( clk ), .D ( new_AGEMA_signal_21756 ), .Q ( new_AGEMA_signal_21757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C ( clk ), .D ( new_AGEMA_signal_21764 ), .Q ( new_AGEMA_signal_21765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C ( clk ), .D ( new_AGEMA_signal_21772 ), .Q ( new_AGEMA_signal_21773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C ( clk ), .D ( new_AGEMA_signal_21780 ), .Q ( new_AGEMA_signal_21781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C ( clk ), .D ( new_AGEMA_signal_21788 ), .Q ( new_AGEMA_signal_21789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C ( clk ), .D ( new_AGEMA_signal_21792 ), .Q ( new_AGEMA_signal_21793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C ( clk ), .D ( new_AGEMA_signal_21796 ), .Q ( new_AGEMA_signal_21797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C ( clk ), .D ( new_AGEMA_signal_21800 ), .Q ( new_AGEMA_signal_21801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C ( clk ), .D ( new_AGEMA_signal_21804 ), .Q ( new_AGEMA_signal_21805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C ( clk ), .D ( new_AGEMA_signal_21808 ), .Q ( new_AGEMA_signal_21809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C ( clk ), .D ( new_AGEMA_signal_21814 ), .Q ( new_AGEMA_signal_21815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C ( clk ), .D ( new_AGEMA_signal_21820 ), .Q ( new_AGEMA_signal_21821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C ( clk ), .D ( new_AGEMA_signal_21826 ), .Q ( new_AGEMA_signal_21827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C ( clk ), .D ( new_AGEMA_signal_21832 ), .Q ( new_AGEMA_signal_21833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C ( clk ), .D ( new_AGEMA_signal_21838 ), .Q ( new_AGEMA_signal_21839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C ( clk ), .D ( new_AGEMA_signal_21844 ), .Q ( new_AGEMA_signal_21845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C ( clk ), .D ( new_AGEMA_signal_21850 ), .Q ( new_AGEMA_signal_21851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C ( clk ), .D ( new_AGEMA_signal_21856 ), .Q ( new_AGEMA_signal_21857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C ( clk ), .D ( new_AGEMA_signal_21862 ), .Q ( new_AGEMA_signal_21863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C ( clk ), .D ( new_AGEMA_signal_21868 ), .Q ( new_AGEMA_signal_21869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C ( clk ), .D ( new_AGEMA_signal_21874 ), .Q ( new_AGEMA_signal_21875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C ( clk ), .D ( new_AGEMA_signal_21880 ), .Q ( new_AGEMA_signal_21881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C ( clk ), .D ( new_AGEMA_signal_21886 ), .Q ( new_AGEMA_signal_21887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C ( clk ), .D ( new_AGEMA_signal_21892 ), .Q ( new_AGEMA_signal_21893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C ( clk ), .D ( new_AGEMA_signal_21898 ), .Q ( new_AGEMA_signal_21899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C ( clk ), .D ( new_AGEMA_signal_21904 ), .Q ( new_AGEMA_signal_21905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C ( clk ), .D ( new_AGEMA_signal_21910 ), .Q ( new_AGEMA_signal_21911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C ( clk ), .D ( new_AGEMA_signal_21916 ), .Q ( new_AGEMA_signal_21917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C ( clk ), .D ( new_AGEMA_signal_21922 ), .Q ( new_AGEMA_signal_21923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C ( clk ), .D ( new_AGEMA_signal_21928 ), .Q ( new_AGEMA_signal_21929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C ( clk ), .D ( new_AGEMA_signal_21934 ), .Q ( new_AGEMA_signal_21935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C ( clk ), .D ( new_AGEMA_signal_21940 ), .Q ( new_AGEMA_signal_21941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C ( clk ), .D ( new_AGEMA_signal_21946 ), .Q ( new_AGEMA_signal_21947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C ( clk ), .D ( new_AGEMA_signal_21952 ), .Q ( new_AGEMA_signal_21953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C ( clk ), .D ( new_AGEMA_signal_21958 ), .Q ( new_AGEMA_signal_21959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C ( clk ), .D ( new_AGEMA_signal_21962 ), .Q ( new_AGEMA_signal_21963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C ( clk ), .D ( new_AGEMA_signal_21966 ), .Q ( new_AGEMA_signal_21967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C ( clk ), .D ( new_AGEMA_signal_21970 ), .Q ( new_AGEMA_signal_21971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C ( clk ), .D ( new_AGEMA_signal_21974 ), .Q ( new_AGEMA_signal_21975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C ( clk ), .D ( new_AGEMA_signal_21978 ), .Q ( new_AGEMA_signal_21979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C ( clk ), .D ( new_AGEMA_signal_21986 ), .Q ( new_AGEMA_signal_21987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C ( clk ), .D ( new_AGEMA_signal_21994 ), .Q ( new_AGEMA_signal_21995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C ( clk ), .D ( new_AGEMA_signal_22002 ), .Q ( new_AGEMA_signal_22003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C ( clk ), .D ( new_AGEMA_signal_22010 ), .Q ( new_AGEMA_signal_22011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C ( clk ), .D ( new_AGEMA_signal_22018 ), .Q ( new_AGEMA_signal_22019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C ( clk ), .D ( new_AGEMA_signal_22022 ), .Q ( new_AGEMA_signal_22023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C ( clk ), .D ( new_AGEMA_signal_22026 ), .Q ( new_AGEMA_signal_22027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C ( clk ), .D ( new_AGEMA_signal_22030 ), .Q ( new_AGEMA_signal_22031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C ( clk ), .D ( new_AGEMA_signal_22034 ), .Q ( new_AGEMA_signal_22035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C ( clk ), .D ( new_AGEMA_signal_22038 ), .Q ( new_AGEMA_signal_22039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C ( clk ), .D ( new_AGEMA_signal_22044 ), .Q ( new_AGEMA_signal_22045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C ( clk ), .D ( new_AGEMA_signal_22050 ), .Q ( new_AGEMA_signal_22051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C ( clk ), .D ( new_AGEMA_signal_22056 ), .Q ( new_AGEMA_signal_22057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C ( clk ), .D ( new_AGEMA_signal_22062 ), .Q ( new_AGEMA_signal_22063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C ( clk ), .D ( new_AGEMA_signal_22068 ), .Q ( new_AGEMA_signal_22069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C ( clk ), .D ( new_AGEMA_signal_22076 ), .Q ( new_AGEMA_signal_22077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C ( clk ), .D ( new_AGEMA_signal_22084 ), .Q ( new_AGEMA_signal_22085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C ( clk ), .D ( new_AGEMA_signal_22092 ), .Q ( new_AGEMA_signal_22093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C ( clk ), .D ( new_AGEMA_signal_22100 ), .Q ( new_AGEMA_signal_22101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C ( clk ), .D ( new_AGEMA_signal_22108 ), .Q ( new_AGEMA_signal_22109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C ( clk ), .D ( new_AGEMA_signal_22124 ), .Q ( new_AGEMA_signal_22125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C ( clk ), .D ( new_AGEMA_signal_22130 ), .Q ( new_AGEMA_signal_22131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C ( clk ), .D ( new_AGEMA_signal_22136 ), .Q ( new_AGEMA_signal_22137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C ( clk ), .D ( new_AGEMA_signal_22142 ), .Q ( new_AGEMA_signal_22143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C ( clk ), .D ( new_AGEMA_signal_22148 ), .Q ( new_AGEMA_signal_22149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C ( clk ), .D ( new_AGEMA_signal_22174 ), .Q ( new_AGEMA_signal_22175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C ( clk ), .D ( new_AGEMA_signal_22180 ), .Q ( new_AGEMA_signal_22181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C ( clk ), .D ( new_AGEMA_signal_22186 ), .Q ( new_AGEMA_signal_22187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C ( clk ), .D ( new_AGEMA_signal_22192 ), .Q ( new_AGEMA_signal_22193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C ( clk ), .D ( new_AGEMA_signal_22198 ), .Q ( new_AGEMA_signal_22199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C ( clk ), .D ( new_AGEMA_signal_22204 ), .Q ( new_AGEMA_signal_22205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C ( clk ), .D ( new_AGEMA_signal_22210 ), .Q ( new_AGEMA_signal_22211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C ( clk ), .D ( new_AGEMA_signal_22216 ), .Q ( new_AGEMA_signal_22217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C ( clk ), .D ( new_AGEMA_signal_22222 ), .Q ( new_AGEMA_signal_22223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C ( clk ), .D ( new_AGEMA_signal_22228 ), .Q ( new_AGEMA_signal_22229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C ( clk ), .D ( new_AGEMA_signal_22236 ), .Q ( new_AGEMA_signal_22237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C ( clk ), .D ( new_AGEMA_signal_22244 ), .Q ( new_AGEMA_signal_22245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C ( clk ), .D ( new_AGEMA_signal_22252 ), .Q ( new_AGEMA_signal_22253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C ( clk ), .D ( new_AGEMA_signal_22260 ), .Q ( new_AGEMA_signal_22261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C ( clk ), .D ( new_AGEMA_signal_22268 ), .Q ( new_AGEMA_signal_22269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C ( clk ), .D ( new_AGEMA_signal_22276 ), .Q ( new_AGEMA_signal_22277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C ( clk ), .D ( new_AGEMA_signal_22284 ), .Q ( new_AGEMA_signal_22285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C ( clk ), .D ( new_AGEMA_signal_22292 ), .Q ( new_AGEMA_signal_22293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C ( clk ), .D ( new_AGEMA_signal_22300 ), .Q ( new_AGEMA_signal_22301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C ( clk ), .D ( new_AGEMA_signal_22308 ), .Q ( new_AGEMA_signal_22309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C ( clk ), .D ( new_AGEMA_signal_22314 ), .Q ( new_AGEMA_signal_22315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C ( clk ), .D ( new_AGEMA_signal_22320 ), .Q ( new_AGEMA_signal_22321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C ( clk ), .D ( new_AGEMA_signal_22326 ), .Q ( new_AGEMA_signal_22327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C ( clk ), .D ( new_AGEMA_signal_22332 ), .Q ( new_AGEMA_signal_22333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C ( clk ), .D ( new_AGEMA_signal_22338 ), .Q ( new_AGEMA_signal_22339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C ( clk ), .D ( new_AGEMA_signal_22344 ), .Q ( new_AGEMA_signal_22345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C ( clk ), .D ( new_AGEMA_signal_22350 ), .Q ( new_AGEMA_signal_22351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C ( clk ), .D ( new_AGEMA_signal_22356 ), .Q ( new_AGEMA_signal_22357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C ( clk ), .D ( new_AGEMA_signal_22362 ), .Q ( new_AGEMA_signal_22363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C ( clk ), .D ( new_AGEMA_signal_22368 ), .Q ( new_AGEMA_signal_22369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C ( clk ), .D ( new_AGEMA_signal_22382 ), .Q ( new_AGEMA_signal_22383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C ( clk ), .D ( new_AGEMA_signal_22386 ), .Q ( new_AGEMA_signal_22387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C ( clk ), .D ( new_AGEMA_signal_22390 ), .Q ( new_AGEMA_signal_22391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C ( clk ), .D ( new_AGEMA_signal_22394 ), .Q ( new_AGEMA_signal_22395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C ( clk ), .D ( new_AGEMA_signal_22398 ), .Q ( new_AGEMA_signal_22399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C ( clk ), .D ( new_AGEMA_signal_22402 ), .Q ( new_AGEMA_signal_22403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C ( clk ), .D ( new_AGEMA_signal_22406 ), .Q ( new_AGEMA_signal_22407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C ( clk ), .D ( new_AGEMA_signal_22410 ), .Q ( new_AGEMA_signal_22411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C ( clk ), .D ( new_AGEMA_signal_22414 ), .Q ( new_AGEMA_signal_22415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C ( clk ), .D ( new_AGEMA_signal_22418 ), .Q ( new_AGEMA_signal_22419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C ( clk ), .D ( new_AGEMA_signal_22422 ), .Q ( new_AGEMA_signal_22423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C ( clk ), .D ( new_AGEMA_signal_22426 ), .Q ( new_AGEMA_signal_22427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C ( clk ), .D ( new_AGEMA_signal_22430 ), .Q ( new_AGEMA_signal_22431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C ( clk ), .D ( new_AGEMA_signal_22434 ), .Q ( new_AGEMA_signal_22435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C ( clk ), .D ( new_AGEMA_signal_22438 ), .Q ( new_AGEMA_signal_22439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C ( clk ), .D ( new_AGEMA_signal_22452 ), .Q ( new_AGEMA_signal_22453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C ( clk ), .D ( new_AGEMA_signal_22458 ), .Q ( new_AGEMA_signal_22459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C ( clk ), .D ( new_AGEMA_signal_22464 ), .Q ( new_AGEMA_signal_22465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C ( clk ), .D ( new_AGEMA_signal_22470 ), .Q ( new_AGEMA_signal_22471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C ( clk ), .D ( new_AGEMA_signal_22476 ), .Q ( new_AGEMA_signal_22477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C ( clk ), .D ( new_AGEMA_signal_22514 ), .Q ( new_AGEMA_signal_22515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C ( clk ), .D ( new_AGEMA_signal_22522 ), .Q ( new_AGEMA_signal_22523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C ( clk ), .D ( new_AGEMA_signal_22530 ), .Q ( new_AGEMA_signal_22531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C ( clk ), .D ( new_AGEMA_signal_22538 ), .Q ( new_AGEMA_signal_22539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C ( clk ), .D ( new_AGEMA_signal_22546 ), .Q ( new_AGEMA_signal_22547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C ( clk ), .D ( new_AGEMA_signal_22554 ), .Q ( new_AGEMA_signal_22555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C ( clk ), .D ( new_AGEMA_signal_22562 ), .Q ( new_AGEMA_signal_22563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C ( clk ), .D ( new_AGEMA_signal_22570 ), .Q ( new_AGEMA_signal_22571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C ( clk ), .D ( new_AGEMA_signal_22578 ), .Q ( new_AGEMA_signal_22579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C ( clk ), .D ( new_AGEMA_signal_22586 ), .Q ( new_AGEMA_signal_22587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C ( clk ), .D ( new_AGEMA_signal_22594 ), .Q ( new_AGEMA_signal_22595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C ( clk ), .D ( new_AGEMA_signal_22602 ), .Q ( new_AGEMA_signal_22603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C ( clk ), .D ( new_AGEMA_signal_22610 ), .Q ( new_AGEMA_signal_22611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C ( clk ), .D ( new_AGEMA_signal_22618 ), .Q ( new_AGEMA_signal_22619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C ( clk ), .D ( new_AGEMA_signal_22626 ), .Q ( new_AGEMA_signal_22627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C ( clk ), .D ( new_AGEMA_signal_22634 ), .Q ( new_AGEMA_signal_22635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C ( clk ), .D ( new_AGEMA_signal_22642 ), .Q ( new_AGEMA_signal_22643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C ( clk ), .D ( new_AGEMA_signal_22650 ), .Q ( new_AGEMA_signal_22651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C ( clk ), .D ( new_AGEMA_signal_22658 ), .Q ( new_AGEMA_signal_22659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C ( clk ), .D ( new_AGEMA_signal_22666 ), .Q ( new_AGEMA_signal_22667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C ( clk ), .D ( new_AGEMA_signal_22672 ), .Q ( new_AGEMA_signal_22673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C ( clk ), .D ( new_AGEMA_signal_22678 ), .Q ( new_AGEMA_signal_22679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C ( clk ), .D ( new_AGEMA_signal_22684 ), .Q ( new_AGEMA_signal_22685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C ( clk ), .D ( new_AGEMA_signal_22690 ), .Q ( new_AGEMA_signal_22691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C ( clk ), .D ( new_AGEMA_signal_22696 ), .Q ( new_AGEMA_signal_22697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C ( clk ), .D ( new_AGEMA_signal_22706 ), .Q ( new_AGEMA_signal_22707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C ( clk ), .D ( new_AGEMA_signal_22716 ), .Q ( new_AGEMA_signal_22717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C ( clk ), .D ( new_AGEMA_signal_22726 ), .Q ( new_AGEMA_signal_22727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C ( clk ), .D ( new_AGEMA_signal_22736 ), .Q ( new_AGEMA_signal_22737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C ( clk ), .D ( new_AGEMA_signal_22746 ), .Q ( new_AGEMA_signal_22747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C ( clk ), .D ( new_AGEMA_signal_22754 ), .Q ( new_AGEMA_signal_22755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C ( clk ), .D ( new_AGEMA_signal_22762 ), .Q ( new_AGEMA_signal_22763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C ( clk ), .D ( new_AGEMA_signal_22770 ), .Q ( new_AGEMA_signal_22771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C ( clk ), .D ( new_AGEMA_signal_22778 ), .Q ( new_AGEMA_signal_22779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C ( clk ), .D ( new_AGEMA_signal_22786 ), .Q ( new_AGEMA_signal_22787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C ( clk ), .D ( new_AGEMA_signal_22794 ), .Q ( new_AGEMA_signal_22795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C ( clk ), .D ( new_AGEMA_signal_22802 ), .Q ( new_AGEMA_signal_22803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C ( clk ), .D ( new_AGEMA_signal_22810 ), .Q ( new_AGEMA_signal_22811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C ( clk ), .D ( new_AGEMA_signal_22818 ), .Q ( new_AGEMA_signal_22819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C ( clk ), .D ( new_AGEMA_signal_22826 ), .Q ( new_AGEMA_signal_22827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C ( clk ), .D ( new_AGEMA_signal_22834 ), .Q ( new_AGEMA_signal_22835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C ( clk ), .D ( new_AGEMA_signal_22842 ), .Q ( new_AGEMA_signal_22843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C ( clk ), .D ( new_AGEMA_signal_22850 ), .Q ( new_AGEMA_signal_22851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C ( clk ), .D ( new_AGEMA_signal_22858 ), .Q ( new_AGEMA_signal_22859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C ( clk ), .D ( new_AGEMA_signal_22866 ), .Q ( new_AGEMA_signal_22867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C ( clk ), .D ( new_AGEMA_signal_22902 ), .Q ( new_AGEMA_signal_22903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C ( clk ), .D ( new_AGEMA_signal_22908 ), .Q ( new_AGEMA_signal_22909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C ( clk ), .D ( new_AGEMA_signal_22914 ), .Q ( new_AGEMA_signal_22915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C ( clk ), .D ( new_AGEMA_signal_22920 ), .Q ( new_AGEMA_signal_22921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C ( clk ), .D ( new_AGEMA_signal_22926 ), .Q ( new_AGEMA_signal_22927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C ( clk ), .D ( new_AGEMA_signal_22956 ), .Q ( new_AGEMA_signal_22957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C ( clk ), .D ( new_AGEMA_signal_22966 ), .Q ( new_AGEMA_signal_22967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C ( clk ), .D ( new_AGEMA_signal_22976 ), .Q ( new_AGEMA_signal_22977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C ( clk ), .D ( new_AGEMA_signal_22986 ), .Q ( new_AGEMA_signal_22987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C ( clk ), .D ( new_AGEMA_signal_22996 ), .Q ( new_AGEMA_signal_22997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C ( clk ), .D ( new_AGEMA_signal_23004 ), .Q ( new_AGEMA_signal_23005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C ( clk ), .D ( new_AGEMA_signal_23012 ), .Q ( new_AGEMA_signal_23013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C ( clk ), .D ( new_AGEMA_signal_23020 ), .Q ( new_AGEMA_signal_23021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C ( clk ), .D ( new_AGEMA_signal_23028 ), .Q ( new_AGEMA_signal_23029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C ( clk ), .D ( new_AGEMA_signal_23036 ), .Q ( new_AGEMA_signal_23037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C ( clk ), .D ( new_AGEMA_signal_23074 ), .Q ( new_AGEMA_signal_23075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C ( clk ), .D ( new_AGEMA_signal_23082 ), .Q ( new_AGEMA_signal_23083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C ( clk ), .D ( new_AGEMA_signal_23090 ), .Q ( new_AGEMA_signal_23091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C ( clk ), .D ( new_AGEMA_signal_23098 ), .Q ( new_AGEMA_signal_23099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C ( clk ), .D ( new_AGEMA_signal_23106 ), .Q ( new_AGEMA_signal_23107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C ( clk ), .D ( new_AGEMA_signal_23114 ), .Q ( new_AGEMA_signal_23115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C ( clk ), .D ( new_AGEMA_signal_23122 ), .Q ( new_AGEMA_signal_23123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C ( clk ), .D ( new_AGEMA_signal_23130 ), .Q ( new_AGEMA_signal_23131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C ( clk ), .D ( new_AGEMA_signal_23138 ), .Q ( new_AGEMA_signal_23139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C ( clk ), .D ( new_AGEMA_signal_23146 ), .Q ( new_AGEMA_signal_23147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C ( clk ), .D ( new_AGEMA_signal_23152 ), .Q ( new_AGEMA_signal_23153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C ( clk ), .D ( new_AGEMA_signal_23158 ), .Q ( new_AGEMA_signal_23159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C ( clk ), .D ( new_AGEMA_signal_23164 ), .Q ( new_AGEMA_signal_23165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C ( clk ), .D ( new_AGEMA_signal_23170 ), .Q ( new_AGEMA_signal_23171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C ( clk ), .D ( new_AGEMA_signal_23176 ), .Q ( new_AGEMA_signal_23177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C ( clk ), .D ( new_AGEMA_signal_23204 ), .Q ( new_AGEMA_signal_23205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C ( clk ), .D ( new_AGEMA_signal_23212 ), .Q ( new_AGEMA_signal_23213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C ( clk ), .D ( new_AGEMA_signal_23220 ), .Q ( new_AGEMA_signal_23221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C ( clk ), .D ( new_AGEMA_signal_23228 ), .Q ( new_AGEMA_signal_23229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C ( clk ), .D ( new_AGEMA_signal_23236 ), .Q ( new_AGEMA_signal_23237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C ( clk ), .D ( new_AGEMA_signal_23362 ), .Q ( new_AGEMA_signal_23363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C ( clk ), .D ( new_AGEMA_signal_23370 ), .Q ( new_AGEMA_signal_23371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C ( clk ), .D ( new_AGEMA_signal_23378 ), .Q ( new_AGEMA_signal_23379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C ( clk ), .D ( new_AGEMA_signal_23386 ), .Q ( new_AGEMA_signal_23387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C ( clk ), .D ( new_AGEMA_signal_23394 ), .Q ( new_AGEMA_signal_23395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C ( clk ), .D ( new_AGEMA_signal_23452 ), .Q ( new_AGEMA_signal_23453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C ( clk ), .D ( new_AGEMA_signal_23460 ), .Q ( new_AGEMA_signal_23461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C ( clk ), .D ( new_AGEMA_signal_23468 ), .Q ( new_AGEMA_signal_23469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C ( clk ), .D ( new_AGEMA_signal_23476 ), .Q ( new_AGEMA_signal_23477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C ( clk ), .D ( new_AGEMA_signal_23484 ), .Q ( new_AGEMA_signal_23485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C ( clk ), .D ( new_AGEMA_signal_23492 ), .Q ( new_AGEMA_signal_23493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C ( clk ), .D ( new_AGEMA_signal_23500 ), .Q ( new_AGEMA_signal_23501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C ( clk ), .D ( new_AGEMA_signal_23508 ), .Q ( new_AGEMA_signal_23509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C ( clk ), .D ( new_AGEMA_signal_23516 ), .Q ( new_AGEMA_signal_23517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C ( clk ), .D ( new_AGEMA_signal_23524 ), .Q ( new_AGEMA_signal_23525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C ( clk ), .D ( new_AGEMA_signal_23534 ), .Q ( new_AGEMA_signal_23535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C ( clk ), .D ( new_AGEMA_signal_23544 ), .Q ( new_AGEMA_signal_23545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C ( clk ), .D ( new_AGEMA_signal_23554 ), .Q ( new_AGEMA_signal_23555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C ( clk ), .D ( new_AGEMA_signal_23564 ), .Q ( new_AGEMA_signal_23565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C ( clk ), .D ( new_AGEMA_signal_23574 ), .Q ( new_AGEMA_signal_23575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C ( clk ), .D ( new_AGEMA_signal_23582 ), .Q ( new_AGEMA_signal_23583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C ( clk ), .D ( new_AGEMA_signal_23590 ), .Q ( new_AGEMA_signal_23591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C ( clk ), .D ( new_AGEMA_signal_23598 ), .Q ( new_AGEMA_signal_23599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C ( clk ), .D ( new_AGEMA_signal_23606 ), .Q ( new_AGEMA_signal_23607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C ( clk ), .D ( new_AGEMA_signal_23614 ), .Q ( new_AGEMA_signal_23615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C ( clk ), .D ( new_AGEMA_signal_23702 ), .Q ( new_AGEMA_signal_23703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C ( clk ), .D ( new_AGEMA_signal_23710 ), .Q ( new_AGEMA_signal_23711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C ( clk ), .D ( new_AGEMA_signal_23718 ), .Q ( new_AGEMA_signal_23719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C ( clk ), .D ( new_AGEMA_signal_23726 ), .Q ( new_AGEMA_signal_23727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C ( clk ), .D ( new_AGEMA_signal_23734 ), .Q ( new_AGEMA_signal_23735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C ( clk ), .D ( new_AGEMA_signal_23782 ), .Q ( new_AGEMA_signal_23783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C ( clk ), .D ( new_AGEMA_signal_23790 ), .Q ( new_AGEMA_signal_23791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C ( clk ), .D ( new_AGEMA_signal_23798 ), .Q ( new_AGEMA_signal_23799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C ( clk ), .D ( new_AGEMA_signal_23806 ), .Q ( new_AGEMA_signal_23807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C ( clk ), .D ( new_AGEMA_signal_23814 ), .Q ( new_AGEMA_signal_23815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C ( clk ), .D ( new_AGEMA_signal_24002 ), .Q ( new_AGEMA_signal_24003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C ( clk ), .D ( new_AGEMA_signal_24012 ), .Q ( new_AGEMA_signal_24013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C ( clk ), .D ( new_AGEMA_signal_24022 ), .Q ( new_AGEMA_signal_24023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C ( clk ), .D ( new_AGEMA_signal_24032 ), .Q ( new_AGEMA_signal_24033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C ( clk ), .D ( new_AGEMA_signal_24042 ), .Q ( new_AGEMA_signal_24043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7678 ( .C ( clk ), .D ( new_AGEMA_signal_24452 ), .Q ( new_AGEMA_signal_24453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7690 ( .C ( clk ), .D ( new_AGEMA_signal_24464 ), .Q ( new_AGEMA_signal_24465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7702 ( .C ( clk ), .D ( new_AGEMA_signal_24476 ), .Q ( new_AGEMA_signal_24477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7714 ( .C ( clk ), .D ( new_AGEMA_signal_24488 ), .Q ( new_AGEMA_signal_24489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7726 ( .C ( clk ), .D ( new_AGEMA_signal_24500 ), .Q ( new_AGEMA_signal_24501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7740 ( .C ( clk ), .D ( new_AGEMA_signal_24514 ), .Q ( new_AGEMA_signal_24515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7754 ( .C ( clk ), .D ( new_AGEMA_signal_24528 ), .Q ( new_AGEMA_signal_24529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7768 ( .C ( clk ), .D ( new_AGEMA_signal_24542 ), .Q ( new_AGEMA_signal_24543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7782 ( .C ( clk ), .D ( new_AGEMA_signal_24556 ), .Q ( new_AGEMA_signal_24557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7796 ( .C ( clk ), .D ( new_AGEMA_signal_24570 ), .Q ( new_AGEMA_signal_24571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7850 ( .C ( clk ), .D ( new_AGEMA_signal_24624 ), .Q ( new_AGEMA_signal_24625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7864 ( .C ( clk ), .D ( new_AGEMA_signal_24638 ), .Q ( new_AGEMA_signal_24639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7878 ( .C ( clk ), .D ( new_AGEMA_signal_24652 ), .Q ( new_AGEMA_signal_24653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7892 ( .C ( clk ), .D ( new_AGEMA_signal_24666 ), .Q ( new_AGEMA_signal_24667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7906 ( .C ( clk ), .D ( new_AGEMA_signal_24680 ), .Q ( new_AGEMA_signal_24681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8030 ( .C ( clk ), .D ( new_AGEMA_signal_24804 ), .Q ( new_AGEMA_signal_24805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8046 ( .C ( clk ), .D ( new_AGEMA_signal_24820 ), .Q ( new_AGEMA_signal_24821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8062 ( .C ( clk ), .D ( new_AGEMA_signal_24836 ), .Q ( new_AGEMA_signal_24837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8078 ( .C ( clk ), .D ( new_AGEMA_signal_24852 ), .Q ( new_AGEMA_signal_24853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8094 ( .C ( clk ), .D ( new_AGEMA_signal_24868 ), .Q ( new_AGEMA_signal_24869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8140 ( .C ( clk ), .D ( new_AGEMA_signal_24914 ), .Q ( new_AGEMA_signal_24915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8156 ( .C ( clk ), .D ( new_AGEMA_signal_24930 ), .Q ( new_AGEMA_signal_24931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8172 ( .C ( clk ), .D ( new_AGEMA_signal_24946 ), .Q ( new_AGEMA_signal_24947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8188 ( .C ( clk ), .D ( new_AGEMA_signal_24962 ), .Q ( new_AGEMA_signal_24963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8204 ( .C ( clk ), .D ( new_AGEMA_signal_24978 ), .Q ( new_AGEMA_signal_24979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8388 ( .C ( clk ), .D ( new_AGEMA_signal_25162 ), .Q ( new_AGEMA_signal_25163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8404 ( .C ( clk ), .D ( new_AGEMA_signal_25178 ), .Q ( new_AGEMA_signal_25179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8420 ( .C ( clk ), .D ( new_AGEMA_signal_25194 ), .Q ( new_AGEMA_signal_25195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8436 ( .C ( clk ), .D ( new_AGEMA_signal_25210 ), .Q ( new_AGEMA_signal_25211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8452 ( .C ( clk ), .D ( new_AGEMA_signal_25226 ), .Q ( new_AGEMA_signal_25227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8520 ( .C ( clk ), .D ( new_AGEMA_signal_25294 ), .Q ( new_AGEMA_signal_25295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8538 ( .C ( clk ), .D ( new_AGEMA_signal_25312 ), .Q ( new_AGEMA_signal_25313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8556 ( .C ( clk ), .D ( new_AGEMA_signal_25330 ), .Q ( new_AGEMA_signal_25331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8574 ( .C ( clk ), .D ( new_AGEMA_signal_25348 ), .Q ( new_AGEMA_signal_25349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8592 ( .C ( clk ), .D ( new_AGEMA_signal_25366 ), .Q ( new_AGEMA_signal_25367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8770 ( .C ( clk ), .D ( new_AGEMA_signal_25544 ), .Q ( new_AGEMA_signal_25545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8790 ( .C ( clk ), .D ( new_AGEMA_signal_25564 ), .Q ( new_AGEMA_signal_25565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8810 ( .C ( clk ), .D ( new_AGEMA_signal_25584 ), .Q ( new_AGEMA_signal_25585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8830 ( .C ( clk ), .D ( new_AGEMA_signal_25604 ), .Q ( new_AGEMA_signal_25605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8850 ( .C ( clk ), .D ( new_AGEMA_signal_25624 ), .Q ( new_AGEMA_signal_25625 ) ) ;

    /* cells in depth 11 */
    buf_clk new_AGEMA_reg_buffer_4797 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_21572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C ( clk ), .D ( new_AGEMA_signal_3514 ), .Q ( new_AGEMA_signal_21574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C ( clk ), .D ( new_AGEMA_signal_3515 ), .Q ( new_AGEMA_signal_21576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C ( clk ), .D ( new_AGEMA_signal_3516 ), .Q ( new_AGEMA_signal_21578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C ( clk ), .D ( new_AGEMA_signal_3517 ), .Q ( new_AGEMA_signal_21580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C ( clk ), .D ( new_AGEMA_signal_21587 ), .Q ( new_AGEMA_signal_21588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C ( clk ), .D ( new_AGEMA_signal_21595 ), .Q ( new_AGEMA_signal_21596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C ( clk ), .D ( new_AGEMA_signal_21603 ), .Q ( new_AGEMA_signal_21604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C ( clk ), .D ( new_AGEMA_signal_21611 ), .Q ( new_AGEMA_signal_21612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C ( clk ), .D ( new_AGEMA_signal_21619 ), .Q ( new_AGEMA_signal_21620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_21622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C ( clk ), .D ( new_AGEMA_signal_3546 ), .Q ( new_AGEMA_signal_21624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C ( clk ), .D ( new_AGEMA_signal_3547 ), .Q ( new_AGEMA_signal_21626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C ( clk ), .D ( new_AGEMA_signal_3548 ), .Q ( new_AGEMA_signal_21628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C ( clk ), .D ( new_AGEMA_signal_3549 ), .Q ( new_AGEMA_signal_21630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C ( clk ), .D ( new_AGEMA_signal_21633 ), .Q ( new_AGEMA_signal_21634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C ( clk ), .D ( new_AGEMA_signal_21637 ), .Q ( new_AGEMA_signal_21638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C ( clk ), .D ( new_AGEMA_signal_21641 ), .Q ( new_AGEMA_signal_21642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C ( clk ), .D ( new_AGEMA_signal_21645 ), .Q ( new_AGEMA_signal_21646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C ( clk ), .D ( new_AGEMA_signal_21649 ), .Q ( new_AGEMA_signal_21650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C ( clk ), .D ( new_AGEMA_signal_21657 ), .Q ( new_AGEMA_signal_21658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C ( clk ), .D ( new_AGEMA_signal_21665 ), .Q ( new_AGEMA_signal_21666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C ( clk ), .D ( new_AGEMA_signal_21673 ), .Q ( new_AGEMA_signal_21674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C ( clk ), .D ( new_AGEMA_signal_21681 ), .Q ( new_AGEMA_signal_21682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C ( clk ), .D ( new_AGEMA_signal_21689 ), .Q ( new_AGEMA_signal_21690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C ( clk ), .D ( new_AGEMA_signal_20509 ), .Q ( new_AGEMA_signal_21692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C ( clk ), .D ( new_AGEMA_signal_20517 ), .Q ( new_AGEMA_signal_21694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C ( clk ), .D ( new_AGEMA_signal_20525 ), .Q ( new_AGEMA_signal_21696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C ( clk ), .D ( new_AGEMA_signal_20533 ), .Q ( new_AGEMA_signal_21698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C ( clk ), .D ( new_AGEMA_signal_20541 ), .Q ( new_AGEMA_signal_21700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C ( clk ), .D ( new_AGEMA_signal_21705 ), .Q ( new_AGEMA_signal_21706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C ( clk ), .D ( new_AGEMA_signal_21711 ), .Q ( new_AGEMA_signal_21712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C ( clk ), .D ( new_AGEMA_signal_21717 ), .Q ( new_AGEMA_signal_21718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C ( clk ), .D ( new_AGEMA_signal_21723 ), .Q ( new_AGEMA_signal_21724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C ( clk ), .D ( new_AGEMA_signal_21729 ), .Q ( new_AGEMA_signal_21730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C ( clk ), .D ( new_AGEMA_signal_21733 ), .Q ( new_AGEMA_signal_21734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C ( clk ), .D ( new_AGEMA_signal_21737 ), .Q ( new_AGEMA_signal_21738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C ( clk ), .D ( new_AGEMA_signal_21741 ), .Q ( new_AGEMA_signal_21742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C ( clk ), .D ( new_AGEMA_signal_21745 ), .Q ( new_AGEMA_signal_21746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C ( clk ), .D ( new_AGEMA_signal_21749 ), .Q ( new_AGEMA_signal_21750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C ( clk ), .D ( new_AGEMA_signal_21757 ), .Q ( new_AGEMA_signal_21758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C ( clk ), .D ( new_AGEMA_signal_21765 ), .Q ( new_AGEMA_signal_21766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C ( clk ), .D ( new_AGEMA_signal_21773 ), .Q ( new_AGEMA_signal_21774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C ( clk ), .D ( new_AGEMA_signal_21781 ), .Q ( new_AGEMA_signal_21782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C ( clk ), .D ( new_AGEMA_signal_21789 ), .Q ( new_AGEMA_signal_21790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C ( clk ), .D ( new_AGEMA_signal_21793 ), .Q ( new_AGEMA_signal_21794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C ( clk ), .D ( new_AGEMA_signal_21797 ), .Q ( new_AGEMA_signal_21798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C ( clk ), .D ( new_AGEMA_signal_21801 ), .Q ( new_AGEMA_signal_21802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C ( clk ), .D ( new_AGEMA_signal_21805 ), .Q ( new_AGEMA_signal_21806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C ( clk ), .D ( new_AGEMA_signal_21809 ), .Q ( new_AGEMA_signal_21810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C ( clk ), .D ( new_AGEMA_signal_21815 ), .Q ( new_AGEMA_signal_21816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C ( clk ), .D ( new_AGEMA_signal_21821 ), .Q ( new_AGEMA_signal_21822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C ( clk ), .D ( new_AGEMA_signal_21827 ), .Q ( new_AGEMA_signal_21828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C ( clk ), .D ( new_AGEMA_signal_21833 ), .Q ( new_AGEMA_signal_21834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C ( clk ), .D ( new_AGEMA_signal_21839 ), .Q ( new_AGEMA_signal_21840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C ( clk ), .D ( new_AGEMA_signal_21845 ), .Q ( new_AGEMA_signal_21846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C ( clk ), .D ( new_AGEMA_signal_21851 ), .Q ( new_AGEMA_signal_21852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C ( clk ), .D ( new_AGEMA_signal_21857 ), .Q ( new_AGEMA_signal_21858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C ( clk ), .D ( new_AGEMA_signal_21863 ), .Q ( new_AGEMA_signal_21864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C ( clk ), .D ( new_AGEMA_signal_21869 ), .Q ( new_AGEMA_signal_21870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C ( clk ), .D ( new_AGEMA_signal_21875 ), .Q ( new_AGEMA_signal_21876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C ( clk ), .D ( new_AGEMA_signal_21881 ), .Q ( new_AGEMA_signal_21882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C ( clk ), .D ( new_AGEMA_signal_21887 ), .Q ( new_AGEMA_signal_21888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C ( clk ), .D ( new_AGEMA_signal_21893 ), .Q ( new_AGEMA_signal_21894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C ( clk ), .D ( new_AGEMA_signal_21899 ), .Q ( new_AGEMA_signal_21900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C ( clk ), .D ( new_AGEMA_signal_21905 ), .Q ( new_AGEMA_signal_21906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C ( clk ), .D ( new_AGEMA_signal_21911 ), .Q ( new_AGEMA_signal_21912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C ( clk ), .D ( new_AGEMA_signal_21917 ), .Q ( new_AGEMA_signal_21918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C ( clk ), .D ( new_AGEMA_signal_21923 ), .Q ( new_AGEMA_signal_21924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C ( clk ), .D ( new_AGEMA_signal_21929 ), .Q ( new_AGEMA_signal_21930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C ( clk ), .D ( new_AGEMA_signal_21935 ), .Q ( new_AGEMA_signal_21936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C ( clk ), .D ( new_AGEMA_signal_21941 ), .Q ( new_AGEMA_signal_21942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C ( clk ), .D ( new_AGEMA_signal_21947 ), .Q ( new_AGEMA_signal_21948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C ( clk ), .D ( new_AGEMA_signal_21953 ), .Q ( new_AGEMA_signal_21954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C ( clk ), .D ( new_AGEMA_signal_21959 ), .Q ( new_AGEMA_signal_21960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C ( clk ), .D ( new_AGEMA_signal_21963 ), .Q ( new_AGEMA_signal_21964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C ( clk ), .D ( new_AGEMA_signal_21967 ), .Q ( new_AGEMA_signal_21968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C ( clk ), .D ( new_AGEMA_signal_21971 ), .Q ( new_AGEMA_signal_21972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C ( clk ), .D ( new_AGEMA_signal_21975 ), .Q ( new_AGEMA_signal_21976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C ( clk ), .D ( new_AGEMA_signal_21979 ), .Q ( new_AGEMA_signal_21980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C ( clk ), .D ( new_AGEMA_signal_21987 ), .Q ( new_AGEMA_signal_21988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C ( clk ), .D ( new_AGEMA_signal_21995 ), .Q ( new_AGEMA_signal_21996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C ( clk ), .D ( new_AGEMA_signal_22003 ), .Q ( new_AGEMA_signal_22004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C ( clk ), .D ( new_AGEMA_signal_22011 ), .Q ( new_AGEMA_signal_22012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C ( clk ), .D ( new_AGEMA_signal_22019 ), .Q ( new_AGEMA_signal_22020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C ( clk ), .D ( new_AGEMA_signal_22023 ), .Q ( new_AGEMA_signal_22024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C ( clk ), .D ( new_AGEMA_signal_22027 ), .Q ( new_AGEMA_signal_22028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C ( clk ), .D ( new_AGEMA_signal_22031 ), .Q ( new_AGEMA_signal_22032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C ( clk ), .D ( new_AGEMA_signal_22035 ), .Q ( new_AGEMA_signal_22036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C ( clk ), .D ( new_AGEMA_signal_22039 ), .Q ( new_AGEMA_signal_22040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C ( clk ), .D ( new_AGEMA_signal_22045 ), .Q ( new_AGEMA_signal_22046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C ( clk ), .D ( new_AGEMA_signal_22051 ), .Q ( new_AGEMA_signal_22052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C ( clk ), .D ( new_AGEMA_signal_22057 ), .Q ( new_AGEMA_signal_22058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C ( clk ), .D ( new_AGEMA_signal_22063 ), .Q ( new_AGEMA_signal_22064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C ( clk ), .D ( new_AGEMA_signal_22069 ), .Q ( new_AGEMA_signal_22070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C ( clk ), .D ( new_AGEMA_signal_22077 ), .Q ( new_AGEMA_signal_22078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C ( clk ), .D ( new_AGEMA_signal_22085 ), .Q ( new_AGEMA_signal_22086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C ( clk ), .D ( new_AGEMA_signal_22093 ), .Q ( new_AGEMA_signal_22094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C ( clk ), .D ( new_AGEMA_signal_22101 ), .Q ( new_AGEMA_signal_22102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C ( clk ), .D ( new_AGEMA_signal_22109 ), .Q ( new_AGEMA_signal_22110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C ( clk ), .D ( new_AGEMA_signal_21213 ), .Q ( new_AGEMA_signal_22112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C ( clk ), .D ( new_AGEMA_signal_21215 ), .Q ( new_AGEMA_signal_22114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C ( clk ), .D ( new_AGEMA_signal_21217 ), .Q ( new_AGEMA_signal_22116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C ( clk ), .D ( new_AGEMA_signal_21219 ), .Q ( new_AGEMA_signal_22118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C ( clk ), .D ( new_AGEMA_signal_21221 ), .Q ( new_AGEMA_signal_22120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C ( clk ), .D ( new_AGEMA_signal_22125 ), .Q ( new_AGEMA_signal_22126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C ( clk ), .D ( new_AGEMA_signal_22131 ), .Q ( new_AGEMA_signal_22132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C ( clk ), .D ( new_AGEMA_signal_22137 ), .Q ( new_AGEMA_signal_22138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C ( clk ), .D ( new_AGEMA_signal_22143 ), .Q ( new_AGEMA_signal_22144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C ( clk ), .D ( new_AGEMA_signal_22149 ), .Q ( new_AGEMA_signal_22150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_22152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C ( clk ), .D ( new_AGEMA_signal_3702 ), .Q ( new_AGEMA_signal_22154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C ( clk ), .D ( new_AGEMA_signal_3703 ), .Q ( new_AGEMA_signal_22156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C ( clk ), .D ( new_AGEMA_signal_3704 ), .Q ( new_AGEMA_signal_22158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C ( clk ), .D ( new_AGEMA_signal_3705 ), .Q ( new_AGEMA_signal_22160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_22162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C ( clk ), .D ( new_AGEMA_signal_3706 ), .Q ( new_AGEMA_signal_22164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C ( clk ), .D ( new_AGEMA_signal_3707 ), .Q ( new_AGEMA_signal_22166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C ( clk ), .D ( new_AGEMA_signal_3708 ), .Q ( new_AGEMA_signal_22168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C ( clk ), .D ( new_AGEMA_signal_3709 ), .Q ( new_AGEMA_signal_22170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C ( clk ), .D ( new_AGEMA_signal_22175 ), .Q ( new_AGEMA_signal_22176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C ( clk ), .D ( new_AGEMA_signal_22181 ), .Q ( new_AGEMA_signal_22182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C ( clk ), .D ( new_AGEMA_signal_22187 ), .Q ( new_AGEMA_signal_22188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C ( clk ), .D ( new_AGEMA_signal_22193 ), .Q ( new_AGEMA_signal_22194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C ( clk ), .D ( new_AGEMA_signal_22199 ), .Q ( new_AGEMA_signal_22200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C ( clk ), .D ( new_AGEMA_signal_22205 ), .Q ( new_AGEMA_signal_22206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C ( clk ), .D ( new_AGEMA_signal_22211 ), .Q ( new_AGEMA_signal_22212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C ( clk ), .D ( new_AGEMA_signal_22217 ), .Q ( new_AGEMA_signal_22218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C ( clk ), .D ( new_AGEMA_signal_22223 ), .Q ( new_AGEMA_signal_22224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C ( clk ), .D ( new_AGEMA_signal_22229 ), .Q ( new_AGEMA_signal_22230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C ( clk ), .D ( new_AGEMA_signal_22237 ), .Q ( new_AGEMA_signal_22238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C ( clk ), .D ( new_AGEMA_signal_22245 ), .Q ( new_AGEMA_signal_22246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C ( clk ), .D ( new_AGEMA_signal_22253 ), .Q ( new_AGEMA_signal_22254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C ( clk ), .D ( new_AGEMA_signal_22261 ), .Q ( new_AGEMA_signal_22262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C ( clk ), .D ( new_AGEMA_signal_22269 ), .Q ( new_AGEMA_signal_22270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C ( clk ), .D ( new_AGEMA_signal_22277 ), .Q ( new_AGEMA_signal_22278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C ( clk ), .D ( new_AGEMA_signal_22285 ), .Q ( new_AGEMA_signal_22286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C ( clk ), .D ( new_AGEMA_signal_22293 ), .Q ( new_AGEMA_signal_22294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C ( clk ), .D ( new_AGEMA_signal_22301 ), .Q ( new_AGEMA_signal_22302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C ( clk ), .D ( new_AGEMA_signal_22309 ), .Q ( new_AGEMA_signal_22310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C ( clk ), .D ( new_AGEMA_signal_22315 ), .Q ( new_AGEMA_signal_22316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C ( clk ), .D ( new_AGEMA_signal_22321 ), .Q ( new_AGEMA_signal_22322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C ( clk ), .D ( new_AGEMA_signal_22327 ), .Q ( new_AGEMA_signal_22328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C ( clk ), .D ( new_AGEMA_signal_22333 ), .Q ( new_AGEMA_signal_22334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C ( clk ), .D ( new_AGEMA_signal_22339 ), .Q ( new_AGEMA_signal_22340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C ( clk ), .D ( new_AGEMA_signal_22345 ), .Q ( new_AGEMA_signal_22346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C ( clk ), .D ( new_AGEMA_signal_22351 ), .Q ( new_AGEMA_signal_22352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C ( clk ), .D ( new_AGEMA_signal_22357 ), .Q ( new_AGEMA_signal_22358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C ( clk ), .D ( new_AGEMA_signal_22363 ), .Q ( new_AGEMA_signal_22364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C ( clk ), .D ( new_AGEMA_signal_22369 ), .Q ( new_AGEMA_signal_22370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C ( clk ), .D ( new_AGEMA_signal_21165 ), .Q ( new_AGEMA_signal_22372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C ( clk ), .D ( new_AGEMA_signal_21169 ), .Q ( new_AGEMA_signal_22374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C ( clk ), .D ( new_AGEMA_signal_21173 ), .Q ( new_AGEMA_signal_22376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C ( clk ), .D ( new_AGEMA_signal_21177 ), .Q ( new_AGEMA_signal_22378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C ( clk ), .D ( new_AGEMA_signal_21181 ), .Q ( new_AGEMA_signal_22380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C ( clk ), .D ( new_AGEMA_signal_22383 ), .Q ( new_AGEMA_signal_22384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C ( clk ), .D ( new_AGEMA_signal_22387 ), .Q ( new_AGEMA_signal_22388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C ( clk ), .D ( new_AGEMA_signal_22391 ), .Q ( new_AGEMA_signal_22392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C ( clk ), .D ( new_AGEMA_signal_22395 ), .Q ( new_AGEMA_signal_22396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C ( clk ), .D ( new_AGEMA_signal_22399 ), .Q ( new_AGEMA_signal_22400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C ( clk ), .D ( new_AGEMA_signal_22403 ), .Q ( new_AGEMA_signal_22404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C ( clk ), .D ( new_AGEMA_signal_22407 ), .Q ( new_AGEMA_signal_22408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C ( clk ), .D ( new_AGEMA_signal_22411 ), .Q ( new_AGEMA_signal_22412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C ( clk ), .D ( new_AGEMA_signal_22415 ), .Q ( new_AGEMA_signal_22416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C ( clk ), .D ( new_AGEMA_signal_22419 ), .Q ( new_AGEMA_signal_22420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C ( clk ), .D ( new_AGEMA_signal_22423 ), .Q ( new_AGEMA_signal_22424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C ( clk ), .D ( new_AGEMA_signal_22427 ), .Q ( new_AGEMA_signal_22428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C ( clk ), .D ( new_AGEMA_signal_22431 ), .Q ( new_AGEMA_signal_22432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C ( clk ), .D ( new_AGEMA_signal_22435 ), .Q ( new_AGEMA_signal_22436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C ( clk ), .D ( new_AGEMA_signal_22439 ), .Q ( new_AGEMA_signal_22440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C ( clk ), .D ( new_AGEMA_signal_20889 ), .Q ( new_AGEMA_signal_22442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C ( clk ), .D ( new_AGEMA_signal_20897 ), .Q ( new_AGEMA_signal_22444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C ( clk ), .D ( new_AGEMA_signal_20905 ), .Q ( new_AGEMA_signal_22446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C ( clk ), .D ( new_AGEMA_signal_20913 ), .Q ( new_AGEMA_signal_22448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C ( clk ), .D ( new_AGEMA_signal_20921 ), .Q ( new_AGEMA_signal_22450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C ( clk ), .D ( new_AGEMA_signal_22453 ), .Q ( new_AGEMA_signal_22454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C ( clk ), .D ( new_AGEMA_signal_22459 ), .Q ( new_AGEMA_signal_22460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C ( clk ), .D ( new_AGEMA_signal_22465 ), .Q ( new_AGEMA_signal_22466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C ( clk ), .D ( new_AGEMA_signal_22471 ), .Q ( new_AGEMA_signal_22472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C ( clk ), .D ( new_AGEMA_signal_22477 ), .Q ( new_AGEMA_signal_22478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_22492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C ( clk ), .D ( new_AGEMA_signal_3850 ), .Q ( new_AGEMA_signal_22496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C ( clk ), .D ( new_AGEMA_signal_3851 ), .Q ( new_AGEMA_signal_22500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C ( clk ), .D ( new_AGEMA_signal_3852 ), .Q ( new_AGEMA_signal_22504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C ( clk ), .D ( new_AGEMA_signal_3853 ), .Q ( new_AGEMA_signal_22508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C ( clk ), .D ( new_AGEMA_signal_22515 ), .Q ( new_AGEMA_signal_22516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C ( clk ), .D ( new_AGEMA_signal_22523 ), .Q ( new_AGEMA_signal_22524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C ( clk ), .D ( new_AGEMA_signal_22531 ), .Q ( new_AGEMA_signal_22532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C ( clk ), .D ( new_AGEMA_signal_22539 ), .Q ( new_AGEMA_signal_22540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C ( clk ), .D ( new_AGEMA_signal_22547 ), .Q ( new_AGEMA_signal_22548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C ( clk ), .D ( new_AGEMA_signal_22555 ), .Q ( new_AGEMA_signal_22556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C ( clk ), .D ( new_AGEMA_signal_22563 ), .Q ( new_AGEMA_signal_22564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C ( clk ), .D ( new_AGEMA_signal_22571 ), .Q ( new_AGEMA_signal_22572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C ( clk ), .D ( new_AGEMA_signal_22579 ), .Q ( new_AGEMA_signal_22580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C ( clk ), .D ( new_AGEMA_signal_22587 ), .Q ( new_AGEMA_signal_22588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C ( clk ), .D ( new_AGEMA_signal_22595 ), .Q ( new_AGEMA_signal_22596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C ( clk ), .D ( new_AGEMA_signal_22603 ), .Q ( new_AGEMA_signal_22604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C ( clk ), .D ( new_AGEMA_signal_22611 ), .Q ( new_AGEMA_signal_22612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C ( clk ), .D ( new_AGEMA_signal_22619 ), .Q ( new_AGEMA_signal_22620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C ( clk ), .D ( new_AGEMA_signal_22627 ), .Q ( new_AGEMA_signal_22628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C ( clk ), .D ( new_AGEMA_signal_22635 ), .Q ( new_AGEMA_signal_22636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C ( clk ), .D ( new_AGEMA_signal_22643 ), .Q ( new_AGEMA_signal_22644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C ( clk ), .D ( new_AGEMA_signal_22651 ), .Q ( new_AGEMA_signal_22652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C ( clk ), .D ( new_AGEMA_signal_22659 ), .Q ( new_AGEMA_signal_22660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C ( clk ), .D ( new_AGEMA_signal_22667 ), .Q ( new_AGEMA_signal_22668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C ( clk ), .D ( new_AGEMA_signal_22673 ), .Q ( new_AGEMA_signal_22674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C ( clk ), .D ( new_AGEMA_signal_22679 ), .Q ( new_AGEMA_signal_22680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C ( clk ), .D ( new_AGEMA_signal_22685 ), .Q ( new_AGEMA_signal_22686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C ( clk ), .D ( new_AGEMA_signal_22691 ), .Q ( new_AGEMA_signal_22692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C ( clk ), .D ( new_AGEMA_signal_22697 ), .Q ( new_AGEMA_signal_22698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C ( clk ), .D ( new_AGEMA_signal_22707 ), .Q ( new_AGEMA_signal_22708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C ( clk ), .D ( new_AGEMA_signal_22717 ), .Q ( new_AGEMA_signal_22718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C ( clk ), .D ( new_AGEMA_signal_22727 ), .Q ( new_AGEMA_signal_22728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C ( clk ), .D ( new_AGEMA_signal_22737 ), .Q ( new_AGEMA_signal_22738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C ( clk ), .D ( new_AGEMA_signal_22747 ), .Q ( new_AGEMA_signal_22748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C ( clk ), .D ( new_AGEMA_signal_22755 ), .Q ( new_AGEMA_signal_22756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C ( clk ), .D ( new_AGEMA_signal_22763 ), .Q ( new_AGEMA_signal_22764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C ( clk ), .D ( new_AGEMA_signal_22771 ), .Q ( new_AGEMA_signal_22772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C ( clk ), .D ( new_AGEMA_signal_22779 ), .Q ( new_AGEMA_signal_22780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C ( clk ), .D ( new_AGEMA_signal_22787 ), .Q ( new_AGEMA_signal_22788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C ( clk ), .D ( new_AGEMA_signal_22795 ), .Q ( new_AGEMA_signal_22796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C ( clk ), .D ( new_AGEMA_signal_22803 ), .Q ( new_AGEMA_signal_22804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C ( clk ), .D ( new_AGEMA_signal_22811 ), .Q ( new_AGEMA_signal_22812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C ( clk ), .D ( new_AGEMA_signal_22819 ), .Q ( new_AGEMA_signal_22820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C ( clk ), .D ( new_AGEMA_signal_22827 ), .Q ( new_AGEMA_signal_22828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C ( clk ), .D ( new_AGEMA_signal_22835 ), .Q ( new_AGEMA_signal_22836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C ( clk ), .D ( new_AGEMA_signal_22843 ), .Q ( new_AGEMA_signal_22844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C ( clk ), .D ( new_AGEMA_signal_22851 ), .Q ( new_AGEMA_signal_22852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C ( clk ), .D ( new_AGEMA_signal_22859 ), .Q ( new_AGEMA_signal_22860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C ( clk ), .D ( new_AGEMA_signal_22867 ), .Q ( new_AGEMA_signal_22868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C ( clk ), .D ( new_AGEMA_signal_21195 ), .Q ( new_AGEMA_signal_22882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C ( clk ), .D ( new_AGEMA_signal_21199 ), .Q ( new_AGEMA_signal_22886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C ( clk ), .D ( new_AGEMA_signal_21203 ), .Q ( new_AGEMA_signal_22890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C ( clk ), .D ( new_AGEMA_signal_21207 ), .Q ( new_AGEMA_signal_22894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C ( clk ), .D ( new_AGEMA_signal_21211 ), .Q ( new_AGEMA_signal_22898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C ( clk ), .D ( new_AGEMA_signal_22903 ), .Q ( new_AGEMA_signal_22904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C ( clk ), .D ( new_AGEMA_signal_22909 ), .Q ( new_AGEMA_signal_22910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C ( clk ), .D ( new_AGEMA_signal_22915 ), .Q ( new_AGEMA_signal_22916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C ( clk ), .D ( new_AGEMA_signal_22921 ), .Q ( new_AGEMA_signal_22922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C ( clk ), .D ( new_AGEMA_signal_22927 ), .Q ( new_AGEMA_signal_22928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C ( clk ), .D ( new_AGEMA_signal_20637 ), .Q ( new_AGEMA_signal_22932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C ( clk ), .D ( new_AGEMA_signal_20643 ), .Q ( new_AGEMA_signal_22936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C ( clk ), .D ( new_AGEMA_signal_20649 ), .Q ( new_AGEMA_signal_22940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C ( clk ), .D ( new_AGEMA_signal_20655 ), .Q ( new_AGEMA_signal_22944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C ( clk ), .D ( new_AGEMA_signal_20661 ), .Q ( new_AGEMA_signal_22948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C ( clk ), .D ( new_AGEMA_signal_22957 ), .Q ( new_AGEMA_signal_22958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C ( clk ), .D ( new_AGEMA_signal_22967 ), .Q ( new_AGEMA_signal_22968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C ( clk ), .D ( new_AGEMA_signal_22977 ), .Q ( new_AGEMA_signal_22978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C ( clk ), .D ( new_AGEMA_signal_22987 ), .Q ( new_AGEMA_signal_22988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C ( clk ), .D ( new_AGEMA_signal_22997 ), .Q ( new_AGEMA_signal_22998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C ( clk ), .D ( new_AGEMA_signal_23005 ), .Q ( new_AGEMA_signal_23006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C ( clk ), .D ( new_AGEMA_signal_23013 ), .Q ( new_AGEMA_signal_23014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C ( clk ), .D ( new_AGEMA_signal_23021 ), .Q ( new_AGEMA_signal_23022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C ( clk ), .D ( new_AGEMA_signal_23029 ), .Q ( new_AGEMA_signal_23030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C ( clk ), .D ( new_AGEMA_signal_23037 ), .Q ( new_AGEMA_signal_23038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_23042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C ( clk ), .D ( new_AGEMA_signal_3386 ), .Q ( new_AGEMA_signal_23046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C ( clk ), .D ( new_AGEMA_signal_3387 ), .Q ( new_AGEMA_signal_23050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C ( clk ), .D ( new_AGEMA_signal_3388 ), .Q ( new_AGEMA_signal_23054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C ( clk ), .D ( new_AGEMA_signal_3389 ), .Q ( new_AGEMA_signal_23058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6301 ( .C ( clk ), .D ( new_AGEMA_signal_23075 ), .Q ( new_AGEMA_signal_23076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C ( clk ), .D ( new_AGEMA_signal_23083 ), .Q ( new_AGEMA_signal_23084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C ( clk ), .D ( new_AGEMA_signal_23091 ), .Q ( new_AGEMA_signal_23092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C ( clk ), .D ( new_AGEMA_signal_23099 ), .Q ( new_AGEMA_signal_23100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C ( clk ), .D ( new_AGEMA_signal_23107 ), .Q ( new_AGEMA_signal_23108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C ( clk ), .D ( new_AGEMA_signal_23115 ), .Q ( new_AGEMA_signal_23116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C ( clk ), .D ( new_AGEMA_signal_23123 ), .Q ( new_AGEMA_signal_23124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C ( clk ), .D ( new_AGEMA_signal_23131 ), .Q ( new_AGEMA_signal_23132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C ( clk ), .D ( new_AGEMA_signal_23139 ), .Q ( new_AGEMA_signal_23140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C ( clk ), .D ( new_AGEMA_signal_23147 ), .Q ( new_AGEMA_signal_23148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C ( clk ), .D ( new_AGEMA_signal_23153 ), .Q ( new_AGEMA_signal_23154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C ( clk ), .D ( new_AGEMA_signal_23159 ), .Q ( new_AGEMA_signal_23160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C ( clk ), .D ( new_AGEMA_signal_23165 ), .Q ( new_AGEMA_signal_23166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C ( clk ), .D ( new_AGEMA_signal_23171 ), .Q ( new_AGEMA_signal_23172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C ( clk ), .D ( new_AGEMA_signal_23177 ), .Q ( new_AGEMA_signal_23178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_23182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C ( clk ), .D ( new_AGEMA_signal_3786 ), .Q ( new_AGEMA_signal_23186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C ( clk ), .D ( new_AGEMA_signal_3787 ), .Q ( new_AGEMA_signal_23190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C ( clk ), .D ( new_AGEMA_signal_3788 ), .Q ( new_AGEMA_signal_23194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C ( clk ), .D ( new_AGEMA_signal_3789 ), .Q ( new_AGEMA_signal_23198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C ( clk ), .D ( new_AGEMA_signal_23205 ), .Q ( new_AGEMA_signal_23206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C ( clk ), .D ( new_AGEMA_signal_23213 ), .Q ( new_AGEMA_signal_23214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C ( clk ), .D ( new_AGEMA_signal_23221 ), .Q ( new_AGEMA_signal_23222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C ( clk ), .D ( new_AGEMA_signal_23229 ), .Q ( new_AGEMA_signal_23230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C ( clk ), .D ( new_AGEMA_signal_23237 ), .Q ( new_AGEMA_signal_23238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_23252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C ( clk ), .D ( new_AGEMA_signal_3522 ), .Q ( new_AGEMA_signal_23258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C ( clk ), .D ( new_AGEMA_signal_3523 ), .Q ( new_AGEMA_signal_23264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C ( clk ), .D ( new_AGEMA_signal_3524 ), .Q ( new_AGEMA_signal_23270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C ( clk ), .D ( new_AGEMA_signal_3525 ), .Q ( new_AGEMA_signal_23276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_23282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C ( clk ), .D ( new_AGEMA_signal_3526 ), .Q ( new_AGEMA_signal_23288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C ( clk ), .D ( new_AGEMA_signal_3527 ), .Q ( new_AGEMA_signal_23294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C ( clk ), .D ( new_AGEMA_signal_3528 ), .Q ( new_AGEMA_signal_23300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C ( clk ), .D ( new_AGEMA_signal_3529 ), .Q ( new_AGEMA_signal_23306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_23312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C ( clk ), .D ( new_AGEMA_signal_3114 ), .Q ( new_AGEMA_signal_23318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C ( clk ), .D ( new_AGEMA_signal_3115 ), .Q ( new_AGEMA_signal_23324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C ( clk ), .D ( new_AGEMA_signal_3116 ), .Q ( new_AGEMA_signal_23330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C ( clk ), .D ( new_AGEMA_signal_3117 ), .Q ( new_AGEMA_signal_23336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C ( clk ), .D ( new_AGEMA_signal_23363 ), .Q ( new_AGEMA_signal_23364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C ( clk ), .D ( new_AGEMA_signal_23371 ), .Q ( new_AGEMA_signal_23372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C ( clk ), .D ( new_AGEMA_signal_23379 ), .Q ( new_AGEMA_signal_23380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C ( clk ), .D ( new_AGEMA_signal_23387 ), .Q ( new_AGEMA_signal_23388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C ( clk ), .D ( new_AGEMA_signal_23395 ), .Q ( new_AGEMA_signal_23396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_23402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C ( clk ), .D ( new_AGEMA_signal_3566 ), .Q ( new_AGEMA_signal_23408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C ( clk ), .D ( new_AGEMA_signal_3567 ), .Q ( new_AGEMA_signal_23414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C ( clk ), .D ( new_AGEMA_signal_3568 ), .Q ( new_AGEMA_signal_23420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C ( clk ), .D ( new_AGEMA_signal_3569 ), .Q ( new_AGEMA_signal_23426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C ( clk ), .D ( new_AGEMA_signal_23453 ), .Q ( new_AGEMA_signal_23454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C ( clk ), .D ( new_AGEMA_signal_23461 ), .Q ( new_AGEMA_signal_23462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C ( clk ), .D ( new_AGEMA_signal_23469 ), .Q ( new_AGEMA_signal_23470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C ( clk ), .D ( new_AGEMA_signal_23477 ), .Q ( new_AGEMA_signal_23478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C ( clk ), .D ( new_AGEMA_signal_23485 ), .Q ( new_AGEMA_signal_23486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C ( clk ), .D ( new_AGEMA_signal_23493 ), .Q ( new_AGEMA_signal_23494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C ( clk ), .D ( new_AGEMA_signal_23501 ), .Q ( new_AGEMA_signal_23502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C ( clk ), .D ( new_AGEMA_signal_23509 ), .Q ( new_AGEMA_signal_23510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C ( clk ), .D ( new_AGEMA_signal_23517 ), .Q ( new_AGEMA_signal_23518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C ( clk ), .D ( new_AGEMA_signal_23525 ), .Q ( new_AGEMA_signal_23526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C ( clk ), .D ( new_AGEMA_signal_23535 ), .Q ( new_AGEMA_signal_23536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C ( clk ), .D ( new_AGEMA_signal_23545 ), .Q ( new_AGEMA_signal_23546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C ( clk ), .D ( new_AGEMA_signal_23555 ), .Q ( new_AGEMA_signal_23556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C ( clk ), .D ( new_AGEMA_signal_23565 ), .Q ( new_AGEMA_signal_23566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C ( clk ), .D ( new_AGEMA_signal_23575 ), .Q ( new_AGEMA_signal_23576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C ( clk ), .D ( new_AGEMA_signal_23583 ), .Q ( new_AGEMA_signal_23584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C ( clk ), .D ( new_AGEMA_signal_23591 ), .Q ( new_AGEMA_signal_23592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C ( clk ), .D ( new_AGEMA_signal_23599 ), .Q ( new_AGEMA_signal_23600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C ( clk ), .D ( new_AGEMA_signal_23607 ), .Q ( new_AGEMA_signal_23608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C ( clk ), .D ( new_AGEMA_signal_23615 ), .Q ( new_AGEMA_signal_23616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_23622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C ( clk ), .D ( new_AGEMA_signal_3646 ), .Q ( new_AGEMA_signal_23628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C ( clk ), .D ( new_AGEMA_signal_3647 ), .Q ( new_AGEMA_signal_23634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C ( clk ), .D ( new_AGEMA_signal_3648 ), .Q ( new_AGEMA_signal_23640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C ( clk ), .D ( new_AGEMA_signal_3649 ), .Q ( new_AGEMA_signal_23646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_23672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C ( clk ), .D ( new_AGEMA_signal_3662 ), .Q ( new_AGEMA_signal_23678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C ( clk ), .D ( new_AGEMA_signal_3663 ), .Q ( new_AGEMA_signal_23684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C ( clk ), .D ( new_AGEMA_signal_3664 ), .Q ( new_AGEMA_signal_23690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C ( clk ), .D ( new_AGEMA_signal_3665 ), .Q ( new_AGEMA_signal_23696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C ( clk ), .D ( new_AGEMA_signal_23703 ), .Q ( new_AGEMA_signal_23704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C ( clk ), .D ( new_AGEMA_signal_23711 ), .Q ( new_AGEMA_signal_23712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C ( clk ), .D ( new_AGEMA_signal_23719 ), .Q ( new_AGEMA_signal_23720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C ( clk ), .D ( new_AGEMA_signal_23727 ), .Q ( new_AGEMA_signal_23728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C ( clk ), .D ( new_AGEMA_signal_23735 ), .Q ( new_AGEMA_signal_23736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_23742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C ( clk ), .D ( new_AGEMA_signal_3718 ), .Q ( new_AGEMA_signal_23748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C ( clk ), .D ( new_AGEMA_signal_3719 ), .Q ( new_AGEMA_signal_23754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C ( clk ), .D ( new_AGEMA_signal_3720 ), .Q ( new_AGEMA_signal_23760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C ( clk ), .D ( new_AGEMA_signal_3721 ), .Q ( new_AGEMA_signal_23766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C ( clk ), .D ( new_AGEMA_signal_23783 ), .Q ( new_AGEMA_signal_23784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C ( clk ), .D ( new_AGEMA_signal_23791 ), .Q ( new_AGEMA_signal_23792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C ( clk ), .D ( new_AGEMA_signal_23799 ), .Q ( new_AGEMA_signal_23800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C ( clk ), .D ( new_AGEMA_signal_23807 ), .Q ( new_AGEMA_signal_23808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C ( clk ), .D ( new_AGEMA_signal_23815 ), .Q ( new_AGEMA_signal_23816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_23842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C ( clk ), .D ( new_AGEMA_signal_3794 ), .Q ( new_AGEMA_signal_23848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C ( clk ), .D ( new_AGEMA_signal_3795 ), .Q ( new_AGEMA_signal_23854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C ( clk ), .D ( new_AGEMA_signal_3796 ), .Q ( new_AGEMA_signal_23860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C ( clk ), .D ( new_AGEMA_signal_3797 ), .Q ( new_AGEMA_signal_23866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_23872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C ( clk ), .D ( new_AGEMA_signal_3802 ), .Q ( new_AGEMA_signal_23878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C ( clk ), .D ( new_AGEMA_signal_3803 ), .Q ( new_AGEMA_signal_23884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C ( clk ), .D ( new_AGEMA_signal_3804 ), .Q ( new_AGEMA_signal_23890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C ( clk ), .D ( new_AGEMA_signal_3805 ), .Q ( new_AGEMA_signal_23896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C ( clk ), .D ( new_AGEMA_signal_24003 ), .Q ( new_AGEMA_signal_24004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C ( clk ), .D ( new_AGEMA_signal_24013 ), .Q ( new_AGEMA_signal_24014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C ( clk ), .D ( new_AGEMA_signal_24023 ), .Q ( new_AGEMA_signal_24024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C ( clk ), .D ( new_AGEMA_signal_24033 ), .Q ( new_AGEMA_signal_24034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C ( clk ), .D ( new_AGEMA_signal_24043 ), .Q ( new_AGEMA_signal_24044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_24152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C ( clk ), .D ( new_AGEMA_signal_3278 ), .Q ( new_AGEMA_signal_24160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C ( clk ), .D ( new_AGEMA_signal_3279 ), .Q ( new_AGEMA_signal_24168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C ( clk ), .D ( new_AGEMA_signal_3280 ), .Q ( new_AGEMA_signal_24176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C ( clk ), .D ( new_AGEMA_signal_3281 ), .Q ( new_AGEMA_signal_24184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C ( clk ), .D ( new_AGEMA_signal_20623 ), .Q ( new_AGEMA_signal_24222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C ( clk ), .D ( new_AGEMA_signal_20625 ), .Q ( new_AGEMA_signal_24230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C ( clk ), .D ( new_AGEMA_signal_20627 ), .Q ( new_AGEMA_signal_24238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C ( clk ), .D ( new_AGEMA_signal_20629 ), .Q ( new_AGEMA_signal_24246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C ( clk ), .D ( new_AGEMA_signal_20631 ), .Q ( new_AGEMA_signal_24254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_24262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C ( clk ), .D ( new_AGEMA_signal_3722 ), .Q ( new_AGEMA_signal_24270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C ( clk ), .D ( new_AGEMA_signal_3723 ), .Q ( new_AGEMA_signal_24278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C ( clk ), .D ( new_AGEMA_signal_3724 ), .Q ( new_AGEMA_signal_24286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C ( clk ), .D ( new_AGEMA_signal_3725 ), .Q ( new_AGEMA_signal_24294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_24352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C ( clk ), .D ( new_AGEMA_signal_3798 ), .Q ( new_AGEMA_signal_24360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C ( clk ), .D ( new_AGEMA_signal_3799 ), .Q ( new_AGEMA_signal_24368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C ( clk ), .D ( new_AGEMA_signal_3800 ), .Q ( new_AGEMA_signal_24376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C ( clk ), .D ( new_AGEMA_signal_3801 ), .Q ( new_AGEMA_signal_24384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7679 ( .C ( clk ), .D ( new_AGEMA_signal_24453 ), .Q ( new_AGEMA_signal_24454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7691 ( .C ( clk ), .D ( new_AGEMA_signal_24465 ), .Q ( new_AGEMA_signal_24466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7703 ( .C ( clk ), .D ( new_AGEMA_signal_24477 ), .Q ( new_AGEMA_signal_24478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7715 ( .C ( clk ), .D ( new_AGEMA_signal_24489 ), .Q ( new_AGEMA_signal_24490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7727 ( .C ( clk ), .D ( new_AGEMA_signal_24501 ), .Q ( new_AGEMA_signal_24502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7741 ( .C ( clk ), .D ( new_AGEMA_signal_24515 ), .Q ( new_AGEMA_signal_24516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7755 ( .C ( clk ), .D ( new_AGEMA_signal_24529 ), .Q ( new_AGEMA_signal_24530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7769 ( .C ( clk ), .D ( new_AGEMA_signal_24543 ), .Q ( new_AGEMA_signal_24544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7783 ( .C ( clk ), .D ( new_AGEMA_signal_24557 ), .Q ( new_AGEMA_signal_24558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7797 ( .C ( clk ), .D ( new_AGEMA_signal_24571 ), .Q ( new_AGEMA_signal_24572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7851 ( .C ( clk ), .D ( new_AGEMA_signal_24625 ), .Q ( new_AGEMA_signal_24626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7865 ( .C ( clk ), .D ( new_AGEMA_signal_24639 ), .Q ( new_AGEMA_signal_24640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7879 ( .C ( clk ), .D ( new_AGEMA_signal_24653 ), .Q ( new_AGEMA_signal_24654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7893 ( .C ( clk ), .D ( new_AGEMA_signal_24667 ), .Q ( new_AGEMA_signal_24668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7907 ( .C ( clk ), .D ( new_AGEMA_signal_24681 ), .Q ( new_AGEMA_signal_24682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8031 ( .C ( clk ), .D ( new_AGEMA_signal_24805 ), .Q ( new_AGEMA_signal_24806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8047 ( .C ( clk ), .D ( new_AGEMA_signal_24821 ), .Q ( new_AGEMA_signal_24822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8063 ( .C ( clk ), .D ( new_AGEMA_signal_24837 ), .Q ( new_AGEMA_signal_24838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8079 ( .C ( clk ), .D ( new_AGEMA_signal_24853 ), .Q ( new_AGEMA_signal_24854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8095 ( .C ( clk ), .D ( new_AGEMA_signal_24869 ), .Q ( new_AGEMA_signal_24870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8141 ( .C ( clk ), .D ( new_AGEMA_signal_24915 ), .Q ( new_AGEMA_signal_24916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8157 ( .C ( clk ), .D ( new_AGEMA_signal_24931 ), .Q ( new_AGEMA_signal_24932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8173 ( .C ( clk ), .D ( new_AGEMA_signal_24947 ), .Q ( new_AGEMA_signal_24948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8189 ( .C ( clk ), .D ( new_AGEMA_signal_24963 ), .Q ( new_AGEMA_signal_24964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8205 ( .C ( clk ), .D ( new_AGEMA_signal_24979 ), .Q ( new_AGEMA_signal_24980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8389 ( .C ( clk ), .D ( new_AGEMA_signal_25163 ), .Q ( new_AGEMA_signal_25164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8405 ( .C ( clk ), .D ( new_AGEMA_signal_25179 ), .Q ( new_AGEMA_signal_25180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8421 ( .C ( clk ), .D ( new_AGEMA_signal_25195 ), .Q ( new_AGEMA_signal_25196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8437 ( .C ( clk ), .D ( new_AGEMA_signal_25211 ), .Q ( new_AGEMA_signal_25212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8453 ( .C ( clk ), .D ( new_AGEMA_signal_25227 ), .Q ( new_AGEMA_signal_25228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8521 ( .C ( clk ), .D ( new_AGEMA_signal_25295 ), .Q ( new_AGEMA_signal_25296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8539 ( .C ( clk ), .D ( new_AGEMA_signal_25313 ), .Q ( new_AGEMA_signal_25314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8557 ( .C ( clk ), .D ( new_AGEMA_signal_25331 ), .Q ( new_AGEMA_signal_25332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8575 ( .C ( clk ), .D ( new_AGEMA_signal_25349 ), .Q ( new_AGEMA_signal_25350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8593 ( .C ( clk ), .D ( new_AGEMA_signal_25367 ), .Q ( new_AGEMA_signal_25368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8771 ( .C ( clk ), .D ( new_AGEMA_signal_25545 ), .Q ( new_AGEMA_signal_25546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8791 ( .C ( clk ), .D ( new_AGEMA_signal_25565 ), .Q ( new_AGEMA_signal_25566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8811 ( .C ( clk ), .D ( new_AGEMA_signal_25585 ), .Q ( new_AGEMA_signal_25586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8831 ( .C ( clk ), .D ( new_AGEMA_signal_25605 ), .Q ( new_AGEMA_signal_25606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8851 ( .C ( clk ), .D ( new_AGEMA_signal_25625 ), .Q ( new_AGEMA_signal_25626 ) ) ;

    /* cells in depth 12 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2001 ( .ina ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, n1932}), .inb ({new_AGEMA_signal_20431, new_AGEMA_signal_20427, new_AGEMA_signal_20423, new_AGEMA_signal_20419, new_AGEMA_signal_20415}), .clk ( clk ), .rnd ({Fresh[9914], Fresh[9913], Fresh[9912], Fresh[9911], Fresh[9910], Fresh[9909], Fresh[9908], Fresh[9907], Fresh[9906], Fresh[9905], Fresh[9904], Fresh[9903], Fresh[9902], Fresh[9901], Fresh[9900]}), .outt ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, n1933}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2051 ( .ina ({new_AGEMA_signal_20451, new_AGEMA_signal_20447, new_AGEMA_signal_20443, new_AGEMA_signal_20439, new_AGEMA_signal_20435}), .inb ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, n1955}), .clk ( clk ), .rnd ({Fresh[9929], Fresh[9928], Fresh[9927], Fresh[9926], Fresh[9925], Fresh[9924], Fresh[9923], Fresh[9922], Fresh[9921], Fresh[9920], Fresh[9919], Fresh[9918], Fresh[9917], Fresh[9916], Fresh[9915]}), .outt ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, n1958}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2067 ( .ina ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n1967}), .inb ({new_AGEMA_signal_20491, new_AGEMA_signal_20483, new_AGEMA_signal_20475, new_AGEMA_signal_20467, new_AGEMA_signal_20459}), .clk ( clk ), .rnd ({Fresh[9944], Fresh[9943], Fresh[9942], Fresh[9941], Fresh[9940], Fresh[9939], Fresh[9938], Fresh[9937], Fresh[9936], Fresh[9935], Fresh[9934], Fresh[9933], Fresh[9932], Fresh[9931], Fresh[9930]}), .outt ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n1990}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2104 ( .ina ({new_AGEMA_signal_20501, new_AGEMA_signal_20499, new_AGEMA_signal_20497, new_AGEMA_signal_20495, new_AGEMA_signal_20493}), .inb ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, new_AGEMA_signal_3542, n1977}), .clk ( clk ), .rnd ({Fresh[9959], Fresh[9958], Fresh[9957], Fresh[9956], Fresh[9955], Fresh[9954], Fresh[9953], Fresh[9952], Fresh[9951], Fresh[9950], Fresh[9949], Fresh[9948], Fresh[9947], Fresh[9946], Fresh[9945]}), .outt ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, new_AGEMA_signal_3854, n1982}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2128 ( .ina ({new_AGEMA_signal_20541, new_AGEMA_signal_20533, new_AGEMA_signal_20525, new_AGEMA_signal_20517, new_AGEMA_signal_20509}), .inb ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, n1998}), .clk ( clk ), .rnd ({Fresh[9974], Fresh[9973], Fresh[9972], Fresh[9971], Fresh[9970], Fresh[9969], Fresh[9968], Fresh[9967], Fresh[9966], Fresh[9965], Fresh[9964], Fresh[9963], Fresh[9962], Fresh[9961], Fresh[9960]}), .outt ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, n1999}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2148 ( .ina ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, n2010}), .inb ({new_AGEMA_signal_20571, new_AGEMA_signal_20565, new_AGEMA_signal_20559, new_AGEMA_signal_20553, new_AGEMA_signal_20547}), .clk ( clk ), .rnd ({Fresh[9989], Fresh[9988], Fresh[9987], Fresh[9986], Fresh[9985], Fresh[9984], Fresh[9983], Fresh[9982], Fresh[9981], Fresh[9980], Fresh[9979], Fresh[9978], Fresh[9977], Fresh[9976], Fresh[9975]}), .outt ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, new_AGEMA_signal_3863, new_AGEMA_signal_3862, n2011}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2165 ( .ina ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, n2024}), .inb ({new_AGEMA_signal_20591, new_AGEMA_signal_20587, new_AGEMA_signal_20583, new_AGEMA_signal_20579, new_AGEMA_signal_20575}), .clk ( clk ), .rnd ({Fresh[10004], Fresh[10003], Fresh[10002], Fresh[10001], Fresh[10000], Fresh[9999], Fresh[9998], Fresh[9997], Fresh[9996], Fresh[9995], Fresh[9994], Fresh[9993], Fresh[9992], Fresh[9991], Fresh[9990]}), .outt ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2025}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2179 ( .ina ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, n2035}), .inb ({new_AGEMA_signal_20621, new_AGEMA_signal_20615, new_AGEMA_signal_20609, new_AGEMA_signal_20603, new_AGEMA_signal_20597}), .clk ( clk ), .rnd ({Fresh[10019], Fresh[10018], Fresh[10017], Fresh[10016], Fresh[10015], Fresh[10014], Fresh[10013], Fresh[10012], Fresh[10011], Fresh[10010], Fresh[10009], Fresh[10008], Fresh[10007], Fresh[10006], Fresh[10005]}), .outt ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, n2036}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2196 ( .ina ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2048}), .inb ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, n2047}), .clk ( clk ), .rnd ({Fresh[10034], Fresh[10033], Fresh[10032], Fresh[10031], Fresh[10030], Fresh[10029], Fresh[10028], Fresh[10027], Fresh[10026], Fresh[10025], Fresh[10024], Fresh[10023], Fresh[10022], Fresh[10021], Fresh[10020]}), .outt ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, new_AGEMA_signal_3875, new_AGEMA_signal_3874, n2049}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2207 ( .ina ({new_AGEMA_signal_20631, new_AGEMA_signal_20629, new_AGEMA_signal_20627, new_AGEMA_signal_20625, new_AGEMA_signal_20623}), .inb ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, new_AGEMA_signal_3578, n2059}), .clk ( clk ), .rnd ({Fresh[10049], Fresh[10048], Fresh[10047], Fresh[10046], Fresh[10045], Fresh[10044], Fresh[10043], Fresh[10042], Fresh[10041], Fresh[10040], Fresh[10039], Fresh[10038], Fresh[10037], Fresh[10036], Fresh[10035]}), .outt ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, new_AGEMA_signal_3879, new_AGEMA_signal_3878, n2072}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2214 ( .ina ({new_AGEMA_signal_20661, new_AGEMA_signal_20655, new_AGEMA_signal_20649, new_AGEMA_signal_20643, new_AGEMA_signal_20637}), .inb ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2064}), .clk ( clk ), .rnd ({Fresh[10064], Fresh[10063], Fresh[10062], Fresh[10061], Fresh[10060], Fresh[10059], Fresh[10058], Fresh[10057], Fresh[10056], Fresh[10055], Fresh[10054], Fresh[10053], Fresh[10052], Fresh[10051], Fresh[10050]}), .outt ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, n2067}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2230 ( .ina ({new_AGEMA_signal_20691, new_AGEMA_signal_20685, new_AGEMA_signal_20679, new_AGEMA_signal_20673, new_AGEMA_signal_20667}), .inb ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, n2077}), .clk ( clk ), .rnd ({Fresh[10079], Fresh[10078], Fresh[10077], Fresh[10076], Fresh[10075], Fresh[10074], Fresh[10073], Fresh[10072], Fresh[10071], Fresh[10070], Fresh[10069], Fresh[10068], Fresh[10067], Fresh[10066], Fresh[10065]}), .outt ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3887, new_AGEMA_signal_3886, n2078}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2250 ( .ina ({new_AGEMA_signal_20701, new_AGEMA_signal_20699, new_AGEMA_signal_20697, new_AGEMA_signal_20695, new_AGEMA_signal_20693}), .inb ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, n2158}), .clk ( clk ), .rnd ({Fresh[10094], Fresh[10093], Fresh[10092], Fresh[10091], Fresh[10090], Fresh[10089], Fresh[10088], Fresh[10087], Fresh[10086], Fresh[10085], Fresh[10084], Fresh[10083], Fresh[10082], Fresh[10081], Fresh[10080]}), .outt ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, new_AGEMA_signal_3890, n2097}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2257 ( .ina ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2095}), .inb ({new_AGEMA_signal_20721, new_AGEMA_signal_20717, new_AGEMA_signal_20713, new_AGEMA_signal_20709, new_AGEMA_signal_20705}), .clk ( clk ), .rnd ({Fresh[10109], Fresh[10108], Fresh[10107], Fresh[10106], Fresh[10105], Fresh[10104], Fresh[10103], Fresh[10102], Fresh[10101], Fresh[10100], Fresh[10099], Fresh[10098], Fresh[10097], Fresh[10096], Fresh[10095]}), .outt ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, n2096}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2275 ( .ina ({new_AGEMA_signal_20751, new_AGEMA_signal_20745, new_AGEMA_signal_20739, new_AGEMA_signal_20733, new_AGEMA_signal_20727}), .inb ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, new_AGEMA_signal_3899, new_AGEMA_signal_3898, n2117}), .clk ( clk ), .rnd ({Fresh[10124], Fresh[10123], Fresh[10122], Fresh[10121], Fresh[10120], Fresh[10119], Fresh[10118], Fresh[10117], Fresh[10116], Fresh[10115], Fresh[10114], Fresh[10113], Fresh[10112], Fresh[10111], Fresh[10110]}), .outt ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, new_AGEMA_signal_4115, new_AGEMA_signal_4114, n2128}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2285 ( .ina ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, n2123}), .inb ({new_AGEMA_signal_20781, new_AGEMA_signal_20775, new_AGEMA_signal_20769, new_AGEMA_signal_20763, new_AGEMA_signal_20757}), .clk ( clk ), .rnd ({Fresh[10139], Fresh[10138], Fresh[10137], Fresh[10136], Fresh[10135], Fresh[10134], Fresh[10133], Fresh[10132], Fresh[10131], Fresh[10130], Fresh[10129], Fresh[10128], Fresh[10127], Fresh[10126], Fresh[10125]}), .outt ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, new_AGEMA_signal_3902, n2124}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2301 ( .ina ({new_AGEMA_signal_20791, new_AGEMA_signal_20789, new_AGEMA_signal_20787, new_AGEMA_signal_20785, new_AGEMA_signal_20783}), .inb ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, n2135}), .clk ( clk ), .rnd ({Fresh[10154], Fresh[10153], Fresh[10152], Fresh[10151], Fresh[10150], Fresh[10149], Fresh[10148], Fresh[10147], Fresh[10146], Fresh[10145], Fresh[10144], Fresh[10143], Fresh[10142], Fresh[10141], Fresh[10140]}), .outt ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2148}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2310 ( .ina ({new_AGEMA_signal_20821, new_AGEMA_signal_20815, new_AGEMA_signal_20809, new_AGEMA_signal_20803, new_AGEMA_signal_20797}), .inb ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, n2141}), .clk ( clk ), .rnd ({Fresh[10169], Fresh[10168], Fresh[10167], Fresh[10166], Fresh[10165], Fresh[10164], Fresh[10163], Fresh[10162], Fresh[10161], Fresh[10160], Fresh[10159], Fresh[10158], Fresh[10157], Fresh[10156], Fresh[10155]}), .outt ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, new_AGEMA_signal_3906, n2142}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2325 ( .ina ({new_AGEMA_signal_20831, new_AGEMA_signal_20829, new_AGEMA_signal_20827, new_AGEMA_signal_20825, new_AGEMA_signal_20823}), .inb ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, n2158}), .clk ( clk ), .rnd ({Fresh[10184], Fresh[10183], Fresh[10182], Fresh[10181], Fresh[10180], Fresh[10179], Fresh[10178], Fresh[10177], Fresh[10176], Fresh[10175], Fresh[10174], Fresh[10173], Fresh[10172], Fresh[10171], Fresh[10170]}), .outt ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, new_AGEMA_signal_3911, new_AGEMA_signal_3910, n2168}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2332 ( .ina ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, n2166}), .inb ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2165}), .clk ( clk ), .rnd ({Fresh[10199], Fresh[10198], Fresh[10197], Fresh[10196], Fresh[10195], Fresh[10194], Fresh[10193], Fresh[10192], Fresh[10191], Fresh[10190], Fresh[10189], Fresh[10188], Fresh[10187], Fresh[10186], Fresh[10185]}), .outt ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, n2167}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2347 ( .ina ({new_AGEMA_signal_20851, new_AGEMA_signal_20847, new_AGEMA_signal_20843, new_AGEMA_signal_20839, new_AGEMA_signal_20835}), .inb ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2180}), .clk ( clk ), .rnd ({Fresh[10214], Fresh[10213], Fresh[10212], Fresh[10211], Fresh[10210], Fresh[10209], Fresh[10208], Fresh[10207], Fresh[10206], Fresh[10205], Fresh[10204], Fresh[10203], Fresh[10202], Fresh[10201], Fresh[10200]}), .outt ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, new_AGEMA_signal_3918, n2184}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2361 ( .ina ({new_AGEMA_signal_20871, new_AGEMA_signal_20867, new_AGEMA_signal_20863, new_AGEMA_signal_20859, new_AGEMA_signal_20855}), .inb ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, n2194}), .clk ( clk ), .rnd ({Fresh[10229], Fresh[10228], Fresh[10227], Fresh[10226], Fresh[10225], Fresh[10224], Fresh[10223], Fresh[10222], Fresh[10221], Fresh[10220], Fresh[10219], Fresh[10218], Fresh[10217], Fresh[10216], Fresh[10215]}), .outt ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, n2197}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2373 ( .ina ({new_AGEMA_signal_20881, new_AGEMA_signal_20879, new_AGEMA_signal_20877, new_AGEMA_signal_20875, new_AGEMA_signal_20873}), .inb ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, new_AGEMA_signal_3927, new_AGEMA_signal_3926, n2204}), .clk ( clk ), .rnd ({Fresh[10244], Fresh[10243], Fresh[10242], Fresh[10241], Fresh[10240], Fresh[10239], Fresh[10238], Fresh[10237], Fresh[10236], Fresh[10235], Fresh[10234], Fresh[10233], Fresh[10232], Fresh[10231], Fresh[10230]}), .outt ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, new_AGEMA_signal_4139, new_AGEMA_signal_4138, n2205}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2390 ( .ina ({new_AGEMA_signal_20921, new_AGEMA_signal_20913, new_AGEMA_signal_20905, new_AGEMA_signal_20897, new_AGEMA_signal_20889}), .inb ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2225}), .clk ( clk ), .rnd ({Fresh[10259], Fresh[10258], Fresh[10257], Fresh[10256], Fresh[10255], Fresh[10254], Fresh[10253], Fresh[10252], Fresh[10251], Fresh[10250], Fresh[10249], Fresh[10248], Fresh[10247], Fresh[10246], Fresh[10245]}), .outt ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, new_AGEMA_signal_3930, n2232}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2395 ( .ina ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, n2230}), .inb ({new_AGEMA_signal_20951, new_AGEMA_signal_20945, new_AGEMA_signal_20939, new_AGEMA_signal_20933, new_AGEMA_signal_20927}), .clk ( clk ), .rnd ({Fresh[10274], Fresh[10273], Fresh[10272], Fresh[10271], Fresh[10270], Fresh[10269], Fresh[10268], Fresh[10267], Fresh[10266], Fresh[10265], Fresh[10264], Fresh[10263], Fresh[10262], Fresh[10261], Fresh[10260]}), .outt ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, n2231}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2401 ( .ina ({new_AGEMA_signal_20971, new_AGEMA_signal_20967, new_AGEMA_signal_20963, new_AGEMA_signal_20959, new_AGEMA_signal_20955}), .inb ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, n2236}), .clk ( clk ), .rnd ({Fresh[10289], Fresh[10288], Fresh[10287], Fresh[10286], Fresh[10285], Fresh[10284], Fresh[10283], Fresh[10282], Fresh[10281], Fresh[10280], Fresh[10279], Fresh[10278], Fresh[10277], Fresh[10276], Fresh[10275]}), .outt ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, new_AGEMA_signal_4146, n2239}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2413 ( .ina ({new_AGEMA_signal_20991, new_AGEMA_signal_20987, new_AGEMA_signal_20983, new_AGEMA_signal_20979, new_AGEMA_signal_20975}), .inb ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2247}), .clk ( clk ), .rnd ({Fresh[10304], Fresh[10303], Fresh[10302], Fresh[10301], Fresh[10300], Fresh[10299], Fresh[10298], Fresh[10297], Fresh[10296], Fresh[10295], Fresh[10294], Fresh[10293], Fresh[10292], Fresh[10291], Fresh[10290]}), .outt ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, new_AGEMA_signal_3938, n2250}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2428 ( .ina ({new_AGEMA_signal_20631, new_AGEMA_signal_20629, new_AGEMA_signal_20627, new_AGEMA_signal_20625, new_AGEMA_signal_20623}), .inb ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, n2264}), .clk ( clk ), .rnd ({Fresh[10319], Fresh[10318], Fresh[10317], Fresh[10316], Fresh[10315], Fresh[10314], Fresh[10313], Fresh[10312], Fresh[10311], Fresh[10310], Fresh[10309], Fresh[10308], Fresh[10307], Fresh[10306], Fresh[10305]}), .outt ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, new_AGEMA_signal_3942, n2276}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2439 ( .ina ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2271}), .inb ({new_AGEMA_signal_21001, new_AGEMA_signal_20999, new_AGEMA_signal_20997, new_AGEMA_signal_20995, new_AGEMA_signal_20993}), .clk ( clk ), .rnd ({Fresh[10334], Fresh[10333], Fresh[10332], Fresh[10331], Fresh[10330], Fresh[10329], Fresh[10328], Fresh[10327], Fresh[10326], Fresh[10325], Fresh[10324], Fresh[10323], Fresh[10322], Fresh[10321], Fresh[10320]}), .outt ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, n2272}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2454 ( .ina ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2286}), .inb ({new_AGEMA_signal_21011, new_AGEMA_signal_21009, new_AGEMA_signal_21007, new_AGEMA_signal_21005, new_AGEMA_signal_21003}), .clk ( clk ), .rnd ({Fresh[10349], Fresh[10348], Fresh[10347], Fresh[10346], Fresh[10345], Fresh[10344], Fresh[10343], Fresh[10342], Fresh[10341], Fresh[10340], Fresh[10339], Fresh[10338], Fresh[10337], Fresh[10336], Fresh[10335]}), .outt ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, n2306}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2468 ( .ina ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2295}), .inb ({new_AGEMA_signal_21031, new_AGEMA_signal_21027, new_AGEMA_signal_21023, new_AGEMA_signal_21019, new_AGEMA_signal_21015}), .clk ( clk ), .rnd ({Fresh[10364], Fresh[10363], Fresh[10362], Fresh[10361], Fresh[10360], Fresh[10359], Fresh[10358], Fresh[10357], Fresh[10356], Fresh[10355], Fresh[10354], Fresh[10353], Fresh[10352], Fresh[10351], Fresh[10350]}), .outt ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, n2296}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2489 ( .ina ({new_AGEMA_signal_21051, new_AGEMA_signal_21047, new_AGEMA_signal_21043, new_AGEMA_signal_21039, new_AGEMA_signal_21035}), .inb ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, n2322}), .clk ( clk ), .rnd ({Fresh[10379], Fresh[10378], Fresh[10377], Fresh[10376], Fresh[10375], Fresh[10374], Fresh[10373], Fresh[10372], Fresh[10371], Fresh[10370], Fresh[10369], Fresh[10368], Fresh[10367], Fresh[10366], Fresh[10365]}), .outt ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, new_AGEMA_signal_3954, n2324}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2500 ( .ina ({new_AGEMA_signal_21061, new_AGEMA_signal_21059, new_AGEMA_signal_21057, new_AGEMA_signal_21055, new_AGEMA_signal_21053}), .inb ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, n2333}), .clk ( clk ), .rnd ({Fresh[10394], Fresh[10393], Fresh[10392], Fresh[10391], Fresh[10390], Fresh[10389], Fresh[10388], Fresh[10387], Fresh[10386], Fresh[10385], Fresh[10384], Fresh[10383], Fresh[10382], Fresh[10381], Fresh[10380]}), .outt ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, new_AGEMA_signal_3958, n2337}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2511 ( .ina ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, n2345}), .inb ({new_AGEMA_signal_21091, new_AGEMA_signal_21085, new_AGEMA_signal_21079, new_AGEMA_signal_21073, new_AGEMA_signal_21067}), .clk ( clk ), .rnd ({Fresh[10409], Fresh[10408], Fresh[10407], Fresh[10406], Fresh[10405], Fresh[10404], Fresh[10403], Fresh[10402], Fresh[10401], Fresh[10400], Fresh[10399], Fresh[10398], Fresh[10397], Fresh[10396], Fresh[10395]}), .outt ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, new_AGEMA_signal_3962, n2350}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2528 ( .ina ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, new_AGEMA_signal_3686, n2361}), .inb ({new_AGEMA_signal_21111, new_AGEMA_signal_21107, new_AGEMA_signal_21103, new_AGEMA_signal_21099, new_AGEMA_signal_21095}), .clk ( clk ), .rnd ({Fresh[10424], Fresh[10423], Fresh[10422], Fresh[10421], Fresh[10420], Fresh[10419], Fresh[10418], Fresh[10417], Fresh[10416], Fresh[10415], Fresh[10414], Fresh[10413], Fresh[10412], Fresh[10411], Fresh[10410]}), .outt ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, new_AGEMA_signal_3966, n2362}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2550 ( .ina ({new_AGEMA_signal_21121, new_AGEMA_signal_21119, new_AGEMA_signal_21117, new_AGEMA_signal_21115, new_AGEMA_signal_21113}), .inb ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, new_AGEMA_signal_3338, n2388}), .clk ( clk ), .rnd ({Fresh[10439], Fresh[10438], Fresh[10437], Fresh[10436], Fresh[10435], Fresh[10434], Fresh[10433], Fresh[10432], Fresh[10431], Fresh[10430], Fresh[10429], Fresh[10428], Fresh[10427], Fresh[10426], Fresh[10425]}), .outt ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2389}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2557 ( .ina ({new_AGEMA_signal_21141, new_AGEMA_signal_21137, new_AGEMA_signal_21133, new_AGEMA_signal_21129, new_AGEMA_signal_21125}), .inb ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, n2393}), .clk ( clk ), .rnd ({Fresh[10454], Fresh[10453], Fresh[10452], Fresh[10451], Fresh[10450], Fresh[10449], Fresh[10448], Fresh[10447], Fresh[10446], Fresh[10445], Fresh[10444], Fresh[10443], Fresh[10442], Fresh[10441], Fresh[10440]}), .outt ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, new_AGEMA_signal_3974, n2397}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2568 ( .ina ({new_AGEMA_signal_21161, new_AGEMA_signal_21157, new_AGEMA_signal_21153, new_AGEMA_signal_21149, new_AGEMA_signal_21145}), .inb ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, n2405}), .clk ( clk ), .rnd ({Fresh[10469], Fresh[10468], Fresh[10467], Fresh[10466], Fresh[10465], Fresh[10464], Fresh[10463], Fresh[10462], Fresh[10461], Fresh[10460], Fresh[10459], Fresh[10458], Fresh[10457], Fresh[10456], Fresh[10455]}), .outt ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, n2411}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2580 ( .ina ({new_AGEMA_signal_21181, new_AGEMA_signal_21177, new_AGEMA_signal_21173, new_AGEMA_signal_21169, new_AGEMA_signal_21165}), .inb ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, n2419}), .clk ( clk ), .rnd ({Fresh[10484], Fresh[10483], Fresh[10482], Fresh[10481], Fresh[10480], Fresh[10479], Fresh[10478], Fresh[10477], Fresh[10476], Fresh[10475], Fresh[10474], Fresh[10473], Fresh[10472], Fresh[10471], Fresh[10470]}), .outt ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, n2420}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2593 ( .ina ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2436}), .inb ({new_AGEMA_signal_21191, new_AGEMA_signal_21189, new_AGEMA_signal_21187, new_AGEMA_signal_21185, new_AGEMA_signal_21183}), .clk ( clk ), .rnd ({Fresh[10499], Fresh[10498], Fresh[10497], Fresh[10496], Fresh[10495], Fresh[10494], Fresh[10493], Fresh[10492], Fresh[10491], Fresh[10490], Fresh[10489], Fresh[10488], Fresh[10487], Fresh[10486], Fresh[10485]}), .outt ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, n2440}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2614 ( .ina ({new_AGEMA_signal_21211, new_AGEMA_signal_21207, new_AGEMA_signal_21203, new_AGEMA_signal_21199, new_AGEMA_signal_21195}), .inb ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, n2461}), .clk ( clk ), .rnd ({Fresh[10514], Fresh[10513], Fresh[10512], Fresh[10511], Fresh[10510], Fresh[10509], Fresh[10508], Fresh[10507], Fresh[10506], Fresh[10505], Fresh[10504], Fresh[10503], Fresh[10502], Fresh[10501], Fresh[10500]}), .outt ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, new_AGEMA_signal_3991, new_AGEMA_signal_3990, n2516}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2621 ( .ins ({new_AGEMA_signal_21221, new_AGEMA_signal_21219, new_AGEMA_signal_21217, new_AGEMA_signal_21215, new_AGEMA_signal_21213}), .inb ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, n2469}), .ina ({new_AGEMA_signal_21251, new_AGEMA_signal_21245, new_AGEMA_signal_21239, new_AGEMA_signal_21233, new_AGEMA_signal_21227}), .clk ( clk ), .rnd ({Fresh[10529], Fresh[10528], Fresh[10527], Fresh[10526], Fresh[10525], Fresh[10524], Fresh[10523], Fresh[10522], Fresh[10521], Fresh[10520], Fresh[10519], Fresh[10518], Fresh[10517], Fresh[10516], Fresh[10515]}), .outt ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, new_AGEMA_signal_3731, new_AGEMA_signal_3730, n2471}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2636 ( .ina ({new_AGEMA_signal_21281, new_AGEMA_signal_21275, new_AGEMA_signal_21269, new_AGEMA_signal_21263, new_AGEMA_signal_21257}), .inb ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, new_AGEMA_signal_3734, n2484}), .clk ( clk ), .rnd ({Fresh[10544], Fresh[10543], Fresh[10542], Fresh[10541], Fresh[10540], Fresh[10539], Fresh[10538], Fresh[10537], Fresh[10536], Fresh[10535], Fresh[10534], Fresh[10533], Fresh[10532], Fresh[10531], Fresh[10530]}), .outt ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, new_AGEMA_signal_3998, n2485}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2644 ( .ina ({new_AGEMA_signal_20661, new_AGEMA_signal_20655, new_AGEMA_signal_20649, new_AGEMA_signal_20643, new_AGEMA_signal_20637}), .inb ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, n2491}), .clk ( clk ), .rnd ({Fresh[10559], Fresh[10558], Fresh[10557], Fresh[10556], Fresh[10555], Fresh[10554], Fresh[10553], Fresh[10552], Fresh[10551], Fresh[10550], Fresh[10549], Fresh[10548], Fresh[10547], Fresh[10546], Fresh[10545]}), .outt ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, n2502}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2651 ( .ina ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, new_AGEMA_signal_3743, new_AGEMA_signal_3742, n2500}), .inb ({new_AGEMA_signal_21301, new_AGEMA_signal_21297, new_AGEMA_signal_21293, new_AGEMA_signal_21289, new_AGEMA_signal_21285}), .clk ( clk ), .rnd ({Fresh[10574], Fresh[10573], Fresh[10572], Fresh[10571], Fresh[10570], Fresh[10569], Fresh[10568], Fresh[10567], Fresh[10566], Fresh[10565], Fresh[10564], Fresh[10563], Fresh[10562], Fresh[10561], Fresh[10560]}), .outt ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, new_AGEMA_signal_4003, new_AGEMA_signal_4002, n2501}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2657 ( .ina ({new_AGEMA_signal_21181, new_AGEMA_signal_21177, new_AGEMA_signal_21173, new_AGEMA_signal_21169, new_AGEMA_signal_21165}), .inb ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, new_AGEMA_signal_4007, new_AGEMA_signal_4006, n2508}), .clk ( clk ), .rnd ({Fresh[10589], Fresh[10588], Fresh[10587], Fresh[10586], Fresh[10585], Fresh[10584], Fresh[10583], Fresh[10582], Fresh[10581], Fresh[10580], Fresh[10579], Fresh[10578], Fresh[10577], Fresh[10576], Fresh[10575]}), .outt ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, new_AGEMA_signal_4203, new_AGEMA_signal_4202, n2509}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2671 ( .ina ({new_AGEMA_signal_21311, new_AGEMA_signal_21309, new_AGEMA_signal_21307, new_AGEMA_signal_21305, new_AGEMA_signal_21303}), .inb ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, new_AGEMA_signal_4010, n2526}), .clk ( clk ), .rnd ({Fresh[10604], Fresh[10603], Fresh[10602], Fresh[10601], Fresh[10600], Fresh[10599], Fresh[10598], Fresh[10597], Fresh[10596], Fresh[10595], Fresh[10594], Fresh[10593], Fresh[10592], Fresh[10591], Fresh[10590]}), .outt ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, new_AGEMA_signal_4206, n2527}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2680 ( .ina ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, new_AGEMA_signal_3755, new_AGEMA_signal_3754, n2539}), .inb ({new_AGEMA_signal_21351, new_AGEMA_signal_21343, new_AGEMA_signal_21335, new_AGEMA_signal_21327, new_AGEMA_signal_21319}), .clk ( clk ), .rnd ({Fresh[10619], Fresh[10618], Fresh[10617], Fresh[10616], Fresh[10615], Fresh[10614], Fresh[10613], Fresh[10612], Fresh[10611], Fresh[10610], Fresh[10609], Fresh[10608], Fresh[10607], Fresh[10606], Fresh[10605]}), .outt ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, new_AGEMA_signal_4015, new_AGEMA_signal_4014, n2550}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2685 ( .ina ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, new_AGEMA_signal_3758, n2548}), .inb ({new_AGEMA_signal_21361, new_AGEMA_signal_21359, new_AGEMA_signal_21357, new_AGEMA_signal_21355, new_AGEMA_signal_21353}), .clk ( clk ), .rnd ({Fresh[10634], Fresh[10633], Fresh[10632], Fresh[10631], Fresh[10630], Fresh[10629], Fresh[10628], Fresh[10627], Fresh[10626], Fresh[10625], Fresh[10624], Fresh[10623], Fresh[10622], Fresh[10621], Fresh[10620]}), .outt ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, new_AGEMA_signal_4019, new_AGEMA_signal_4018, n2549}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2701 ( .ina ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, n2568}), .inb ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, new_AGEMA_signal_3767, new_AGEMA_signal_3766, n2567}), .clk ( clk ), .rnd ({Fresh[10649], Fresh[10648], Fresh[10647], Fresh[10646], Fresh[10645], Fresh[10644], Fresh[10643], Fresh[10642], Fresh[10641], Fresh[10640], Fresh[10639], Fresh[10638], Fresh[10637], Fresh[10636], Fresh[10635]}), .outt ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, n2569}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2712 ( .ina ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3770, n2583}), .inb ({new_AGEMA_signal_21381, new_AGEMA_signal_21377, new_AGEMA_signal_21373, new_AGEMA_signal_21369, new_AGEMA_signal_21365}), .clk ( clk ), .rnd ({Fresh[10664], Fresh[10663], Fresh[10662], Fresh[10661], Fresh[10660], Fresh[10659], Fresh[10658], Fresh[10657], Fresh[10656], Fresh[10655], Fresh[10654], Fresh[10653], Fresh[10652], Fresh[10651], Fresh[10650]}), .outt ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, n2584}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2729 ( .ina ({new_AGEMA_signal_21401, new_AGEMA_signal_21397, new_AGEMA_signal_21393, new_AGEMA_signal_21389, new_AGEMA_signal_21385}), .inb ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2604}), .clk ( clk ), .rnd ({Fresh[10679], Fresh[10678], Fresh[10677], Fresh[10676], Fresh[10675], Fresh[10674], Fresh[10673], Fresh[10672], Fresh[10671], Fresh[10670], Fresh[10669], Fresh[10668], Fresh[10667], Fresh[10666], Fresh[10665]}), .outt ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, n2606}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2740 ( .ina ({new_AGEMA_signal_20661, new_AGEMA_signal_20655, new_AGEMA_signal_20649, new_AGEMA_signal_20643, new_AGEMA_signal_20637}), .inb ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, new_AGEMA_signal_3779, new_AGEMA_signal_3778, n2621}), .clk ( clk ), .rnd ({Fresh[10694], Fresh[10693], Fresh[10692], Fresh[10691], Fresh[10690], Fresh[10689], Fresh[10688], Fresh[10687], Fresh[10686], Fresh[10685], Fresh[10684], Fresh[10683], Fresh[10682], Fresh[10681], Fresh[10680]}), .outt ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, new_AGEMA_signal_4035, new_AGEMA_signal_4034, n2622}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2747 ( .ina ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, new_AGEMA_signal_3783, new_AGEMA_signal_3782, n2633}), .inb ({new_AGEMA_signal_21421, new_AGEMA_signal_21417, new_AGEMA_signal_21413, new_AGEMA_signal_21409, new_AGEMA_signal_21405}), .clk ( clk ), .rnd ({Fresh[10709], Fresh[10708], Fresh[10707], Fresh[10706], Fresh[10705], Fresh[10704], Fresh[10703], Fresh[10702], Fresh[10701], Fresh[10700], Fresh[10699], Fresh[10698], Fresh[10697], Fresh[10696], Fresh[10695]}), .outt ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, n2634}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2761 ( .ina ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_3791, new_AGEMA_signal_3790, n2656}), .inb ({new_AGEMA_signal_21441, new_AGEMA_signal_21437, new_AGEMA_signal_21433, new_AGEMA_signal_21429, new_AGEMA_signal_21425}), .clk ( clk ), .rnd ({Fresh[10724], Fresh[10723], Fresh[10722], Fresh[10721], Fresh[10720], Fresh[10719], Fresh[10718], Fresh[10717], Fresh[10716], Fresh[10715], Fresh[10714], Fresh[10713], Fresh[10712], Fresh[10711], Fresh[10710]}), .outt ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, new_AGEMA_signal_4043, new_AGEMA_signal_4042, n2657}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2783 ( .ina ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, new_AGEMA_signal_3807, new_AGEMA_signal_3806, n2696}), .inb ({new_AGEMA_signal_21461, new_AGEMA_signal_21457, new_AGEMA_signal_21453, new_AGEMA_signal_21449, new_AGEMA_signal_21445}), .clk ( clk ), .rnd ({Fresh[10739], Fresh[10738], Fresh[10737], Fresh[10736], Fresh[10735], Fresh[10734], Fresh[10733], Fresh[10732], Fresh[10731], Fresh[10730], Fresh[10729], Fresh[10728], Fresh[10727], Fresh[10726], Fresh[10725]}), .outt ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, new_AGEMA_signal_4047, new_AGEMA_signal_4046, n2697}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2795 ( .ina ({new_AGEMA_signal_20631, new_AGEMA_signal_20629, new_AGEMA_signal_20627, new_AGEMA_signal_20625, new_AGEMA_signal_20623}), .inb ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, n2718}), .clk ( clk ), .rnd ({Fresh[10754], Fresh[10753], Fresh[10752], Fresh[10751], Fresh[10750], Fresh[10749], Fresh[10748], Fresh[10747], Fresh[10746], Fresh[10745], Fresh[10744], Fresh[10743], Fresh[10742], Fresh[10741], Fresh[10740]}), .outt ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, new_AGEMA_signal_4051, new_AGEMA_signal_4050, n2808}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2802 ( .ina ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, new_AGEMA_signal_3815, new_AGEMA_signal_3814, n2730}), .inb ({new_AGEMA_signal_21501, new_AGEMA_signal_21493, new_AGEMA_signal_21485, new_AGEMA_signal_21477, new_AGEMA_signal_21469}), .clk ( clk ), .rnd ({Fresh[10769], Fresh[10768], Fresh[10767], Fresh[10766], Fresh[10765], Fresh[10764], Fresh[10763], Fresh[10762], Fresh[10761], Fresh[10760], Fresh[10759], Fresh[10758], Fresh[10757], Fresh[10756], Fresh[10755]}), .outt ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, new_AGEMA_signal_4055, new_AGEMA_signal_4054, n2747}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2810 ( .ina ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, new_AGEMA_signal_3819, new_AGEMA_signal_3818, n2745}), .inb ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, n2744}), .clk ( clk ), .rnd ({Fresh[10784], Fresh[10783], Fresh[10782], Fresh[10781], Fresh[10780], Fresh[10779], Fresh[10778], Fresh[10777], Fresh[10776], Fresh[10775], Fresh[10774], Fresh[10773], Fresh[10772], Fresh[10771], Fresh[10770]}), .outt ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, n2746}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2818 ( .ina ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, new_AGEMA_signal_3827, new_AGEMA_signal_3826, n2759}), .inb ({new_AGEMA_signal_21511, new_AGEMA_signal_21509, new_AGEMA_signal_21507, new_AGEMA_signal_21505, new_AGEMA_signal_21503}), .clk ( clk ), .rnd ({Fresh[10799], Fresh[10798], Fresh[10797], Fresh[10796], Fresh[10795], Fresh[10794], Fresh[10793], Fresh[10792], Fresh[10791], Fresh[10790], Fresh[10789], Fresh[10788], Fresh[10787], Fresh[10786], Fresh[10785]}), .outt ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, new_AGEMA_signal_4063, new_AGEMA_signal_4062, n2804}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2824 ( .ina ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, new_AGEMA_signal_3831, new_AGEMA_signal_3830, n2771}), .inb ({new_AGEMA_signal_21531, new_AGEMA_signal_21527, new_AGEMA_signal_21523, new_AGEMA_signal_21519, new_AGEMA_signal_21515}), .clk ( clk ), .rnd ({Fresh[10814], Fresh[10813], Fresh[10812], Fresh[10811], Fresh[10810], Fresh[10809], Fresh[10808], Fresh[10807], Fresh[10806], Fresh[10805], Fresh[10804], Fresh[10803], Fresh[10802], Fresh[10801], Fresh[10800]}), .outt ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, new_AGEMA_signal_4067, new_AGEMA_signal_4066, n2802}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2838 ( .ina ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, n2798}), .inb ({new_AGEMA_signal_21541, new_AGEMA_signal_21539, new_AGEMA_signal_21537, new_AGEMA_signal_21535, new_AGEMA_signal_21533}), .clk ( clk ), .rnd ({Fresh[10829], Fresh[10828], Fresh[10827], Fresh[10826], Fresh[10825], Fresh[10824], Fresh[10823], Fresh[10822], Fresh[10821], Fresh[10820], Fresh[10819], Fresh[10818], Fresh[10817], Fresh[10816], Fresh[10815]}), .outt ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, n2799}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2852 ( .ina ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, new_AGEMA_signal_3839, new_AGEMA_signal_3838, n2826}), .inb ({new_AGEMA_signal_21571, new_AGEMA_signal_21565, new_AGEMA_signal_21559, new_AGEMA_signal_21553, new_AGEMA_signal_21547}), .clk ( clk ), .rnd ({Fresh[10844], Fresh[10843], Fresh[10842], Fresh[10841], Fresh[10840], Fresh[10839], Fresh[10838], Fresh[10837], Fresh[10836], Fresh[10835], Fresh[10834], Fresh[10833], Fresh[10832], Fresh[10831], Fresh[10830]}), .outt ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, new_AGEMA_signal_4074, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C ( clk ), .D ( new_AGEMA_signal_21572 ), .Q ( new_AGEMA_signal_21573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C ( clk ), .D ( new_AGEMA_signal_21574 ), .Q ( new_AGEMA_signal_21575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C ( clk ), .D ( new_AGEMA_signal_21576 ), .Q ( new_AGEMA_signal_21577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C ( clk ), .D ( new_AGEMA_signal_21578 ), .Q ( new_AGEMA_signal_21579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C ( clk ), .D ( new_AGEMA_signal_21580 ), .Q ( new_AGEMA_signal_21581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C ( clk ), .D ( new_AGEMA_signal_21588 ), .Q ( new_AGEMA_signal_21589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C ( clk ), .D ( new_AGEMA_signal_21596 ), .Q ( new_AGEMA_signal_21597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C ( clk ), .D ( new_AGEMA_signal_21604 ), .Q ( new_AGEMA_signal_21605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C ( clk ), .D ( new_AGEMA_signal_21612 ), .Q ( new_AGEMA_signal_21613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C ( clk ), .D ( new_AGEMA_signal_21620 ), .Q ( new_AGEMA_signal_21621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C ( clk ), .D ( new_AGEMA_signal_21622 ), .Q ( new_AGEMA_signal_21623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C ( clk ), .D ( new_AGEMA_signal_21624 ), .Q ( new_AGEMA_signal_21625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C ( clk ), .D ( new_AGEMA_signal_21626 ), .Q ( new_AGEMA_signal_21627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C ( clk ), .D ( new_AGEMA_signal_21628 ), .Q ( new_AGEMA_signal_21629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C ( clk ), .D ( new_AGEMA_signal_21630 ), .Q ( new_AGEMA_signal_21631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C ( clk ), .D ( new_AGEMA_signal_21634 ), .Q ( new_AGEMA_signal_21635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C ( clk ), .D ( new_AGEMA_signal_21638 ), .Q ( new_AGEMA_signal_21639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C ( clk ), .D ( new_AGEMA_signal_21642 ), .Q ( new_AGEMA_signal_21643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C ( clk ), .D ( new_AGEMA_signal_21646 ), .Q ( new_AGEMA_signal_21647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C ( clk ), .D ( new_AGEMA_signal_21650 ), .Q ( new_AGEMA_signal_21651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C ( clk ), .D ( new_AGEMA_signal_21658 ), .Q ( new_AGEMA_signal_21659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C ( clk ), .D ( new_AGEMA_signal_21666 ), .Q ( new_AGEMA_signal_21667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C ( clk ), .D ( new_AGEMA_signal_21674 ), .Q ( new_AGEMA_signal_21675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C ( clk ), .D ( new_AGEMA_signal_21682 ), .Q ( new_AGEMA_signal_21683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C ( clk ), .D ( new_AGEMA_signal_21690 ), .Q ( new_AGEMA_signal_21691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C ( clk ), .D ( new_AGEMA_signal_21692 ), .Q ( new_AGEMA_signal_21693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C ( clk ), .D ( new_AGEMA_signal_21694 ), .Q ( new_AGEMA_signal_21695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C ( clk ), .D ( new_AGEMA_signal_21696 ), .Q ( new_AGEMA_signal_21697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C ( clk ), .D ( new_AGEMA_signal_21698 ), .Q ( new_AGEMA_signal_21699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C ( clk ), .D ( new_AGEMA_signal_21700 ), .Q ( new_AGEMA_signal_21701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C ( clk ), .D ( new_AGEMA_signal_21706 ), .Q ( new_AGEMA_signal_21707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C ( clk ), .D ( new_AGEMA_signal_21712 ), .Q ( new_AGEMA_signal_21713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C ( clk ), .D ( new_AGEMA_signal_21718 ), .Q ( new_AGEMA_signal_21719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C ( clk ), .D ( new_AGEMA_signal_21724 ), .Q ( new_AGEMA_signal_21725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C ( clk ), .D ( new_AGEMA_signal_21730 ), .Q ( new_AGEMA_signal_21731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C ( clk ), .D ( new_AGEMA_signal_21734 ), .Q ( new_AGEMA_signal_21735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C ( clk ), .D ( new_AGEMA_signal_21738 ), .Q ( new_AGEMA_signal_21739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C ( clk ), .D ( new_AGEMA_signal_21742 ), .Q ( new_AGEMA_signal_21743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C ( clk ), .D ( new_AGEMA_signal_21746 ), .Q ( new_AGEMA_signal_21747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C ( clk ), .D ( new_AGEMA_signal_21750 ), .Q ( new_AGEMA_signal_21751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C ( clk ), .D ( new_AGEMA_signal_21758 ), .Q ( new_AGEMA_signal_21759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C ( clk ), .D ( new_AGEMA_signal_21766 ), .Q ( new_AGEMA_signal_21767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C ( clk ), .D ( new_AGEMA_signal_21774 ), .Q ( new_AGEMA_signal_21775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C ( clk ), .D ( new_AGEMA_signal_21782 ), .Q ( new_AGEMA_signal_21783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C ( clk ), .D ( new_AGEMA_signal_21790 ), .Q ( new_AGEMA_signal_21791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C ( clk ), .D ( new_AGEMA_signal_21794 ), .Q ( new_AGEMA_signal_21795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C ( clk ), .D ( new_AGEMA_signal_21798 ), .Q ( new_AGEMA_signal_21799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C ( clk ), .D ( new_AGEMA_signal_21802 ), .Q ( new_AGEMA_signal_21803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C ( clk ), .D ( new_AGEMA_signal_21806 ), .Q ( new_AGEMA_signal_21807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C ( clk ), .D ( new_AGEMA_signal_21810 ), .Q ( new_AGEMA_signal_21811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C ( clk ), .D ( new_AGEMA_signal_21816 ), .Q ( new_AGEMA_signal_21817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C ( clk ), .D ( new_AGEMA_signal_21822 ), .Q ( new_AGEMA_signal_21823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C ( clk ), .D ( new_AGEMA_signal_21828 ), .Q ( new_AGEMA_signal_21829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C ( clk ), .D ( new_AGEMA_signal_21834 ), .Q ( new_AGEMA_signal_21835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C ( clk ), .D ( new_AGEMA_signal_21840 ), .Q ( new_AGEMA_signal_21841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C ( clk ), .D ( new_AGEMA_signal_21846 ), .Q ( new_AGEMA_signal_21847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C ( clk ), .D ( new_AGEMA_signal_21852 ), .Q ( new_AGEMA_signal_21853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C ( clk ), .D ( new_AGEMA_signal_21858 ), .Q ( new_AGEMA_signal_21859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C ( clk ), .D ( new_AGEMA_signal_21864 ), .Q ( new_AGEMA_signal_21865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C ( clk ), .D ( new_AGEMA_signal_21870 ), .Q ( new_AGEMA_signal_21871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C ( clk ), .D ( new_AGEMA_signal_21876 ), .Q ( new_AGEMA_signal_21877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C ( clk ), .D ( new_AGEMA_signal_21882 ), .Q ( new_AGEMA_signal_21883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C ( clk ), .D ( new_AGEMA_signal_21888 ), .Q ( new_AGEMA_signal_21889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C ( clk ), .D ( new_AGEMA_signal_21894 ), .Q ( new_AGEMA_signal_21895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C ( clk ), .D ( new_AGEMA_signal_21900 ), .Q ( new_AGEMA_signal_21901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C ( clk ), .D ( new_AGEMA_signal_21906 ), .Q ( new_AGEMA_signal_21907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C ( clk ), .D ( new_AGEMA_signal_21912 ), .Q ( new_AGEMA_signal_21913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C ( clk ), .D ( new_AGEMA_signal_21918 ), .Q ( new_AGEMA_signal_21919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C ( clk ), .D ( new_AGEMA_signal_21924 ), .Q ( new_AGEMA_signal_21925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C ( clk ), .D ( new_AGEMA_signal_21930 ), .Q ( new_AGEMA_signal_21931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C ( clk ), .D ( new_AGEMA_signal_21936 ), .Q ( new_AGEMA_signal_21937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C ( clk ), .D ( new_AGEMA_signal_21942 ), .Q ( new_AGEMA_signal_21943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C ( clk ), .D ( new_AGEMA_signal_21948 ), .Q ( new_AGEMA_signal_21949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C ( clk ), .D ( new_AGEMA_signal_21954 ), .Q ( new_AGEMA_signal_21955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C ( clk ), .D ( new_AGEMA_signal_21960 ), .Q ( new_AGEMA_signal_21961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C ( clk ), .D ( new_AGEMA_signal_21964 ), .Q ( new_AGEMA_signal_21965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C ( clk ), .D ( new_AGEMA_signal_21968 ), .Q ( new_AGEMA_signal_21969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C ( clk ), .D ( new_AGEMA_signal_21972 ), .Q ( new_AGEMA_signal_21973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C ( clk ), .D ( new_AGEMA_signal_21976 ), .Q ( new_AGEMA_signal_21977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C ( clk ), .D ( new_AGEMA_signal_21980 ), .Q ( new_AGEMA_signal_21981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C ( clk ), .D ( new_AGEMA_signal_21988 ), .Q ( new_AGEMA_signal_21989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C ( clk ), .D ( new_AGEMA_signal_21996 ), .Q ( new_AGEMA_signal_21997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C ( clk ), .D ( new_AGEMA_signal_22004 ), .Q ( new_AGEMA_signal_22005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C ( clk ), .D ( new_AGEMA_signal_22012 ), .Q ( new_AGEMA_signal_22013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C ( clk ), .D ( new_AGEMA_signal_22020 ), .Q ( new_AGEMA_signal_22021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C ( clk ), .D ( new_AGEMA_signal_22024 ), .Q ( new_AGEMA_signal_22025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C ( clk ), .D ( new_AGEMA_signal_22028 ), .Q ( new_AGEMA_signal_22029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C ( clk ), .D ( new_AGEMA_signal_22032 ), .Q ( new_AGEMA_signal_22033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C ( clk ), .D ( new_AGEMA_signal_22036 ), .Q ( new_AGEMA_signal_22037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C ( clk ), .D ( new_AGEMA_signal_22040 ), .Q ( new_AGEMA_signal_22041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C ( clk ), .D ( new_AGEMA_signal_22046 ), .Q ( new_AGEMA_signal_22047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C ( clk ), .D ( new_AGEMA_signal_22052 ), .Q ( new_AGEMA_signal_22053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C ( clk ), .D ( new_AGEMA_signal_22058 ), .Q ( new_AGEMA_signal_22059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C ( clk ), .D ( new_AGEMA_signal_22064 ), .Q ( new_AGEMA_signal_22065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C ( clk ), .D ( new_AGEMA_signal_22070 ), .Q ( new_AGEMA_signal_22071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C ( clk ), .D ( new_AGEMA_signal_22078 ), .Q ( new_AGEMA_signal_22079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C ( clk ), .D ( new_AGEMA_signal_22086 ), .Q ( new_AGEMA_signal_22087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C ( clk ), .D ( new_AGEMA_signal_22094 ), .Q ( new_AGEMA_signal_22095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C ( clk ), .D ( new_AGEMA_signal_22102 ), .Q ( new_AGEMA_signal_22103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C ( clk ), .D ( new_AGEMA_signal_22110 ), .Q ( new_AGEMA_signal_22111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C ( clk ), .D ( new_AGEMA_signal_22112 ), .Q ( new_AGEMA_signal_22113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C ( clk ), .D ( new_AGEMA_signal_22114 ), .Q ( new_AGEMA_signal_22115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C ( clk ), .D ( new_AGEMA_signal_22116 ), .Q ( new_AGEMA_signal_22117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C ( clk ), .D ( new_AGEMA_signal_22118 ), .Q ( new_AGEMA_signal_22119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C ( clk ), .D ( new_AGEMA_signal_22120 ), .Q ( new_AGEMA_signal_22121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C ( clk ), .D ( new_AGEMA_signal_22126 ), .Q ( new_AGEMA_signal_22127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C ( clk ), .D ( new_AGEMA_signal_22132 ), .Q ( new_AGEMA_signal_22133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C ( clk ), .D ( new_AGEMA_signal_22138 ), .Q ( new_AGEMA_signal_22139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C ( clk ), .D ( new_AGEMA_signal_22144 ), .Q ( new_AGEMA_signal_22145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C ( clk ), .D ( new_AGEMA_signal_22150 ), .Q ( new_AGEMA_signal_22151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C ( clk ), .D ( new_AGEMA_signal_22152 ), .Q ( new_AGEMA_signal_22153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C ( clk ), .D ( new_AGEMA_signal_22154 ), .Q ( new_AGEMA_signal_22155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C ( clk ), .D ( new_AGEMA_signal_22156 ), .Q ( new_AGEMA_signal_22157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C ( clk ), .D ( new_AGEMA_signal_22158 ), .Q ( new_AGEMA_signal_22159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C ( clk ), .D ( new_AGEMA_signal_22160 ), .Q ( new_AGEMA_signal_22161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C ( clk ), .D ( new_AGEMA_signal_22162 ), .Q ( new_AGEMA_signal_22163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C ( clk ), .D ( new_AGEMA_signal_22164 ), .Q ( new_AGEMA_signal_22165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C ( clk ), .D ( new_AGEMA_signal_22166 ), .Q ( new_AGEMA_signal_22167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C ( clk ), .D ( new_AGEMA_signal_22168 ), .Q ( new_AGEMA_signal_22169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C ( clk ), .D ( new_AGEMA_signal_22170 ), .Q ( new_AGEMA_signal_22171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C ( clk ), .D ( new_AGEMA_signal_22176 ), .Q ( new_AGEMA_signal_22177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C ( clk ), .D ( new_AGEMA_signal_22182 ), .Q ( new_AGEMA_signal_22183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C ( clk ), .D ( new_AGEMA_signal_22188 ), .Q ( new_AGEMA_signal_22189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C ( clk ), .D ( new_AGEMA_signal_22194 ), .Q ( new_AGEMA_signal_22195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C ( clk ), .D ( new_AGEMA_signal_22200 ), .Q ( new_AGEMA_signal_22201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C ( clk ), .D ( new_AGEMA_signal_22206 ), .Q ( new_AGEMA_signal_22207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C ( clk ), .D ( new_AGEMA_signal_22212 ), .Q ( new_AGEMA_signal_22213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C ( clk ), .D ( new_AGEMA_signal_22218 ), .Q ( new_AGEMA_signal_22219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C ( clk ), .D ( new_AGEMA_signal_22224 ), .Q ( new_AGEMA_signal_22225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C ( clk ), .D ( new_AGEMA_signal_22230 ), .Q ( new_AGEMA_signal_22231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C ( clk ), .D ( new_AGEMA_signal_22238 ), .Q ( new_AGEMA_signal_22239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C ( clk ), .D ( new_AGEMA_signal_22246 ), .Q ( new_AGEMA_signal_22247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C ( clk ), .D ( new_AGEMA_signal_22254 ), .Q ( new_AGEMA_signal_22255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C ( clk ), .D ( new_AGEMA_signal_22262 ), .Q ( new_AGEMA_signal_22263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C ( clk ), .D ( new_AGEMA_signal_22270 ), .Q ( new_AGEMA_signal_22271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C ( clk ), .D ( new_AGEMA_signal_22278 ), .Q ( new_AGEMA_signal_22279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C ( clk ), .D ( new_AGEMA_signal_22286 ), .Q ( new_AGEMA_signal_22287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C ( clk ), .D ( new_AGEMA_signal_22294 ), .Q ( new_AGEMA_signal_22295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C ( clk ), .D ( new_AGEMA_signal_22302 ), .Q ( new_AGEMA_signal_22303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C ( clk ), .D ( new_AGEMA_signal_22310 ), .Q ( new_AGEMA_signal_22311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C ( clk ), .D ( new_AGEMA_signal_22316 ), .Q ( new_AGEMA_signal_22317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C ( clk ), .D ( new_AGEMA_signal_22322 ), .Q ( new_AGEMA_signal_22323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C ( clk ), .D ( new_AGEMA_signal_22328 ), .Q ( new_AGEMA_signal_22329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C ( clk ), .D ( new_AGEMA_signal_22334 ), .Q ( new_AGEMA_signal_22335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C ( clk ), .D ( new_AGEMA_signal_22340 ), .Q ( new_AGEMA_signal_22341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C ( clk ), .D ( new_AGEMA_signal_22346 ), .Q ( new_AGEMA_signal_22347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C ( clk ), .D ( new_AGEMA_signal_22352 ), .Q ( new_AGEMA_signal_22353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C ( clk ), .D ( new_AGEMA_signal_22358 ), .Q ( new_AGEMA_signal_22359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C ( clk ), .D ( new_AGEMA_signal_22364 ), .Q ( new_AGEMA_signal_22365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C ( clk ), .D ( new_AGEMA_signal_22370 ), .Q ( new_AGEMA_signal_22371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C ( clk ), .D ( new_AGEMA_signal_22372 ), .Q ( new_AGEMA_signal_22373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C ( clk ), .D ( new_AGEMA_signal_22374 ), .Q ( new_AGEMA_signal_22375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C ( clk ), .D ( new_AGEMA_signal_22376 ), .Q ( new_AGEMA_signal_22377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C ( clk ), .D ( new_AGEMA_signal_22378 ), .Q ( new_AGEMA_signal_22379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C ( clk ), .D ( new_AGEMA_signal_22380 ), .Q ( new_AGEMA_signal_22381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C ( clk ), .D ( new_AGEMA_signal_22384 ), .Q ( new_AGEMA_signal_22385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C ( clk ), .D ( new_AGEMA_signal_22388 ), .Q ( new_AGEMA_signal_22389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C ( clk ), .D ( new_AGEMA_signal_22392 ), .Q ( new_AGEMA_signal_22393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C ( clk ), .D ( new_AGEMA_signal_22396 ), .Q ( new_AGEMA_signal_22397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C ( clk ), .D ( new_AGEMA_signal_22400 ), .Q ( new_AGEMA_signal_22401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C ( clk ), .D ( new_AGEMA_signal_22404 ), .Q ( new_AGEMA_signal_22405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C ( clk ), .D ( new_AGEMA_signal_22408 ), .Q ( new_AGEMA_signal_22409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C ( clk ), .D ( new_AGEMA_signal_22412 ), .Q ( new_AGEMA_signal_22413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C ( clk ), .D ( new_AGEMA_signal_22416 ), .Q ( new_AGEMA_signal_22417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C ( clk ), .D ( new_AGEMA_signal_22420 ), .Q ( new_AGEMA_signal_22421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C ( clk ), .D ( new_AGEMA_signal_22424 ), .Q ( new_AGEMA_signal_22425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C ( clk ), .D ( new_AGEMA_signal_22428 ), .Q ( new_AGEMA_signal_22429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C ( clk ), .D ( new_AGEMA_signal_22432 ), .Q ( new_AGEMA_signal_22433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C ( clk ), .D ( new_AGEMA_signal_22436 ), .Q ( new_AGEMA_signal_22437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C ( clk ), .D ( new_AGEMA_signal_22440 ), .Q ( new_AGEMA_signal_22441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C ( clk ), .D ( new_AGEMA_signal_22442 ), .Q ( new_AGEMA_signal_22443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C ( clk ), .D ( new_AGEMA_signal_22444 ), .Q ( new_AGEMA_signal_22445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C ( clk ), .D ( new_AGEMA_signal_22446 ), .Q ( new_AGEMA_signal_22447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C ( clk ), .D ( new_AGEMA_signal_22448 ), .Q ( new_AGEMA_signal_22449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C ( clk ), .D ( new_AGEMA_signal_22450 ), .Q ( new_AGEMA_signal_22451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C ( clk ), .D ( new_AGEMA_signal_22454 ), .Q ( new_AGEMA_signal_22455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C ( clk ), .D ( new_AGEMA_signal_22460 ), .Q ( new_AGEMA_signal_22461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C ( clk ), .D ( new_AGEMA_signal_22466 ), .Q ( new_AGEMA_signal_22467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C ( clk ), .D ( new_AGEMA_signal_22472 ), .Q ( new_AGEMA_signal_22473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C ( clk ), .D ( new_AGEMA_signal_22478 ), .Q ( new_AGEMA_signal_22479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C ( clk ), .D ( new_AGEMA_signal_22492 ), .Q ( new_AGEMA_signal_22493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C ( clk ), .D ( new_AGEMA_signal_22496 ), .Q ( new_AGEMA_signal_22497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C ( clk ), .D ( new_AGEMA_signal_22500 ), .Q ( new_AGEMA_signal_22501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C ( clk ), .D ( new_AGEMA_signal_22504 ), .Q ( new_AGEMA_signal_22505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C ( clk ), .D ( new_AGEMA_signal_22508 ), .Q ( new_AGEMA_signal_22509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C ( clk ), .D ( new_AGEMA_signal_22516 ), .Q ( new_AGEMA_signal_22517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C ( clk ), .D ( new_AGEMA_signal_22524 ), .Q ( new_AGEMA_signal_22525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C ( clk ), .D ( new_AGEMA_signal_22532 ), .Q ( new_AGEMA_signal_22533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C ( clk ), .D ( new_AGEMA_signal_22540 ), .Q ( new_AGEMA_signal_22541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C ( clk ), .D ( new_AGEMA_signal_22548 ), .Q ( new_AGEMA_signal_22549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C ( clk ), .D ( new_AGEMA_signal_22556 ), .Q ( new_AGEMA_signal_22557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C ( clk ), .D ( new_AGEMA_signal_22564 ), .Q ( new_AGEMA_signal_22565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C ( clk ), .D ( new_AGEMA_signal_22572 ), .Q ( new_AGEMA_signal_22573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C ( clk ), .D ( new_AGEMA_signal_22580 ), .Q ( new_AGEMA_signal_22581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C ( clk ), .D ( new_AGEMA_signal_22588 ), .Q ( new_AGEMA_signal_22589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C ( clk ), .D ( new_AGEMA_signal_22596 ), .Q ( new_AGEMA_signal_22597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C ( clk ), .D ( new_AGEMA_signal_22604 ), .Q ( new_AGEMA_signal_22605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C ( clk ), .D ( new_AGEMA_signal_22612 ), .Q ( new_AGEMA_signal_22613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C ( clk ), .D ( new_AGEMA_signal_22620 ), .Q ( new_AGEMA_signal_22621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C ( clk ), .D ( new_AGEMA_signal_22628 ), .Q ( new_AGEMA_signal_22629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C ( clk ), .D ( new_AGEMA_signal_22636 ), .Q ( new_AGEMA_signal_22637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C ( clk ), .D ( new_AGEMA_signal_22644 ), .Q ( new_AGEMA_signal_22645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C ( clk ), .D ( new_AGEMA_signal_22652 ), .Q ( new_AGEMA_signal_22653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C ( clk ), .D ( new_AGEMA_signal_22660 ), .Q ( new_AGEMA_signal_22661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C ( clk ), .D ( new_AGEMA_signal_22668 ), .Q ( new_AGEMA_signal_22669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C ( clk ), .D ( new_AGEMA_signal_22674 ), .Q ( new_AGEMA_signal_22675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C ( clk ), .D ( new_AGEMA_signal_22680 ), .Q ( new_AGEMA_signal_22681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C ( clk ), .D ( new_AGEMA_signal_22686 ), .Q ( new_AGEMA_signal_22687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C ( clk ), .D ( new_AGEMA_signal_22692 ), .Q ( new_AGEMA_signal_22693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C ( clk ), .D ( new_AGEMA_signal_22698 ), .Q ( new_AGEMA_signal_22699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C ( clk ), .D ( new_AGEMA_signal_22708 ), .Q ( new_AGEMA_signal_22709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C ( clk ), .D ( new_AGEMA_signal_22718 ), .Q ( new_AGEMA_signal_22719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C ( clk ), .D ( new_AGEMA_signal_22728 ), .Q ( new_AGEMA_signal_22729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C ( clk ), .D ( new_AGEMA_signal_22738 ), .Q ( new_AGEMA_signal_22739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C ( clk ), .D ( new_AGEMA_signal_22748 ), .Q ( new_AGEMA_signal_22749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C ( clk ), .D ( new_AGEMA_signal_22756 ), .Q ( new_AGEMA_signal_22757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C ( clk ), .D ( new_AGEMA_signal_22764 ), .Q ( new_AGEMA_signal_22765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C ( clk ), .D ( new_AGEMA_signal_22772 ), .Q ( new_AGEMA_signal_22773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C ( clk ), .D ( new_AGEMA_signal_22780 ), .Q ( new_AGEMA_signal_22781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C ( clk ), .D ( new_AGEMA_signal_22788 ), .Q ( new_AGEMA_signal_22789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C ( clk ), .D ( new_AGEMA_signal_22796 ), .Q ( new_AGEMA_signal_22797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C ( clk ), .D ( new_AGEMA_signal_22804 ), .Q ( new_AGEMA_signal_22805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C ( clk ), .D ( new_AGEMA_signal_22812 ), .Q ( new_AGEMA_signal_22813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C ( clk ), .D ( new_AGEMA_signal_22820 ), .Q ( new_AGEMA_signal_22821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C ( clk ), .D ( new_AGEMA_signal_22828 ), .Q ( new_AGEMA_signal_22829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C ( clk ), .D ( new_AGEMA_signal_22836 ), .Q ( new_AGEMA_signal_22837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C ( clk ), .D ( new_AGEMA_signal_22844 ), .Q ( new_AGEMA_signal_22845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C ( clk ), .D ( new_AGEMA_signal_22852 ), .Q ( new_AGEMA_signal_22853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C ( clk ), .D ( new_AGEMA_signal_22860 ), .Q ( new_AGEMA_signal_22861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C ( clk ), .D ( new_AGEMA_signal_22868 ), .Q ( new_AGEMA_signal_22869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C ( clk ), .D ( new_AGEMA_signal_22882 ), .Q ( new_AGEMA_signal_22883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C ( clk ), .D ( new_AGEMA_signal_22886 ), .Q ( new_AGEMA_signal_22887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C ( clk ), .D ( new_AGEMA_signal_22890 ), .Q ( new_AGEMA_signal_22891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C ( clk ), .D ( new_AGEMA_signal_22894 ), .Q ( new_AGEMA_signal_22895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C ( clk ), .D ( new_AGEMA_signal_22898 ), .Q ( new_AGEMA_signal_22899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C ( clk ), .D ( new_AGEMA_signal_22904 ), .Q ( new_AGEMA_signal_22905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C ( clk ), .D ( new_AGEMA_signal_22910 ), .Q ( new_AGEMA_signal_22911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C ( clk ), .D ( new_AGEMA_signal_22916 ), .Q ( new_AGEMA_signal_22917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C ( clk ), .D ( new_AGEMA_signal_22922 ), .Q ( new_AGEMA_signal_22923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C ( clk ), .D ( new_AGEMA_signal_22928 ), .Q ( new_AGEMA_signal_22929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C ( clk ), .D ( new_AGEMA_signal_22932 ), .Q ( new_AGEMA_signal_22933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C ( clk ), .D ( new_AGEMA_signal_22936 ), .Q ( new_AGEMA_signal_22937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C ( clk ), .D ( new_AGEMA_signal_22940 ), .Q ( new_AGEMA_signal_22941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C ( clk ), .D ( new_AGEMA_signal_22944 ), .Q ( new_AGEMA_signal_22945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C ( clk ), .D ( new_AGEMA_signal_22948 ), .Q ( new_AGEMA_signal_22949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C ( clk ), .D ( new_AGEMA_signal_22958 ), .Q ( new_AGEMA_signal_22959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C ( clk ), .D ( new_AGEMA_signal_22968 ), .Q ( new_AGEMA_signal_22969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C ( clk ), .D ( new_AGEMA_signal_22978 ), .Q ( new_AGEMA_signal_22979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C ( clk ), .D ( new_AGEMA_signal_22988 ), .Q ( new_AGEMA_signal_22989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C ( clk ), .D ( new_AGEMA_signal_22998 ), .Q ( new_AGEMA_signal_22999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C ( clk ), .D ( new_AGEMA_signal_23006 ), .Q ( new_AGEMA_signal_23007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C ( clk ), .D ( new_AGEMA_signal_23014 ), .Q ( new_AGEMA_signal_23015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C ( clk ), .D ( new_AGEMA_signal_23022 ), .Q ( new_AGEMA_signal_23023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C ( clk ), .D ( new_AGEMA_signal_23030 ), .Q ( new_AGEMA_signal_23031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C ( clk ), .D ( new_AGEMA_signal_23038 ), .Q ( new_AGEMA_signal_23039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C ( clk ), .D ( new_AGEMA_signal_23042 ), .Q ( new_AGEMA_signal_23043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C ( clk ), .D ( new_AGEMA_signal_23046 ), .Q ( new_AGEMA_signal_23047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C ( clk ), .D ( new_AGEMA_signal_23050 ), .Q ( new_AGEMA_signal_23051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C ( clk ), .D ( new_AGEMA_signal_23054 ), .Q ( new_AGEMA_signal_23055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C ( clk ), .D ( new_AGEMA_signal_23058 ), .Q ( new_AGEMA_signal_23059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C ( clk ), .D ( new_AGEMA_signal_23076 ), .Q ( new_AGEMA_signal_23077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C ( clk ), .D ( new_AGEMA_signal_23084 ), .Q ( new_AGEMA_signal_23085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C ( clk ), .D ( new_AGEMA_signal_23092 ), .Q ( new_AGEMA_signal_23093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C ( clk ), .D ( new_AGEMA_signal_23100 ), .Q ( new_AGEMA_signal_23101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C ( clk ), .D ( new_AGEMA_signal_23108 ), .Q ( new_AGEMA_signal_23109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C ( clk ), .D ( new_AGEMA_signal_23116 ), .Q ( new_AGEMA_signal_23117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C ( clk ), .D ( new_AGEMA_signal_23124 ), .Q ( new_AGEMA_signal_23125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C ( clk ), .D ( new_AGEMA_signal_23132 ), .Q ( new_AGEMA_signal_23133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C ( clk ), .D ( new_AGEMA_signal_23140 ), .Q ( new_AGEMA_signal_23141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C ( clk ), .D ( new_AGEMA_signal_23148 ), .Q ( new_AGEMA_signal_23149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C ( clk ), .D ( new_AGEMA_signal_23154 ), .Q ( new_AGEMA_signal_23155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C ( clk ), .D ( new_AGEMA_signal_23160 ), .Q ( new_AGEMA_signal_23161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C ( clk ), .D ( new_AGEMA_signal_23166 ), .Q ( new_AGEMA_signal_23167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C ( clk ), .D ( new_AGEMA_signal_23172 ), .Q ( new_AGEMA_signal_23173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C ( clk ), .D ( new_AGEMA_signal_23178 ), .Q ( new_AGEMA_signal_23179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C ( clk ), .D ( new_AGEMA_signal_23182 ), .Q ( new_AGEMA_signal_23183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C ( clk ), .D ( new_AGEMA_signal_23186 ), .Q ( new_AGEMA_signal_23187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C ( clk ), .D ( new_AGEMA_signal_23190 ), .Q ( new_AGEMA_signal_23191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C ( clk ), .D ( new_AGEMA_signal_23194 ), .Q ( new_AGEMA_signal_23195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C ( clk ), .D ( new_AGEMA_signal_23198 ), .Q ( new_AGEMA_signal_23199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C ( clk ), .D ( new_AGEMA_signal_23206 ), .Q ( new_AGEMA_signal_23207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C ( clk ), .D ( new_AGEMA_signal_23214 ), .Q ( new_AGEMA_signal_23215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C ( clk ), .D ( new_AGEMA_signal_23222 ), .Q ( new_AGEMA_signal_23223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C ( clk ), .D ( new_AGEMA_signal_23230 ), .Q ( new_AGEMA_signal_23231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C ( clk ), .D ( new_AGEMA_signal_23238 ), .Q ( new_AGEMA_signal_23239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C ( clk ), .D ( new_AGEMA_signal_23252 ), .Q ( new_AGEMA_signal_23253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C ( clk ), .D ( new_AGEMA_signal_23258 ), .Q ( new_AGEMA_signal_23259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C ( clk ), .D ( new_AGEMA_signal_23264 ), .Q ( new_AGEMA_signal_23265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C ( clk ), .D ( new_AGEMA_signal_23270 ), .Q ( new_AGEMA_signal_23271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C ( clk ), .D ( new_AGEMA_signal_23276 ), .Q ( new_AGEMA_signal_23277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C ( clk ), .D ( new_AGEMA_signal_23282 ), .Q ( new_AGEMA_signal_23283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C ( clk ), .D ( new_AGEMA_signal_23288 ), .Q ( new_AGEMA_signal_23289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C ( clk ), .D ( new_AGEMA_signal_23294 ), .Q ( new_AGEMA_signal_23295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C ( clk ), .D ( new_AGEMA_signal_23300 ), .Q ( new_AGEMA_signal_23301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C ( clk ), .D ( new_AGEMA_signal_23306 ), .Q ( new_AGEMA_signal_23307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C ( clk ), .D ( new_AGEMA_signal_23312 ), .Q ( new_AGEMA_signal_23313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C ( clk ), .D ( new_AGEMA_signal_23318 ), .Q ( new_AGEMA_signal_23319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C ( clk ), .D ( new_AGEMA_signal_23324 ), .Q ( new_AGEMA_signal_23325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C ( clk ), .D ( new_AGEMA_signal_23330 ), .Q ( new_AGEMA_signal_23331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C ( clk ), .D ( new_AGEMA_signal_23336 ), .Q ( new_AGEMA_signal_23337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C ( clk ), .D ( new_AGEMA_signal_23364 ), .Q ( new_AGEMA_signal_23365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C ( clk ), .D ( new_AGEMA_signal_23372 ), .Q ( new_AGEMA_signal_23373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C ( clk ), .D ( new_AGEMA_signal_23380 ), .Q ( new_AGEMA_signal_23381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C ( clk ), .D ( new_AGEMA_signal_23388 ), .Q ( new_AGEMA_signal_23389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C ( clk ), .D ( new_AGEMA_signal_23396 ), .Q ( new_AGEMA_signal_23397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C ( clk ), .D ( new_AGEMA_signal_23402 ), .Q ( new_AGEMA_signal_23403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C ( clk ), .D ( new_AGEMA_signal_23408 ), .Q ( new_AGEMA_signal_23409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C ( clk ), .D ( new_AGEMA_signal_23414 ), .Q ( new_AGEMA_signal_23415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C ( clk ), .D ( new_AGEMA_signal_23420 ), .Q ( new_AGEMA_signal_23421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C ( clk ), .D ( new_AGEMA_signal_23426 ), .Q ( new_AGEMA_signal_23427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C ( clk ), .D ( new_AGEMA_signal_23454 ), .Q ( new_AGEMA_signal_23455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C ( clk ), .D ( new_AGEMA_signal_23462 ), .Q ( new_AGEMA_signal_23463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C ( clk ), .D ( new_AGEMA_signal_23470 ), .Q ( new_AGEMA_signal_23471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C ( clk ), .D ( new_AGEMA_signal_23478 ), .Q ( new_AGEMA_signal_23479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C ( clk ), .D ( new_AGEMA_signal_23486 ), .Q ( new_AGEMA_signal_23487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C ( clk ), .D ( new_AGEMA_signal_23494 ), .Q ( new_AGEMA_signal_23495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C ( clk ), .D ( new_AGEMA_signal_23502 ), .Q ( new_AGEMA_signal_23503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C ( clk ), .D ( new_AGEMA_signal_23510 ), .Q ( new_AGEMA_signal_23511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C ( clk ), .D ( new_AGEMA_signal_23518 ), .Q ( new_AGEMA_signal_23519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C ( clk ), .D ( new_AGEMA_signal_23526 ), .Q ( new_AGEMA_signal_23527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C ( clk ), .D ( new_AGEMA_signal_23536 ), .Q ( new_AGEMA_signal_23537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C ( clk ), .D ( new_AGEMA_signal_23546 ), .Q ( new_AGEMA_signal_23547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C ( clk ), .D ( new_AGEMA_signal_23556 ), .Q ( new_AGEMA_signal_23557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C ( clk ), .D ( new_AGEMA_signal_23566 ), .Q ( new_AGEMA_signal_23567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C ( clk ), .D ( new_AGEMA_signal_23576 ), .Q ( new_AGEMA_signal_23577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C ( clk ), .D ( new_AGEMA_signal_23584 ), .Q ( new_AGEMA_signal_23585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C ( clk ), .D ( new_AGEMA_signal_23592 ), .Q ( new_AGEMA_signal_23593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C ( clk ), .D ( new_AGEMA_signal_23600 ), .Q ( new_AGEMA_signal_23601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C ( clk ), .D ( new_AGEMA_signal_23608 ), .Q ( new_AGEMA_signal_23609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C ( clk ), .D ( new_AGEMA_signal_23616 ), .Q ( new_AGEMA_signal_23617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C ( clk ), .D ( new_AGEMA_signal_23622 ), .Q ( new_AGEMA_signal_23623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C ( clk ), .D ( new_AGEMA_signal_23628 ), .Q ( new_AGEMA_signal_23629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C ( clk ), .D ( new_AGEMA_signal_23634 ), .Q ( new_AGEMA_signal_23635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C ( clk ), .D ( new_AGEMA_signal_23640 ), .Q ( new_AGEMA_signal_23641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C ( clk ), .D ( new_AGEMA_signal_23646 ), .Q ( new_AGEMA_signal_23647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C ( clk ), .D ( new_AGEMA_signal_23672 ), .Q ( new_AGEMA_signal_23673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C ( clk ), .D ( new_AGEMA_signal_23678 ), .Q ( new_AGEMA_signal_23679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C ( clk ), .D ( new_AGEMA_signal_23684 ), .Q ( new_AGEMA_signal_23685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C ( clk ), .D ( new_AGEMA_signal_23690 ), .Q ( new_AGEMA_signal_23691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C ( clk ), .D ( new_AGEMA_signal_23696 ), .Q ( new_AGEMA_signal_23697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C ( clk ), .D ( new_AGEMA_signal_23704 ), .Q ( new_AGEMA_signal_23705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C ( clk ), .D ( new_AGEMA_signal_23712 ), .Q ( new_AGEMA_signal_23713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C ( clk ), .D ( new_AGEMA_signal_23720 ), .Q ( new_AGEMA_signal_23721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C ( clk ), .D ( new_AGEMA_signal_23728 ), .Q ( new_AGEMA_signal_23729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C ( clk ), .D ( new_AGEMA_signal_23736 ), .Q ( new_AGEMA_signal_23737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C ( clk ), .D ( new_AGEMA_signal_23742 ), .Q ( new_AGEMA_signal_23743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C ( clk ), .D ( new_AGEMA_signal_23748 ), .Q ( new_AGEMA_signal_23749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C ( clk ), .D ( new_AGEMA_signal_23754 ), .Q ( new_AGEMA_signal_23755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C ( clk ), .D ( new_AGEMA_signal_23760 ), .Q ( new_AGEMA_signal_23761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C ( clk ), .D ( new_AGEMA_signal_23766 ), .Q ( new_AGEMA_signal_23767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C ( clk ), .D ( new_AGEMA_signal_23784 ), .Q ( new_AGEMA_signal_23785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C ( clk ), .D ( new_AGEMA_signal_23792 ), .Q ( new_AGEMA_signal_23793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C ( clk ), .D ( new_AGEMA_signal_23800 ), .Q ( new_AGEMA_signal_23801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C ( clk ), .D ( new_AGEMA_signal_23808 ), .Q ( new_AGEMA_signal_23809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C ( clk ), .D ( new_AGEMA_signal_23816 ), .Q ( new_AGEMA_signal_23817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C ( clk ), .D ( new_AGEMA_signal_23842 ), .Q ( new_AGEMA_signal_23843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C ( clk ), .D ( new_AGEMA_signal_23848 ), .Q ( new_AGEMA_signal_23849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C ( clk ), .D ( new_AGEMA_signal_23854 ), .Q ( new_AGEMA_signal_23855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C ( clk ), .D ( new_AGEMA_signal_23860 ), .Q ( new_AGEMA_signal_23861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C ( clk ), .D ( new_AGEMA_signal_23866 ), .Q ( new_AGEMA_signal_23867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C ( clk ), .D ( new_AGEMA_signal_23872 ), .Q ( new_AGEMA_signal_23873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C ( clk ), .D ( new_AGEMA_signal_23878 ), .Q ( new_AGEMA_signal_23879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C ( clk ), .D ( new_AGEMA_signal_23884 ), .Q ( new_AGEMA_signal_23885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C ( clk ), .D ( new_AGEMA_signal_23890 ), .Q ( new_AGEMA_signal_23891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C ( clk ), .D ( new_AGEMA_signal_23896 ), .Q ( new_AGEMA_signal_23897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C ( clk ), .D ( new_AGEMA_signal_24004 ), .Q ( new_AGEMA_signal_24005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C ( clk ), .D ( new_AGEMA_signal_24014 ), .Q ( new_AGEMA_signal_24015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C ( clk ), .D ( new_AGEMA_signal_24024 ), .Q ( new_AGEMA_signal_24025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C ( clk ), .D ( new_AGEMA_signal_24034 ), .Q ( new_AGEMA_signal_24035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C ( clk ), .D ( new_AGEMA_signal_24044 ), .Q ( new_AGEMA_signal_24045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C ( clk ), .D ( new_AGEMA_signal_24152 ), .Q ( new_AGEMA_signal_24153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C ( clk ), .D ( new_AGEMA_signal_24160 ), .Q ( new_AGEMA_signal_24161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C ( clk ), .D ( new_AGEMA_signal_24168 ), .Q ( new_AGEMA_signal_24169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C ( clk ), .D ( new_AGEMA_signal_24176 ), .Q ( new_AGEMA_signal_24177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C ( clk ), .D ( new_AGEMA_signal_24184 ), .Q ( new_AGEMA_signal_24185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C ( clk ), .D ( new_AGEMA_signal_24222 ), .Q ( new_AGEMA_signal_24223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C ( clk ), .D ( new_AGEMA_signal_24230 ), .Q ( new_AGEMA_signal_24231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C ( clk ), .D ( new_AGEMA_signal_24238 ), .Q ( new_AGEMA_signal_24239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C ( clk ), .D ( new_AGEMA_signal_24246 ), .Q ( new_AGEMA_signal_24247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C ( clk ), .D ( new_AGEMA_signal_24254 ), .Q ( new_AGEMA_signal_24255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C ( clk ), .D ( new_AGEMA_signal_24262 ), .Q ( new_AGEMA_signal_24263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C ( clk ), .D ( new_AGEMA_signal_24270 ), .Q ( new_AGEMA_signal_24271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C ( clk ), .D ( new_AGEMA_signal_24278 ), .Q ( new_AGEMA_signal_24279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C ( clk ), .D ( new_AGEMA_signal_24286 ), .Q ( new_AGEMA_signal_24287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C ( clk ), .D ( new_AGEMA_signal_24294 ), .Q ( new_AGEMA_signal_24295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C ( clk ), .D ( new_AGEMA_signal_24352 ), .Q ( new_AGEMA_signal_24353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C ( clk ), .D ( new_AGEMA_signal_24360 ), .Q ( new_AGEMA_signal_24361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C ( clk ), .D ( new_AGEMA_signal_24368 ), .Q ( new_AGEMA_signal_24369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C ( clk ), .D ( new_AGEMA_signal_24376 ), .Q ( new_AGEMA_signal_24377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C ( clk ), .D ( new_AGEMA_signal_24384 ), .Q ( new_AGEMA_signal_24385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7680 ( .C ( clk ), .D ( new_AGEMA_signal_24454 ), .Q ( new_AGEMA_signal_24455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7692 ( .C ( clk ), .D ( new_AGEMA_signal_24466 ), .Q ( new_AGEMA_signal_24467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7704 ( .C ( clk ), .D ( new_AGEMA_signal_24478 ), .Q ( new_AGEMA_signal_24479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7716 ( .C ( clk ), .D ( new_AGEMA_signal_24490 ), .Q ( new_AGEMA_signal_24491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7728 ( .C ( clk ), .D ( new_AGEMA_signal_24502 ), .Q ( new_AGEMA_signal_24503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7742 ( .C ( clk ), .D ( new_AGEMA_signal_24516 ), .Q ( new_AGEMA_signal_24517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7756 ( .C ( clk ), .D ( new_AGEMA_signal_24530 ), .Q ( new_AGEMA_signal_24531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7770 ( .C ( clk ), .D ( new_AGEMA_signal_24544 ), .Q ( new_AGEMA_signal_24545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7784 ( .C ( clk ), .D ( new_AGEMA_signal_24558 ), .Q ( new_AGEMA_signal_24559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7798 ( .C ( clk ), .D ( new_AGEMA_signal_24572 ), .Q ( new_AGEMA_signal_24573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7852 ( .C ( clk ), .D ( new_AGEMA_signal_24626 ), .Q ( new_AGEMA_signal_24627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7866 ( .C ( clk ), .D ( new_AGEMA_signal_24640 ), .Q ( new_AGEMA_signal_24641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7880 ( .C ( clk ), .D ( new_AGEMA_signal_24654 ), .Q ( new_AGEMA_signal_24655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7894 ( .C ( clk ), .D ( new_AGEMA_signal_24668 ), .Q ( new_AGEMA_signal_24669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7908 ( .C ( clk ), .D ( new_AGEMA_signal_24682 ), .Q ( new_AGEMA_signal_24683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8032 ( .C ( clk ), .D ( new_AGEMA_signal_24806 ), .Q ( new_AGEMA_signal_24807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8048 ( .C ( clk ), .D ( new_AGEMA_signal_24822 ), .Q ( new_AGEMA_signal_24823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8064 ( .C ( clk ), .D ( new_AGEMA_signal_24838 ), .Q ( new_AGEMA_signal_24839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8080 ( .C ( clk ), .D ( new_AGEMA_signal_24854 ), .Q ( new_AGEMA_signal_24855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8096 ( .C ( clk ), .D ( new_AGEMA_signal_24870 ), .Q ( new_AGEMA_signal_24871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8142 ( .C ( clk ), .D ( new_AGEMA_signal_24916 ), .Q ( new_AGEMA_signal_24917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8158 ( .C ( clk ), .D ( new_AGEMA_signal_24932 ), .Q ( new_AGEMA_signal_24933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8174 ( .C ( clk ), .D ( new_AGEMA_signal_24948 ), .Q ( new_AGEMA_signal_24949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8190 ( .C ( clk ), .D ( new_AGEMA_signal_24964 ), .Q ( new_AGEMA_signal_24965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8206 ( .C ( clk ), .D ( new_AGEMA_signal_24980 ), .Q ( new_AGEMA_signal_24981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8390 ( .C ( clk ), .D ( new_AGEMA_signal_25164 ), .Q ( new_AGEMA_signal_25165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8406 ( .C ( clk ), .D ( new_AGEMA_signal_25180 ), .Q ( new_AGEMA_signal_25181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8422 ( .C ( clk ), .D ( new_AGEMA_signal_25196 ), .Q ( new_AGEMA_signal_25197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8438 ( .C ( clk ), .D ( new_AGEMA_signal_25212 ), .Q ( new_AGEMA_signal_25213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8454 ( .C ( clk ), .D ( new_AGEMA_signal_25228 ), .Q ( new_AGEMA_signal_25229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8522 ( .C ( clk ), .D ( new_AGEMA_signal_25296 ), .Q ( new_AGEMA_signal_25297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8540 ( .C ( clk ), .D ( new_AGEMA_signal_25314 ), .Q ( new_AGEMA_signal_25315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8558 ( .C ( clk ), .D ( new_AGEMA_signal_25332 ), .Q ( new_AGEMA_signal_25333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8576 ( .C ( clk ), .D ( new_AGEMA_signal_25350 ), .Q ( new_AGEMA_signal_25351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8594 ( .C ( clk ), .D ( new_AGEMA_signal_25368 ), .Q ( new_AGEMA_signal_25369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8772 ( .C ( clk ), .D ( new_AGEMA_signal_25546 ), .Q ( new_AGEMA_signal_25547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8792 ( .C ( clk ), .D ( new_AGEMA_signal_25566 ), .Q ( new_AGEMA_signal_25567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8812 ( .C ( clk ), .D ( new_AGEMA_signal_25586 ), .Q ( new_AGEMA_signal_25587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8832 ( .C ( clk ), .D ( new_AGEMA_signal_25606 ), .Q ( new_AGEMA_signal_25607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8852 ( .C ( clk ), .D ( new_AGEMA_signal_25626 ), .Q ( new_AGEMA_signal_25627 ) ) ;

    /* cells in depth 13 */
    buf_clk new_AGEMA_reg_buffer_5681 ( .C ( clk ), .D ( new_AGEMA_signal_22455 ), .Q ( new_AGEMA_signal_22456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C ( clk ), .D ( new_AGEMA_signal_22461 ), .Q ( new_AGEMA_signal_22462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C ( clk ), .D ( new_AGEMA_signal_22467 ), .Q ( new_AGEMA_signal_22468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C ( clk ), .D ( new_AGEMA_signal_22473 ), .Q ( new_AGEMA_signal_22474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C ( clk ), .D ( new_AGEMA_signal_22479 ), .Q ( new_AGEMA_signal_22480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C ( clk ), .D ( new_AGEMA_signal_22385 ), .Q ( new_AGEMA_signal_22482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C ( clk ), .D ( new_AGEMA_signal_22389 ), .Q ( new_AGEMA_signal_22484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C ( clk ), .D ( new_AGEMA_signal_22393 ), .Q ( new_AGEMA_signal_22486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C ( clk ), .D ( new_AGEMA_signal_22397 ), .Q ( new_AGEMA_signal_22488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C ( clk ), .D ( new_AGEMA_signal_22401 ), .Q ( new_AGEMA_signal_22490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C ( clk ), .D ( new_AGEMA_signal_22493 ), .Q ( new_AGEMA_signal_22494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C ( clk ), .D ( new_AGEMA_signal_22497 ), .Q ( new_AGEMA_signal_22498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C ( clk ), .D ( new_AGEMA_signal_22501 ), .Q ( new_AGEMA_signal_22502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C ( clk ), .D ( new_AGEMA_signal_22505 ), .Q ( new_AGEMA_signal_22506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C ( clk ), .D ( new_AGEMA_signal_22509 ), .Q ( new_AGEMA_signal_22510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C ( clk ), .D ( new_AGEMA_signal_22517 ), .Q ( new_AGEMA_signal_22518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C ( clk ), .D ( new_AGEMA_signal_22525 ), .Q ( new_AGEMA_signal_22526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C ( clk ), .D ( new_AGEMA_signal_22533 ), .Q ( new_AGEMA_signal_22534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C ( clk ), .D ( new_AGEMA_signal_22541 ), .Q ( new_AGEMA_signal_22542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C ( clk ), .D ( new_AGEMA_signal_22549 ), .Q ( new_AGEMA_signal_22550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C ( clk ), .D ( new_AGEMA_signal_22557 ), .Q ( new_AGEMA_signal_22558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C ( clk ), .D ( new_AGEMA_signal_22565 ), .Q ( new_AGEMA_signal_22566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C ( clk ), .D ( new_AGEMA_signal_22573 ), .Q ( new_AGEMA_signal_22574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C ( clk ), .D ( new_AGEMA_signal_22581 ), .Q ( new_AGEMA_signal_22582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C ( clk ), .D ( new_AGEMA_signal_22589 ), .Q ( new_AGEMA_signal_22590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C ( clk ), .D ( new_AGEMA_signal_22597 ), .Q ( new_AGEMA_signal_22598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C ( clk ), .D ( new_AGEMA_signal_22605 ), .Q ( new_AGEMA_signal_22606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C ( clk ), .D ( new_AGEMA_signal_22613 ), .Q ( new_AGEMA_signal_22614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C ( clk ), .D ( new_AGEMA_signal_22621 ), .Q ( new_AGEMA_signal_22622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C ( clk ), .D ( new_AGEMA_signal_22629 ), .Q ( new_AGEMA_signal_22630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C ( clk ), .D ( new_AGEMA_signal_22637 ), .Q ( new_AGEMA_signal_22638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C ( clk ), .D ( new_AGEMA_signal_22645 ), .Q ( new_AGEMA_signal_22646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C ( clk ), .D ( new_AGEMA_signal_22653 ), .Q ( new_AGEMA_signal_22654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C ( clk ), .D ( new_AGEMA_signal_22661 ), .Q ( new_AGEMA_signal_22662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C ( clk ), .D ( new_AGEMA_signal_22669 ), .Q ( new_AGEMA_signal_22670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C ( clk ), .D ( new_AGEMA_signal_22675 ), .Q ( new_AGEMA_signal_22676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C ( clk ), .D ( new_AGEMA_signal_22681 ), .Q ( new_AGEMA_signal_22682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C ( clk ), .D ( new_AGEMA_signal_22687 ), .Q ( new_AGEMA_signal_22688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C ( clk ), .D ( new_AGEMA_signal_22693 ), .Q ( new_AGEMA_signal_22694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C ( clk ), .D ( new_AGEMA_signal_22699 ), .Q ( new_AGEMA_signal_22700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C ( clk ), .D ( new_AGEMA_signal_22709 ), .Q ( new_AGEMA_signal_22710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C ( clk ), .D ( new_AGEMA_signal_22719 ), .Q ( new_AGEMA_signal_22720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C ( clk ), .D ( new_AGEMA_signal_22729 ), .Q ( new_AGEMA_signal_22730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C ( clk ), .D ( new_AGEMA_signal_22739 ), .Q ( new_AGEMA_signal_22740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C ( clk ), .D ( new_AGEMA_signal_22749 ), .Q ( new_AGEMA_signal_22750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C ( clk ), .D ( new_AGEMA_signal_22757 ), .Q ( new_AGEMA_signal_22758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C ( clk ), .D ( new_AGEMA_signal_22765 ), .Q ( new_AGEMA_signal_22766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C ( clk ), .D ( new_AGEMA_signal_22773 ), .Q ( new_AGEMA_signal_22774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C ( clk ), .D ( new_AGEMA_signal_22781 ), .Q ( new_AGEMA_signal_22782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C ( clk ), .D ( new_AGEMA_signal_22789 ), .Q ( new_AGEMA_signal_22790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C ( clk ), .D ( new_AGEMA_signal_22797 ), .Q ( new_AGEMA_signal_22798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C ( clk ), .D ( new_AGEMA_signal_22805 ), .Q ( new_AGEMA_signal_22806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C ( clk ), .D ( new_AGEMA_signal_22813 ), .Q ( new_AGEMA_signal_22814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C ( clk ), .D ( new_AGEMA_signal_22821 ), .Q ( new_AGEMA_signal_22822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C ( clk ), .D ( new_AGEMA_signal_22829 ), .Q ( new_AGEMA_signal_22830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C ( clk ), .D ( new_AGEMA_signal_22837 ), .Q ( new_AGEMA_signal_22838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C ( clk ), .D ( new_AGEMA_signal_22845 ), .Q ( new_AGEMA_signal_22846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C ( clk ), .D ( new_AGEMA_signal_22853 ), .Q ( new_AGEMA_signal_22854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C ( clk ), .D ( new_AGEMA_signal_22861 ), .Q ( new_AGEMA_signal_22862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C ( clk ), .D ( new_AGEMA_signal_22869 ), .Q ( new_AGEMA_signal_22870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C ( clk ), .D ( new_AGEMA_signal_21693 ), .Q ( new_AGEMA_signal_22872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C ( clk ), .D ( new_AGEMA_signal_21695 ), .Q ( new_AGEMA_signal_22874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C ( clk ), .D ( new_AGEMA_signal_21697 ), .Q ( new_AGEMA_signal_22876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C ( clk ), .D ( new_AGEMA_signal_21699 ), .Q ( new_AGEMA_signal_22878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C ( clk ), .D ( new_AGEMA_signal_21701 ), .Q ( new_AGEMA_signal_22880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C ( clk ), .D ( new_AGEMA_signal_22883 ), .Q ( new_AGEMA_signal_22884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C ( clk ), .D ( new_AGEMA_signal_22887 ), .Q ( new_AGEMA_signal_22888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C ( clk ), .D ( new_AGEMA_signal_22891 ), .Q ( new_AGEMA_signal_22892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C ( clk ), .D ( new_AGEMA_signal_22895 ), .Q ( new_AGEMA_signal_22896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C ( clk ), .D ( new_AGEMA_signal_22899 ), .Q ( new_AGEMA_signal_22900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C ( clk ), .D ( new_AGEMA_signal_22905 ), .Q ( new_AGEMA_signal_22906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C ( clk ), .D ( new_AGEMA_signal_22911 ), .Q ( new_AGEMA_signal_22912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C ( clk ), .D ( new_AGEMA_signal_22917 ), .Q ( new_AGEMA_signal_22918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C ( clk ), .D ( new_AGEMA_signal_22923 ), .Q ( new_AGEMA_signal_22924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C ( clk ), .D ( new_AGEMA_signal_22929 ), .Q ( new_AGEMA_signal_22930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C ( clk ), .D ( new_AGEMA_signal_22933 ), .Q ( new_AGEMA_signal_22934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C ( clk ), .D ( new_AGEMA_signal_22937 ), .Q ( new_AGEMA_signal_22938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C ( clk ), .D ( new_AGEMA_signal_22941 ), .Q ( new_AGEMA_signal_22942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C ( clk ), .D ( new_AGEMA_signal_22945 ), .Q ( new_AGEMA_signal_22946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C ( clk ), .D ( new_AGEMA_signal_22949 ), .Q ( new_AGEMA_signal_22950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C ( clk ), .D ( new_AGEMA_signal_22959 ), .Q ( new_AGEMA_signal_22960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C ( clk ), .D ( new_AGEMA_signal_22969 ), .Q ( new_AGEMA_signal_22970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C ( clk ), .D ( new_AGEMA_signal_22979 ), .Q ( new_AGEMA_signal_22980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C ( clk ), .D ( new_AGEMA_signal_22989 ), .Q ( new_AGEMA_signal_22990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C ( clk ), .D ( new_AGEMA_signal_22999 ), .Q ( new_AGEMA_signal_23000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C ( clk ), .D ( new_AGEMA_signal_23007 ), .Q ( new_AGEMA_signal_23008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C ( clk ), .D ( new_AGEMA_signal_23015 ), .Q ( new_AGEMA_signal_23016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C ( clk ), .D ( new_AGEMA_signal_23023 ), .Q ( new_AGEMA_signal_23024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C ( clk ), .D ( new_AGEMA_signal_23031 ), .Q ( new_AGEMA_signal_23032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C ( clk ), .D ( new_AGEMA_signal_23039 ), .Q ( new_AGEMA_signal_23040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C ( clk ), .D ( new_AGEMA_signal_23043 ), .Q ( new_AGEMA_signal_23044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C ( clk ), .D ( new_AGEMA_signal_23047 ), .Q ( new_AGEMA_signal_23048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C ( clk ), .D ( new_AGEMA_signal_23051 ), .Q ( new_AGEMA_signal_23052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C ( clk ), .D ( new_AGEMA_signal_23055 ), .Q ( new_AGEMA_signal_23056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C ( clk ), .D ( new_AGEMA_signal_23059 ), .Q ( new_AGEMA_signal_23060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_23062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C ( clk ), .D ( new_AGEMA_signal_4202 ), .Q ( new_AGEMA_signal_23064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C ( clk ), .D ( new_AGEMA_signal_4203 ), .Q ( new_AGEMA_signal_23066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C ( clk ), .D ( new_AGEMA_signal_4204 ), .Q ( new_AGEMA_signal_23068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C ( clk ), .D ( new_AGEMA_signal_4205 ), .Q ( new_AGEMA_signal_23070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C ( clk ), .D ( new_AGEMA_signal_23077 ), .Q ( new_AGEMA_signal_23078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C ( clk ), .D ( new_AGEMA_signal_23085 ), .Q ( new_AGEMA_signal_23086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C ( clk ), .D ( new_AGEMA_signal_23093 ), .Q ( new_AGEMA_signal_23094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C ( clk ), .D ( new_AGEMA_signal_23101 ), .Q ( new_AGEMA_signal_23102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C ( clk ), .D ( new_AGEMA_signal_23109 ), .Q ( new_AGEMA_signal_23110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C ( clk ), .D ( new_AGEMA_signal_23117 ), .Q ( new_AGEMA_signal_23118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C ( clk ), .D ( new_AGEMA_signal_23125 ), .Q ( new_AGEMA_signal_23126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C ( clk ), .D ( new_AGEMA_signal_23133 ), .Q ( new_AGEMA_signal_23134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C ( clk ), .D ( new_AGEMA_signal_23141 ), .Q ( new_AGEMA_signal_23142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C ( clk ), .D ( new_AGEMA_signal_23149 ), .Q ( new_AGEMA_signal_23150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C ( clk ), .D ( new_AGEMA_signal_23155 ), .Q ( new_AGEMA_signal_23156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C ( clk ), .D ( new_AGEMA_signal_23161 ), .Q ( new_AGEMA_signal_23162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C ( clk ), .D ( new_AGEMA_signal_23167 ), .Q ( new_AGEMA_signal_23168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C ( clk ), .D ( new_AGEMA_signal_23173 ), .Q ( new_AGEMA_signal_23174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C ( clk ), .D ( new_AGEMA_signal_23179 ), .Q ( new_AGEMA_signal_23180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C ( clk ), .D ( new_AGEMA_signal_23183 ), .Q ( new_AGEMA_signal_23184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C ( clk ), .D ( new_AGEMA_signal_23187 ), .Q ( new_AGEMA_signal_23188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C ( clk ), .D ( new_AGEMA_signal_23191 ), .Q ( new_AGEMA_signal_23192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C ( clk ), .D ( new_AGEMA_signal_23195 ), .Q ( new_AGEMA_signal_23196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C ( clk ), .D ( new_AGEMA_signal_23199 ), .Q ( new_AGEMA_signal_23200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C ( clk ), .D ( new_AGEMA_signal_23207 ), .Q ( new_AGEMA_signal_23208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C ( clk ), .D ( new_AGEMA_signal_23215 ), .Q ( new_AGEMA_signal_23216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C ( clk ), .D ( new_AGEMA_signal_23223 ), .Q ( new_AGEMA_signal_23224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C ( clk ), .D ( new_AGEMA_signal_23231 ), .Q ( new_AGEMA_signal_23232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C ( clk ), .D ( new_AGEMA_signal_23239 ), .Q ( new_AGEMA_signal_23240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_23242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C ( clk ), .D ( new_AGEMA_signal_4066 ), .Q ( new_AGEMA_signal_23244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C ( clk ), .D ( new_AGEMA_signal_4067 ), .Q ( new_AGEMA_signal_23246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C ( clk ), .D ( new_AGEMA_signal_4068 ), .Q ( new_AGEMA_signal_23248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C ( clk ), .D ( new_AGEMA_signal_4069 ), .Q ( new_AGEMA_signal_23250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C ( clk ), .D ( new_AGEMA_signal_23253 ), .Q ( new_AGEMA_signal_23254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C ( clk ), .D ( new_AGEMA_signal_23259 ), .Q ( new_AGEMA_signal_23260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C ( clk ), .D ( new_AGEMA_signal_23265 ), .Q ( new_AGEMA_signal_23266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C ( clk ), .D ( new_AGEMA_signal_23271 ), .Q ( new_AGEMA_signal_23272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C ( clk ), .D ( new_AGEMA_signal_23277 ), .Q ( new_AGEMA_signal_23278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C ( clk ), .D ( new_AGEMA_signal_23283 ), .Q ( new_AGEMA_signal_23284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C ( clk ), .D ( new_AGEMA_signal_23289 ), .Q ( new_AGEMA_signal_23290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C ( clk ), .D ( new_AGEMA_signal_23295 ), .Q ( new_AGEMA_signal_23296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C ( clk ), .D ( new_AGEMA_signal_23301 ), .Q ( new_AGEMA_signal_23302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C ( clk ), .D ( new_AGEMA_signal_23307 ), .Q ( new_AGEMA_signal_23308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C ( clk ), .D ( new_AGEMA_signal_23313 ), .Q ( new_AGEMA_signal_23314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C ( clk ), .D ( new_AGEMA_signal_23319 ), .Q ( new_AGEMA_signal_23320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C ( clk ), .D ( new_AGEMA_signal_23325 ), .Q ( new_AGEMA_signal_23326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C ( clk ), .D ( new_AGEMA_signal_23331 ), .Q ( new_AGEMA_signal_23332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C ( clk ), .D ( new_AGEMA_signal_23337 ), .Q ( new_AGEMA_signal_23338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C ( clk ), .D ( new_AGEMA_signal_22443 ), .Q ( new_AGEMA_signal_23342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C ( clk ), .D ( new_AGEMA_signal_22445 ), .Q ( new_AGEMA_signal_23346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C ( clk ), .D ( new_AGEMA_signal_22447 ), .Q ( new_AGEMA_signal_23350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C ( clk ), .D ( new_AGEMA_signal_22449 ), .Q ( new_AGEMA_signal_23354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C ( clk ), .D ( new_AGEMA_signal_22451 ), .Q ( new_AGEMA_signal_23358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C ( clk ), .D ( new_AGEMA_signal_23365 ), .Q ( new_AGEMA_signal_23366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C ( clk ), .D ( new_AGEMA_signal_23373 ), .Q ( new_AGEMA_signal_23374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C ( clk ), .D ( new_AGEMA_signal_23381 ), .Q ( new_AGEMA_signal_23382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C ( clk ), .D ( new_AGEMA_signal_23389 ), .Q ( new_AGEMA_signal_23390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C ( clk ), .D ( new_AGEMA_signal_23397 ), .Q ( new_AGEMA_signal_23398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C ( clk ), .D ( new_AGEMA_signal_23403 ), .Q ( new_AGEMA_signal_23404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C ( clk ), .D ( new_AGEMA_signal_23409 ), .Q ( new_AGEMA_signal_23410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C ( clk ), .D ( new_AGEMA_signal_23415 ), .Q ( new_AGEMA_signal_23416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C ( clk ), .D ( new_AGEMA_signal_23421 ), .Q ( new_AGEMA_signal_23422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C ( clk ), .D ( new_AGEMA_signal_23427 ), .Q ( new_AGEMA_signal_23428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_23432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C ( clk ), .D ( new_AGEMA_signal_3878 ), .Q ( new_AGEMA_signal_23436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C ( clk ), .D ( new_AGEMA_signal_3879 ), .Q ( new_AGEMA_signal_23440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C ( clk ), .D ( new_AGEMA_signal_3880 ), .Q ( new_AGEMA_signal_23444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C ( clk ), .D ( new_AGEMA_signal_3881 ), .Q ( new_AGEMA_signal_23448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C ( clk ), .D ( new_AGEMA_signal_23455 ), .Q ( new_AGEMA_signal_23456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C ( clk ), .D ( new_AGEMA_signal_23463 ), .Q ( new_AGEMA_signal_23464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C ( clk ), .D ( new_AGEMA_signal_23471 ), .Q ( new_AGEMA_signal_23472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C ( clk ), .D ( new_AGEMA_signal_23479 ), .Q ( new_AGEMA_signal_23480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C ( clk ), .D ( new_AGEMA_signal_23487 ), .Q ( new_AGEMA_signal_23488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C ( clk ), .D ( new_AGEMA_signal_23495 ), .Q ( new_AGEMA_signal_23496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C ( clk ), .D ( new_AGEMA_signal_23503 ), .Q ( new_AGEMA_signal_23504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C ( clk ), .D ( new_AGEMA_signal_23511 ), .Q ( new_AGEMA_signal_23512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C ( clk ), .D ( new_AGEMA_signal_23519 ), .Q ( new_AGEMA_signal_23520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C ( clk ), .D ( new_AGEMA_signal_23527 ), .Q ( new_AGEMA_signal_23528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C ( clk ), .D ( new_AGEMA_signal_23537 ), .Q ( new_AGEMA_signal_23538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C ( clk ), .D ( new_AGEMA_signal_23547 ), .Q ( new_AGEMA_signal_23548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C ( clk ), .D ( new_AGEMA_signal_23557 ), .Q ( new_AGEMA_signal_23558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C ( clk ), .D ( new_AGEMA_signal_23567 ), .Q ( new_AGEMA_signal_23568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C ( clk ), .D ( new_AGEMA_signal_23577 ), .Q ( new_AGEMA_signal_23578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C ( clk ), .D ( new_AGEMA_signal_23585 ), .Q ( new_AGEMA_signal_23586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C ( clk ), .D ( new_AGEMA_signal_23593 ), .Q ( new_AGEMA_signal_23594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C ( clk ), .D ( new_AGEMA_signal_23601 ), .Q ( new_AGEMA_signal_23602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C ( clk ), .D ( new_AGEMA_signal_23609 ), .Q ( new_AGEMA_signal_23610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C ( clk ), .D ( new_AGEMA_signal_23617 ), .Q ( new_AGEMA_signal_23618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C ( clk ), .D ( new_AGEMA_signal_23623 ), .Q ( new_AGEMA_signal_23624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C ( clk ), .D ( new_AGEMA_signal_23629 ), .Q ( new_AGEMA_signal_23630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C ( clk ), .D ( new_AGEMA_signal_23635 ), .Q ( new_AGEMA_signal_23636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C ( clk ), .D ( new_AGEMA_signal_23641 ), .Q ( new_AGEMA_signal_23642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C ( clk ), .D ( new_AGEMA_signal_23647 ), .Q ( new_AGEMA_signal_23648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_23652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C ( clk ), .D ( new_AGEMA_signal_3942 ), .Q ( new_AGEMA_signal_23656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C ( clk ), .D ( new_AGEMA_signal_3943 ), .Q ( new_AGEMA_signal_23660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C ( clk ), .D ( new_AGEMA_signal_3944 ), .Q ( new_AGEMA_signal_23664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C ( clk ), .D ( new_AGEMA_signal_3945 ), .Q ( new_AGEMA_signal_23668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C ( clk ), .D ( new_AGEMA_signal_23673 ), .Q ( new_AGEMA_signal_23674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C ( clk ), .D ( new_AGEMA_signal_23679 ), .Q ( new_AGEMA_signal_23680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C ( clk ), .D ( new_AGEMA_signal_23685 ), .Q ( new_AGEMA_signal_23686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C ( clk ), .D ( new_AGEMA_signal_23691 ), .Q ( new_AGEMA_signal_23692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C ( clk ), .D ( new_AGEMA_signal_23697 ), .Q ( new_AGEMA_signal_23698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C ( clk ), .D ( new_AGEMA_signal_23705 ), .Q ( new_AGEMA_signal_23706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C ( clk ), .D ( new_AGEMA_signal_23713 ), .Q ( new_AGEMA_signal_23714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C ( clk ), .D ( new_AGEMA_signal_23721 ), .Q ( new_AGEMA_signal_23722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C ( clk ), .D ( new_AGEMA_signal_23729 ), .Q ( new_AGEMA_signal_23730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C ( clk ), .D ( new_AGEMA_signal_23737 ), .Q ( new_AGEMA_signal_23738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C ( clk ), .D ( new_AGEMA_signal_23743 ), .Q ( new_AGEMA_signal_23744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C ( clk ), .D ( new_AGEMA_signal_23749 ), .Q ( new_AGEMA_signal_23750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C ( clk ), .D ( new_AGEMA_signal_23755 ), .Q ( new_AGEMA_signal_23756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C ( clk ), .D ( new_AGEMA_signal_23761 ), .Q ( new_AGEMA_signal_23762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C ( clk ), .D ( new_AGEMA_signal_23767 ), .Q ( new_AGEMA_signal_23768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C ( clk ), .D ( new_AGEMA_signal_23785 ), .Q ( new_AGEMA_signal_23786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C ( clk ), .D ( new_AGEMA_signal_23793 ), .Q ( new_AGEMA_signal_23794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C ( clk ), .D ( new_AGEMA_signal_23801 ), .Q ( new_AGEMA_signal_23802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C ( clk ), .D ( new_AGEMA_signal_23809 ), .Q ( new_AGEMA_signal_23810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C ( clk ), .D ( new_AGEMA_signal_23817 ), .Q ( new_AGEMA_signal_23818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_23822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C ( clk ), .D ( new_AGEMA_signal_4034 ), .Q ( new_AGEMA_signal_23826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C ( clk ), .D ( new_AGEMA_signal_4035 ), .Q ( new_AGEMA_signal_23830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C ( clk ), .D ( new_AGEMA_signal_4036 ), .Q ( new_AGEMA_signal_23834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C ( clk ), .D ( new_AGEMA_signal_4037 ), .Q ( new_AGEMA_signal_23838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C ( clk ), .D ( new_AGEMA_signal_23843 ), .Q ( new_AGEMA_signal_23844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C ( clk ), .D ( new_AGEMA_signal_23849 ), .Q ( new_AGEMA_signal_23850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C ( clk ), .D ( new_AGEMA_signal_23855 ), .Q ( new_AGEMA_signal_23856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C ( clk ), .D ( new_AGEMA_signal_23861 ), .Q ( new_AGEMA_signal_23862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C ( clk ), .D ( new_AGEMA_signal_23867 ), .Q ( new_AGEMA_signal_23868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C ( clk ), .D ( new_AGEMA_signal_23873 ), .Q ( new_AGEMA_signal_23874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C ( clk ), .D ( new_AGEMA_signal_23879 ), .Q ( new_AGEMA_signal_23880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C ( clk ), .D ( new_AGEMA_signal_23885 ), .Q ( new_AGEMA_signal_23886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C ( clk ), .D ( new_AGEMA_signal_23891 ), .Q ( new_AGEMA_signal_23892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C ( clk ), .D ( new_AGEMA_signal_23897 ), .Q ( new_AGEMA_signal_23898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_23902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C ( clk ), .D ( new_AGEMA_signal_4062 ), .Q ( new_AGEMA_signal_23906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C ( clk ), .D ( new_AGEMA_signal_4063 ), .Q ( new_AGEMA_signal_23910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C ( clk ), .D ( new_AGEMA_signal_4064 ), .Q ( new_AGEMA_signal_23914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C ( clk ), .D ( new_AGEMA_signal_4065 ), .Q ( new_AGEMA_signal_23918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_23922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C ( clk ), .D ( new_AGEMA_signal_3534 ), .Q ( new_AGEMA_signal_23928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C ( clk ), .D ( new_AGEMA_signal_3535 ), .Q ( new_AGEMA_signal_23934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C ( clk ), .D ( new_AGEMA_signal_3536 ), .Q ( new_AGEMA_signal_23940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C ( clk ), .D ( new_AGEMA_signal_3537 ), .Q ( new_AGEMA_signal_23946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_23972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C ( clk ), .D ( new_AGEMA_signal_3886 ), .Q ( new_AGEMA_signal_23978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C ( clk ), .D ( new_AGEMA_signal_3887 ), .Q ( new_AGEMA_signal_23984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C ( clk ), .D ( new_AGEMA_signal_3888 ), .Q ( new_AGEMA_signal_23990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C ( clk ), .D ( new_AGEMA_signal_3889 ), .Q ( new_AGEMA_signal_23996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C ( clk ), .D ( new_AGEMA_signal_24005 ), .Q ( new_AGEMA_signal_24006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C ( clk ), .D ( new_AGEMA_signal_24015 ), .Q ( new_AGEMA_signal_24016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C ( clk ), .D ( new_AGEMA_signal_24025 ), .Q ( new_AGEMA_signal_24026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C ( clk ), .D ( new_AGEMA_signal_24035 ), .Q ( new_AGEMA_signal_24036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C ( clk ), .D ( new_AGEMA_signal_24045 ), .Q ( new_AGEMA_signal_24046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_24052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C ( clk ), .D ( new_AGEMA_signal_4114 ), .Q ( new_AGEMA_signal_24058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C ( clk ), .D ( new_AGEMA_signal_4115 ), .Q ( new_AGEMA_signal_24064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C ( clk ), .D ( new_AGEMA_signal_4116 ), .Q ( new_AGEMA_signal_24070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C ( clk ), .D ( new_AGEMA_signal_4117 ), .Q ( new_AGEMA_signal_24076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_24082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C ( clk ), .D ( new_AGEMA_signal_3606 ), .Q ( new_AGEMA_signal_24088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C ( clk ), .D ( new_AGEMA_signal_3607 ), .Q ( new_AGEMA_signal_24094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C ( clk ), .D ( new_AGEMA_signal_3608 ), .Q ( new_AGEMA_signal_24100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C ( clk ), .D ( new_AGEMA_signal_3609 ), .Q ( new_AGEMA_signal_24106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C ( clk ), .D ( new_AGEMA_signal_24153 ), .Q ( new_AGEMA_signal_24154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C ( clk ), .D ( new_AGEMA_signal_24161 ), .Q ( new_AGEMA_signal_24162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C ( clk ), .D ( new_AGEMA_signal_24169 ), .Q ( new_AGEMA_signal_24170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C ( clk ), .D ( new_AGEMA_signal_24177 ), .Q ( new_AGEMA_signal_24178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C ( clk ), .D ( new_AGEMA_signal_24185 ), .Q ( new_AGEMA_signal_24186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_24192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C ( clk ), .D ( new_AGEMA_signal_3658 ), .Q ( new_AGEMA_signal_24198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C ( clk ), .D ( new_AGEMA_signal_3659 ), .Q ( new_AGEMA_signal_24204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C ( clk ), .D ( new_AGEMA_signal_3660 ), .Q ( new_AGEMA_signal_24210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C ( clk ), .D ( new_AGEMA_signal_3661 ), .Q ( new_AGEMA_signal_24216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C ( clk ), .D ( new_AGEMA_signal_24223 ), .Q ( new_AGEMA_signal_24224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C ( clk ), .D ( new_AGEMA_signal_24231 ), .Q ( new_AGEMA_signal_24232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C ( clk ), .D ( new_AGEMA_signal_24239 ), .Q ( new_AGEMA_signal_24240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C ( clk ), .D ( new_AGEMA_signal_24247 ), .Q ( new_AGEMA_signal_24248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C ( clk ), .D ( new_AGEMA_signal_24255 ), .Q ( new_AGEMA_signal_24256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C ( clk ), .D ( new_AGEMA_signal_24263 ), .Q ( new_AGEMA_signal_24264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C ( clk ), .D ( new_AGEMA_signal_24271 ), .Q ( new_AGEMA_signal_24272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C ( clk ), .D ( new_AGEMA_signal_24279 ), .Q ( new_AGEMA_signal_24280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C ( clk ), .D ( new_AGEMA_signal_24287 ), .Q ( new_AGEMA_signal_24288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C ( clk ), .D ( new_AGEMA_signal_24295 ), .Q ( new_AGEMA_signal_24296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C ( clk ), .D ( new_AGEMA_signal_24353 ), .Q ( new_AGEMA_signal_24354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C ( clk ), .D ( new_AGEMA_signal_24361 ), .Q ( new_AGEMA_signal_24362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C ( clk ), .D ( new_AGEMA_signal_24369 ), .Q ( new_AGEMA_signal_24370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C ( clk ), .D ( new_AGEMA_signal_24377 ), .Q ( new_AGEMA_signal_24378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C ( clk ), .D ( new_AGEMA_signal_24385 ), .Q ( new_AGEMA_signal_24386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_24412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C ( clk ), .D ( new_AGEMA_signal_3858 ), .Q ( new_AGEMA_signal_24420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C ( clk ), .D ( new_AGEMA_signal_3859 ), .Q ( new_AGEMA_signal_24428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C ( clk ), .D ( new_AGEMA_signal_3860 ), .Q ( new_AGEMA_signal_24436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7669 ( .C ( clk ), .D ( new_AGEMA_signal_3861 ), .Q ( new_AGEMA_signal_24444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7681 ( .C ( clk ), .D ( new_AGEMA_signal_24455 ), .Q ( new_AGEMA_signal_24456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7693 ( .C ( clk ), .D ( new_AGEMA_signal_24467 ), .Q ( new_AGEMA_signal_24468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7705 ( .C ( clk ), .D ( new_AGEMA_signal_24479 ), .Q ( new_AGEMA_signal_24480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7717 ( .C ( clk ), .D ( new_AGEMA_signal_24491 ), .Q ( new_AGEMA_signal_24492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7729 ( .C ( clk ), .D ( new_AGEMA_signal_24503 ), .Q ( new_AGEMA_signal_24504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7743 ( .C ( clk ), .D ( new_AGEMA_signal_24517 ), .Q ( new_AGEMA_signal_24518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7757 ( .C ( clk ), .D ( new_AGEMA_signal_24531 ), .Q ( new_AGEMA_signal_24532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7771 ( .C ( clk ), .D ( new_AGEMA_signal_24545 ), .Q ( new_AGEMA_signal_24546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7785 ( .C ( clk ), .D ( new_AGEMA_signal_24559 ), .Q ( new_AGEMA_signal_24560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7799 ( .C ( clk ), .D ( new_AGEMA_signal_24573 ), .Q ( new_AGEMA_signal_24574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7807 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_24582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7815 ( .C ( clk ), .D ( new_AGEMA_signal_4138 ), .Q ( new_AGEMA_signal_24590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7823 ( .C ( clk ), .D ( new_AGEMA_signal_4139 ), .Q ( new_AGEMA_signal_24598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7831 ( .C ( clk ), .D ( new_AGEMA_signal_4140 ), .Q ( new_AGEMA_signal_24606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7839 ( .C ( clk ), .D ( new_AGEMA_signal_4141 ), .Q ( new_AGEMA_signal_24614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7853 ( .C ( clk ), .D ( new_AGEMA_signal_24627 ), .Q ( new_AGEMA_signal_24628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7867 ( .C ( clk ), .D ( new_AGEMA_signal_24641 ), .Q ( new_AGEMA_signal_24642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7881 ( .C ( clk ), .D ( new_AGEMA_signal_24655 ), .Q ( new_AGEMA_signal_24656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7895 ( .C ( clk ), .D ( new_AGEMA_signal_24669 ), .Q ( new_AGEMA_signal_24670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7909 ( .C ( clk ), .D ( new_AGEMA_signal_24683 ), .Q ( new_AGEMA_signal_24684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7917 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_24692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7925 ( .C ( clk ), .D ( new_AGEMA_signal_3990 ), .Q ( new_AGEMA_signal_24700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7933 ( .C ( clk ), .D ( new_AGEMA_signal_3991 ), .Q ( new_AGEMA_signal_24708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7941 ( .C ( clk ), .D ( new_AGEMA_signal_3992 ), .Q ( new_AGEMA_signal_24716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7949 ( .C ( clk ), .D ( new_AGEMA_signal_3993 ), .Q ( new_AGEMA_signal_24724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7957 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_24732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7965 ( .C ( clk ), .D ( new_AGEMA_signal_4050 ), .Q ( new_AGEMA_signal_24740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7973 ( .C ( clk ), .D ( new_AGEMA_signal_4051 ), .Q ( new_AGEMA_signal_24748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7981 ( .C ( clk ), .D ( new_AGEMA_signal_4052 ), .Q ( new_AGEMA_signal_24756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7989 ( .C ( clk ), .D ( new_AGEMA_signal_4053 ), .Q ( new_AGEMA_signal_24764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8033 ( .C ( clk ), .D ( new_AGEMA_signal_24807 ), .Q ( new_AGEMA_signal_24808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8049 ( .C ( clk ), .D ( new_AGEMA_signal_24823 ), .Q ( new_AGEMA_signal_24824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8065 ( .C ( clk ), .D ( new_AGEMA_signal_24839 ), .Q ( new_AGEMA_signal_24840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8081 ( .C ( clk ), .D ( new_AGEMA_signal_24855 ), .Q ( new_AGEMA_signal_24856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8097 ( .C ( clk ), .D ( new_AGEMA_signal_24871 ), .Q ( new_AGEMA_signal_24872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8143 ( .C ( clk ), .D ( new_AGEMA_signal_24917 ), .Q ( new_AGEMA_signal_24918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8159 ( .C ( clk ), .D ( new_AGEMA_signal_24933 ), .Q ( new_AGEMA_signal_24934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8175 ( .C ( clk ), .D ( new_AGEMA_signal_24949 ), .Q ( new_AGEMA_signal_24950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8191 ( .C ( clk ), .D ( new_AGEMA_signal_24965 ), .Q ( new_AGEMA_signal_24966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8207 ( .C ( clk ), .D ( new_AGEMA_signal_24981 ), .Q ( new_AGEMA_signal_24982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8217 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_24992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8227 ( .C ( clk ), .D ( new_AGEMA_signal_4206 ), .Q ( new_AGEMA_signal_25002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8237 ( .C ( clk ), .D ( new_AGEMA_signal_4207 ), .Q ( new_AGEMA_signal_25012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8247 ( .C ( clk ), .D ( new_AGEMA_signal_4208 ), .Q ( new_AGEMA_signal_25022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8257 ( .C ( clk ), .D ( new_AGEMA_signal_4209 ), .Q ( new_AGEMA_signal_25032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8391 ( .C ( clk ), .D ( new_AGEMA_signal_25165 ), .Q ( new_AGEMA_signal_25166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8407 ( .C ( clk ), .D ( new_AGEMA_signal_25181 ), .Q ( new_AGEMA_signal_25182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8423 ( .C ( clk ), .D ( new_AGEMA_signal_25197 ), .Q ( new_AGEMA_signal_25198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8439 ( .C ( clk ), .D ( new_AGEMA_signal_25213 ), .Q ( new_AGEMA_signal_25214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8455 ( .C ( clk ), .D ( new_AGEMA_signal_25229 ), .Q ( new_AGEMA_signal_25230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8523 ( .C ( clk ), .D ( new_AGEMA_signal_25297 ), .Q ( new_AGEMA_signal_25298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8541 ( .C ( clk ), .D ( new_AGEMA_signal_25315 ), .Q ( new_AGEMA_signal_25316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8559 ( .C ( clk ), .D ( new_AGEMA_signal_25333 ), .Q ( new_AGEMA_signal_25334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8577 ( .C ( clk ), .D ( new_AGEMA_signal_25351 ), .Q ( new_AGEMA_signal_25352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8595 ( .C ( clk ), .D ( new_AGEMA_signal_25369 ), .Q ( new_AGEMA_signal_25370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8773 ( .C ( clk ), .D ( new_AGEMA_signal_25547 ), .Q ( new_AGEMA_signal_25548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8793 ( .C ( clk ), .D ( new_AGEMA_signal_25567 ), .Q ( new_AGEMA_signal_25568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8813 ( .C ( clk ), .D ( new_AGEMA_signal_25587 ), .Q ( new_AGEMA_signal_25588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8833 ( .C ( clk ), .D ( new_AGEMA_signal_25607 ), .Q ( new_AGEMA_signal_25608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8853 ( .C ( clk ), .D ( new_AGEMA_signal_25627 ), .Q ( new_AGEMA_signal_25628 ) ) ;

    /* cells in depth 14 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2002 ( .ina ({new_AGEMA_signal_21581, new_AGEMA_signal_21579, new_AGEMA_signal_21577, new_AGEMA_signal_21575, new_AGEMA_signal_21573}), .inb ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, new_AGEMA_signal_3843, new_AGEMA_signal_3842, n1933}), .clk ( clk ), .rnd ({Fresh[10859], Fresh[10858], Fresh[10857], Fresh[10856], Fresh[10855], Fresh[10854], Fresh[10853], Fresh[10852], Fresh[10851], Fresh[10850], Fresh[10849], Fresh[10848], Fresh[10847], Fresh[10846], Fresh[10845]}), .outt ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, new_AGEMA_signal_4079, new_AGEMA_signal_4078, n1935}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2054 ( .ina ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, n1958}), .inb ({new_AGEMA_signal_21621, new_AGEMA_signal_21613, new_AGEMA_signal_21605, new_AGEMA_signal_21597, new_AGEMA_signal_21589}), .clk ( clk ), .rnd ({Fresh[10874], Fresh[10873], Fresh[10872], Fresh[10871], Fresh[10870], Fresh[10869], Fresh[10868], Fresh[10867], Fresh[10866], Fresh[10865], Fresh[10864], Fresh[10863], Fresh[10862], Fresh[10861], Fresh[10860]}), .outt ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, new_AGEMA_signal_4083, new_AGEMA_signal_4082, n1959}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2109 ( .ina ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, new_AGEMA_signal_3854, n1982}), .inb ({new_AGEMA_signal_21631, new_AGEMA_signal_21629, new_AGEMA_signal_21627, new_AGEMA_signal_21625, new_AGEMA_signal_21623}), .clk ( clk ), .rnd ({Fresh[10889], Fresh[10888], Fresh[10887], Fresh[10886], Fresh[10885], Fresh[10884], Fresh[10883], Fresh[10882], Fresh[10881], Fresh[10880], Fresh[10879], Fresh[10878], Fresh[10877], Fresh[10876], Fresh[10875]}), .outt ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, new_AGEMA_signal_4086, n1983}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2149 ( .ina ({new_AGEMA_signal_21651, new_AGEMA_signal_21647, new_AGEMA_signal_21643, new_AGEMA_signal_21639, new_AGEMA_signal_21635}), .inb ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, new_AGEMA_signal_3863, new_AGEMA_signal_3862, n2011}), .clk ( clk ), .rnd ({Fresh[10904], Fresh[10903], Fresh[10902], Fresh[10901], Fresh[10900], Fresh[10899], Fresh[10898], Fresh[10897], Fresh[10896], Fresh[10895], Fresh[10894], Fresh[10893], Fresh[10892], Fresh[10891], Fresh[10890]}), .outt ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, new_AGEMA_signal_4091, new_AGEMA_signal_4090, n2014}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2166 ( .ina ({new_AGEMA_signal_21691, new_AGEMA_signal_21683, new_AGEMA_signal_21675, new_AGEMA_signal_21667, new_AGEMA_signal_21659}), .inb ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2025}), .clk ( clk ), .rnd ({Fresh[10919], Fresh[10918], Fresh[10917], Fresh[10916], Fresh[10915], Fresh[10914], Fresh[10913], Fresh[10912], Fresh[10911], Fresh[10910], Fresh[10909], Fresh[10908], Fresh[10907], Fresh[10906], Fresh[10905]}), .outt ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, new_AGEMA_signal_3866, n2029}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2180 ( .ina ({new_AGEMA_signal_21701, new_AGEMA_signal_21699, new_AGEMA_signal_21697, new_AGEMA_signal_21695, new_AGEMA_signal_21693}), .inb ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, n2036}), .clk ( clk ), .rnd ({Fresh[10934], Fresh[10933], Fresh[10932], Fresh[10931], Fresh[10930], Fresh[10929], Fresh[10928], Fresh[10927], Fresh[10926], Fresh[10925], Fresh[10924], Fresh[10923], Fresh[10922], Fresh[10921], Fresh[10920]}), .outt ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, new_AGEMA_signal_4099, new_AGEMA_signal_4098, n2037}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2197 ( .ina ({new_AGEMA_signal_21731, new_AGEMA_signal_21725, new_AGEMA_signal_21719, new_AGEMA_signal_21713, new_AGEMA_signal_21707}), .inb ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, new_AGEMA_signal_3875, new_AGEMA_signal_3874, n2049}), .clk ( clk ), .rnd ({Fresh[10949], Fresh[10948], Fresh[10947], Fresh[10946], Fresh[10945], Fresh[10944], Fresh[10943], Fresh[10942], Fresh[10941], Fresh[10940], Fresh[10939], Fresh[10938], Fresh[10937], Fresh[10936], Fresh[10935]}), .outt ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, new_AGEMA_signal_4102, n2052}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2219 ( .ina ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, n2067}), .inb ({new_AGEMA_signal_21751, new_AGEMA_signal_21747, new_AGEMA_signal_21743, new_AGEMA_signal_21739, new_AGEMA_signal_21735}), .clk ( clk ), .rnd ({Fresh[10964], Fresh[10963], Fresh[10962], Fresh[10961], Fresh[10960], Fresh[10959], Fresh[10958], Fresh[10957], Fresh[10956], Fresh[10955], Fresh[10954], Fresh[10953], Fresh[10952], Fresh[10951], Fresh[10950]}), .outt ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, new_AGEMA_signal_4107, new_AGEMA_signal_4106, n2070}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2258 ( .ina ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, new_AGEMA_signal_3890, n2097}), .inb ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, n2096}), .clk ( clk ), .rnd ({Fresh[10979], Fresh[10978], Fresh[10977], Fresh[10976], Fresh[10975], Fresh[10974], Fresh[10973], Fresh[10972], Fresh[10971], Fresh[10970], Fresh[10969], Fresh[10968], Fresh[10967], Fresh[10966], Fresh[10965]}), .outt ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, new_AGEMA_signal_4110, n2098}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2287 ( .ina ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, new_AGEMA_signal_3902, n2124}), .inb ({new_AGEMA_signal_21791, new_AGEMA_signal_21783, new_AGEMA_signal_21775, new_AGEMA_signal_21767, new_AGEMA_signal_21759}), .clk ( clk ), .rnd ({Fresh[10994], Fresh[10993], Fresh[10992], Fresh[10991], Fresh[10990], Fresh[10989], Fresh[10988], Fresh[10987], Fresh[10986], Fresh[10985], Fresh[10984], Fresh[10983], Fresh[10982], Fresh[10981], Fresh[10980]}), .outt ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, new_AGEMA_signal_4119, new_AGEMA_signal_4118, n2125}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2311 ( .ina ({new_AGEMA_signal_21811, new_AGEMA_signal_21807, new_AGEMA_signal_21803, new_AGEMA_signal_21799, new_AGEMA_signal_21795}), .inb ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, new_AGEMA_signal_3906, n2142}), .clk ( clk ), .rnd ({Fresh[11009], Fresh[11008], Fresh[11007], Fresh[11006], Fresh[11005], Fresh[11004], Fresh[11003], Fresh[11002], Fresh[11001], Fresh[11000], Fresh[10999], Fresh[10998], Fresh[10997], Fresh[10996], Fresh[10995]}), .outt ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, new_AGEMA_signal_4122, n2145}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2333 ( .ina ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, new_AGEMA_signal_3911, new_AGEMA_signal_3910, n2168}), .inb ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, new_AGEMA_signal_3914, n2167}), .clk ( clk ), .rnd ({Fresh[11024], Fresh[11023], Fresh[11022], Fresh[11021], Fresh[11020], Fresh[11019], Fresh[11018], Fresh[11017], Fresh[11016], Fresh[11015], Fresh[11014], Fresh[11013], Fresh[11012], Fresh[11011], Fresh[11010]}), .outt ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, new_AGEMA_signal_4127, new_AGEMA_signal_4126, n2169}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2350 ( .ina ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, new_AGEMA_signal_3918, n2184}), .inb ({new_AGEMA_signal_21841, new_AGEMA_signal_21835, new_AGEMA_signal_21829, new_AGEMA_signal_21823, new_AGEMA_signal_21817}), .clk ( clk ), .rnd ({Fresh[11039], Fresh[11038], Fresh[11037], Fresh[11036], Fresh[11035], Fresh[11034], Fresh[11033], Fresh[11032], Fresh[11031], Fresh[11030], Fresh[11029], Fresh[11028], Fresh[11027], Fresh[11026], Fresh[11025]}), .outt ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, n2185}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2365 ( .ina ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, n2197}), .inb ({new_AGEMA_signal_21871, new_AGEMA_signal_21865, new_AGEMA_signal_21859, new_AGEMA_signal_21853, new_AGEMA_signal_21847}), .clk ( clk ), .rnd ({Fresh[11054], Fresh[11053], Fresh[11052], Fresh[11051], Fresh[11050], Fresh[11049], Fresh[11048], Fresh[11047], Fresh[11046], Fresh[11045], Fresh[11044], Fresh[11043], Fresh[11042], Fresh[11041], Fresh[11040]}), .outt ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, new_AGEMA_signal_4135, new_AGEMA_signal_4134, n2198}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2396 ( .ina ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, new_AGEMA_signal_3930, n2232}), .inb ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, n2231}), .clk ( clk ), .rnd ({Fresh[11069], Fresh[11068], Fresh[11067], Fresh[11066], Fresh[11065], Fresh[11064], Fresh[11063], Fresh[11062], Fresh[11061], Fresh[11060], Fresh[11059], Fresh[11058], Fresh[11057], Fresh[11056], Fresh[11055]}), .outt ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, new_AGEMA_signal_4143, new_AGEMA_signal_4142, n2312}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2404 ( .ina ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, new_AGEMA_signal_4146, n2239}), .inb ({new_AGEMA_signal_21901, new_AGEMA_signal_21895, new_AGEMA_signal_21889, new_AGEMA_signal_21883, new_AGEMA_signal_21877}), .clk ( clk ), .rnd ({Fresh[11084], Fresh[11083], Fresh[11082], Fresh[11081], Fresh[11080], Fresh[11079], Fresh[11078], Fresh[11077], Fresh[11076], Fresh[11075], Fresh[11074], Fresh[11073], Fresh[11072], Fresh[11071], Fresh[11070]}), .outt ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, new_AGEMA_signal_4299, new_AGEMA_signal_4298, n2258}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2415 ( .ina ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, new_AGEMA_signal_3938, n2250}), .inb ({new_AGEMA_signal_21931, new_AGEMA_signal_21925, new_AGEMA_signal_21919, new_AGEMA_signal_21913, new_AGEMA_signal_21907}), .clk ( clk ), .rnd ({Fresh[11099], Fresh[11098], Fresh[11097], Fresh[11096], Fresh[11095], Fresh[11094], Fresh[11093], Fresh[11092], Fresh[11091], Fresh[11090], Fresh[11089], Fresh[11088], Fresh[11087], Fresh[11086], Fresh[11085]}), .outt ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, new_AGEMA_signal_4151, new_AGEMA_signal_4150, n2251}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2440 ( .ina ({new_AGEMA_signal_21961, new_AGEMA_signal_21955, new_AGEMA_signal_21949, new_AGEMA_signal_21943, new_AGEMA_signal_21937}), .inb ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, n2272}), .clk ( clk ), .rnd ({Fresh[11114], Fresh[11113], Fresh[11112], Fresh[11111], Fresh[11110], Fresh[11109], Fresh[11108], Fresh[11107], Fresh[11106], Fresh[11105], Fresh[11104], Fresh[11103], Fresh[11102], Fresh[11101], Fresh[11100]}), .outt ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, new_AGEMA_signal_4155, new_AGEMA_signal_4154, n2274}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2469 ( .ina ({new_AGEMA_signal_21981, new_AGEMA_signal_21977, new_AGEMA_signal_21973, new_AGEMA_signal_21969, new_AGEMA_signal_21965}), .inb ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, new_AGEMA_signal_3950, n2296}), .clk ( clk ), .rnd ({Fresh[11129], Fresh[11128], Fresh[11127], Fresh[11126], Fresh[11125], Fresh[11124], Fresh[11123], Fresh[11122], Fresh[11121], Fresh[11120], Fresh[11119], Fresh[11118], Fresh[11117], Fresh[11116], Fresh[11115]}), .outt ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, new_AGEMA_signal_4158, n2302}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2490 ( .ina ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, new_AGEMA_signal_3954, n2324}), .inb ({new_AGEMA_signal_22021, new_AGEMA_signal_22013, new_AGEMA_signal_22005, new_AGEMA_signal_21997, new_AGEMA_signal_21989}), .clk ( clk ), .rnd ({Fresh[11144], Fresh[11143], Fresh[11142], Fresh[11141], Fresh[11140], Fresh[11139], Fresh[11138], Fresh[11137], Fresh[11136], Fresh[11135], Fresh[11134], Fresh[11133], Fresh[11132], Fresh[11131], Fresh[11130]}), .outt ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, new_AGEMA_signal_4163, new_AGEMA_signal_4162, n2339}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2503 ( .ina ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, new_AGEMA_signal_3959, new_AGEMA_signal_3958, n2337}), .inb ({new_AGEMA_signal_22041, new_AGEMA_signal_22037, new_AGEMA_signal_22033, new_AGEMA_signal_22029, new_AGEMA_signal_22025}), .clk ( clk ), .rnd ({Fresh[11159], Fresh[11158], Fresh[11157], Fresh[11156], Fresh[11155], Fresh[11154], Fresh[11153], Fresh[11152], Fresh[11151], Fresh[11150], Fresh[11149], Fresh[11148], Fresh[11147], Fresh[11146], Fresh[11145]}), .outt ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, n2338}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2515 ( .ina ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, new_AGEMA_signal_3962, n2350}), .inb ({new_AGEMA_signal_22071, new_AGEMA_signal_22065, new_AGEMA_signal_22059, new_AGEMA_signal_22053, new_AGEMA_signal_22047}), .clk ( clk ), .rnd ({Fresh[11174], Fresh[11173], Fresh[11172], Fresh[11171], Fresh[11170], Fresh[11169], Fresh[11168], Fresh[11167], Fresh[11166], Fresh[11165], Fresh[11164], Fresh[11163], Fresh[11162], Fresh[11161], Fresh[11160]}), .outt ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, new_AGEMA_signal_4170, n2351}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2529 ( .ina ({new_AGEMA_signal_22111, new_AGEMA_signal_22103, new_AGEMA_signal_22095, new_AGEMA_signal_22087, new_AGEMA_signal_22079}), .inb ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, new_AGEMA_signal_3966, n2362}), .clk ( clk ), .rnd ({Fresh[11189], Fresh[11188], Fresh[11187], Fresh[11186], Fresh[11185], Fresh[11184], Fresh[11183], Fresh[11182], Fresh[11181], Fresh[11180], Fresh[11179], Fresh[11178], Fresh[11177], Fresh[11176], Fresh[11175]}), .outt ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, new_AGEMA_signal_4174, n2365}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2551 ( .ina ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2389}), .inb ({new_AGEMA_signal_22121, new_AGEMA_signal_22119, new_AGEMA_signal_22117, new_AGEMA_signal_22115, new_AGEMA_signal_22113}), .clk ( clk ), .rnd ({Fresh[11204], Fresh[11203], Fresh[11202], Fresh[11201], Fresh[11200], Fresh[11199], Fresh[11198], Fresh[11197], Fresh[11196], Fresh[11195], Fresh[11194], Fresh[11193], Fresh[11192], Fresh[11191], Fresh[11190]}), .outt ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, new_AGEMA_signal_3971, new_AGEMA_signal_3970, n2399}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2560 ( .ina ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, new_AGEMA_signal_3974, n2397}), .inb ({new_AGEMA_signal_22151, new_AGEMA_signal_22145, new_AGEMA_signal_22139, new_AGEMA_signal_22133, new_AGEMA_signal_22127}), .clk ( clk ), .rnd ({Fresh[11219], Fresh[11218], Fresh[11217], Fresh[11216], Fresh[11215], Fresh[11214], Fresh[11213], Fresh[11212], Fresh[11211], Fresh[11210], Fresh[11209], Fresh[11208], Fresh[11207], Fresh[11206], Fresh[11205]}), .outt ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, new_AGEMA_signal_4179, new_AGEMA_signal_4178, n2398}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2572 ( .ina ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, n2411}), .inb ({new_AGEMA_signal_22161, new_AGEMA_signal_22159, new_AGEMA_signal_22157, new_AGEMA_signal_22155, new_AGEMA_signal_22153}), .clk ( clk ), .rnd ({Fresh[11234], Fresh[11233], Fresh[11232], Fresh[11231], Fresh[11230], Fresh[11229], Fresh[11228], Fresh[11227], Fresh[11226], Fresh[11225], Fresh[11224], Fresh[11223], Fresh[11222], Fresh[11221], Fresh[11220]}), .outt ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, new_AGEMA_signal_3979, new_AGEMA_signal_3978, n2423}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2581 ( .ina ({new_AGEMA_signal_22171, new_AGEMA_signal_22169, new_AGEMA_signal_22167, new_AGEMA_signal_22165, new_AGEMA_signal_22163}), .inb ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, n2420}), .clk ( clk ), .rnd ({Fresh[11249], Fresh[11248], Fresh[11247], Fresh[11246], Fresh[11245], Fresh[11244], Fresh[11243], Fresh[11242], Fresh[11241], Fresh[11240], Fresh[11239], Fresh[11238], Fresh[11237], Fresh[11236], Fresh[11235]}), .outt ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, new_AGEMA_signal_3983, new_AGEMA_signal_3982, n2422}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2596 ( .ina ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, new_AGEMA_signal_3986, n2440}), .inb ({new_AGEMA_signal_22201, new_AGEMA_signal_22195, new_AGEMA_signal_22189, new_AGEMA_signal_22183, new_AGEMA_signal_22177}), .clk ( clk ), .rnd ({Fresh[11264], Fresh[11263], Fresh[11262], Fresh[11261], Fresh[11260], Fresh[11259], Fresh[11258], Fresh[11257], Fresh[11256], Fresh[11255], Fresh[11254], Fresh[11253], Fresh[11252], Fresh[11251], Fresh[11250]}), .outt ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, new_AGEMA_signal_4187, new_AGEMA_signal_4186, n2441}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2623 ( .ina ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, new_AGEMA_signal_3731, new_AGEMA_signal_3730, n2471}), .inb ({new_AGEMA_signal_22231, new_AGEMA_signal_22225, new_AGEMA_signal_22219, new_AGEMA_signal_22213, new_AGEMA_signal_22207}), .clk ( clk ), .rnd ({Fresh[11279], Fresh[11278], Fresh[11277], Fresh[11276], Fresh[11275], Fresh[11274], Fresh[11273], Fresh[11272], Fresh[11271], Fresh[11270], Fresh[11269], Fresh[11268], Fresh[11267], Fresh[11266], Fresh[11265]}), .outt ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, new_AGEMA_signal_3994, n2479}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2637 ( .ina ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, new_AGEMA_signal_3998, n2485}), .inb ({new_AGEMA_signal_22271, new_AGEMA_signal_22263, new_AGEMA_signal_22255, new_AGEMA_signal_22247, new_AGEMA_signal_22239}), .clk ( clk ), .rnd ({Fresh[11294], Fresh[11293], Fresh[11292], Fresh[11291], Fresh[11290], Fresh[11289], Fresh[11288], Fresh[11287], Fresh[11286], Fresh[11285], Fresh[11284], Fresh[11283], Fresh[11282], Fresh[11281], Fresh[11280]}), .outt ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, new_AGEMA_signal_4194, n2512}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2652 ( .ina ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, n2502}), .inb ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, new_AGEMA_signal_4003, new_AGEMA_signal_4002, n2501}), .clk ( clk ), .rnd ({Fresh[11309], Fresh[11308], Fresh[11307], Fresh[11306], Fresh[11305], Fresh[11304], Fresh[11303], Fresh[11302], Fresh[11301], Fresh[11300], Fresh[11299], Fresh[11298], Fresh[11297], Fresh[11296], Fresh[11295]}), .outt ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, new_AGEMA_signal_4199, new_AGEMA_signal_4198, n2510}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2686 ( .ina ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, new_AGEMA_signal_4015, new_AGEMA_signal_4014, n2550}), .inb ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, new_AGEMA_signal_4019, new_AGEMA_signal_4018, n2549}), .clk ( clk ), .rnd ({Fresh[11324], Fresh[11323], Fresh[11322], Fresh[11321], Fresh[11320], Fresh[11319], Fresh[11318], Fresh[11317], Fresh[11316], Fresh[11315], Fresh[11314], Fresh[11313], Fresh[11312], Fresh[11311], Fresh[11310]}), .outt ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, new_AGEMA_signal_4210, n2552}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2702 ( .ina ({new_AGEMA_signal_22311, new_AGEMA_signal_22303, new_AGEMA_signal_22295, new_AGEMA_signal_22287, new_AGEMA_signal_22279}), .inb ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, new_AGEMA_signal_4022, n2569}), .clk ( clk ), .rnd ({Fresh[11339], Fresh[11338], Fresh[11337], Fresh[11336], Fresh[11335], Fresh[11334], Fresh[11333], Fresh[11332], Fresh[11331], Fresh[11330], Fresh[11329], Fresh[11328], Fresh[11327], Fresh[11326], Fresh[11325]}), .outt ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, new_AGEMA_signal_4215, new_AGEMA_signal_4214, n2593}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2713 ( .ina ({new_AGEMA_signal_22341, new_AGEMA_signal_22335, new_AGEMA_signal_22329, new_AGEMA_signal_22323, new_AGEMA_signal_22317}), .inb ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, n2584}), .clk ( clk ), .rnd ({Fresh[11354], Fresh[11353], Fresh[11352], Fresh[11351], Fresh[11350], Fresh[11349], Fresh[11348], Fresh[11347], Fresh[11346], Fresh[11345], Fresh[11344], Fresh[11343], Fresh[11342], Fresh[11341], Fresh[11340]}), .outt ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, new_AGEMA_signal_4218, n2589}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2730 ( .ina ({new_AGEMA_signal_22371, new_AGEMA_signal_22365, new_AGEMA_signal_22359, new_AGEMA_signal_22353, new_AGEMA_signal_22347}), .inb ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, n2606}), .clk ( clk ), .rnd ({Fresh[11369], Fresh[11368], Fresh[11367], Fresh[11366], Fresh[11365], Fresh[11364], Fresh[11363], Fresh[11362], Fresh[11361], Fresh[11360], Fresh[11359], Fresh[11358], Fresh[11357], Fresh[11356], Fresh[11355]}), .outt ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, new_AGEMA_signal_4030, n2608}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2748 ( .ina ({new_AGEMA_signal_22381, new_AGEMA_signal_22379, new_AGEMA_signal_22377, new_AGEMA_signal_22375, new_AGEMA_signal_22373}), .inb ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, n2634}), .clk ( clk ), .rnd ({Fresh[11384], Fresh[11383], Fresh[11382], Fresh[11381], Fresh[11380], Fresh[11379], Fresh[11378], Fresh[11377], Fresh[11376], Fresh[11375], Fresh[11374], Fresh[11373], Fresh[11372], Fresh[11371], Fresh[11370]}), .outt ({new_AGEMA_signal_4229, new_AGEMA_signal_4228, new_AGEMA_signal_4227, new_AGEMA_signal_4226, n2636}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2762 ( .ina ({new_AGEMA_signal_22401, new_AGEMA_signal_22397, new_AGEMA_signal_22393, new_AGEMA_signal_22389, new_AGEMA_signal_22385}), .inb ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, new_AGEMA_signal_4043, new_AGEMA_signal_4042, n2657}), .clk ( clk ), .rnd ({Fresh[11399], Fresh[11398], Fresh[11397], Fresh[11396], Fresh[11395], Fresh[11394], Fresh[11393], Fresh[11392], Fresh[11391], Fresh[11390], Fresh[11389], Fresh[11388], Fresh[11387], Fresh[11386], Fresh[11385]}), .outt ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, new_AGEMA_signal_4230, n2659}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2784 ( .ina ({new_AGEMA_signal_22421, new_AGEMA_signal_22417, new_AGEMA_signal_22413, new_AGEMA_signal_22409, new_AGEMA_signal_22405}), .inb ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, new_AGEMA_signal_4047, new_AGEMA_signal_4046, n2697}), .clk ( clk ), .rnd ({Fresh[11414], Fresh[11413], Fresh[11412], Fresh[11411], Fresh[11410], Fresh[11409], Fresh[11408], Fresh[11407], Fresh[11406], Fresh[11405], Fresh[11404], Fresh[11403], Fresh[11402], Fresh[11401], Fresh[11400]}), .outt ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, new_AGEMA_signal_4235, new_AGEMA_signal_4234, n2702}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2811 ( .ina ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, new_AGEMA_signal_4055, new_AGEMA_signal_4054, n2747}), .inb ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, new_AGEMA_signal_4059, new_AGEMA_signal_4058, n2746}), .clk ( clk ), .rnd ({Fresh[11429], Fresh[11428], Fresh[11427], Fresh[11426], Fresh[11425], Fresh[11424], Fresh[11423], Fresh[11422], Fresh[11421], Fresh[11420], Fresh[11419], Fresh[11418], Fresh[11417], Fresh[11416], Fresh[11415]}), .outt ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, new_AGEMA_signal_4239, new_AGEMA_signal_4238, n2806}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2839 ( .ina ({new_AGEMA_signal_22441, new_AGEMA_signal_22437, new_AGEMA_signal_22433, new_AGEMA_signal_22429, new_AGEMA_signal_22425}), .inb ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, n2799}), .clk ( clk ), .rnd ({Fresh[11444], Fresh[11443], Fresh[11442], Fresh[11441], Fresh[11440], Fresh[11439], Fresh[11438], Fresh[11437], Fresh[11436], Fresh[11435], Fresh[11434], Fresh[11433], Fresh[11432], Fresh[11431], Fresh[11430]}), .outt ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, new_AGEMA_signal_4071, new_AGEMA_signal_4070, n2801}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2853 ( .ina ({new_AGEMA_signal_22451, new_AGEMA_signal_22449, new_AGEMA_signal_22447, new_AGEMA_signal_22445, new_AGEMA_signal_22443}), .inb ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, new_AGEMA_signal_4074, n2827}), .clk ( clk ), .rnd ({Fresh[11459], Fresh[11458], Fresh[11457], Fresh[11456], Fresh[11455], Fresh[11454], Fresh[11453], Fresh[11452], Fresh[11451], Fresh[11450], Fresh[11449], Fresh[11448], Fresh[11447], Fresh[11446], Fresh[11445]}), .outt ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, new_AGEMA_signal_4247, new_AGEMA_signal_4246, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C ( clk ), .D ( new_AGEMA_signal_22456 ), .Q ( new_AGEMA_signal_22457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C ( clk ), .D ( new_AGEMA_signal_22462 ), .Q ( new_AGEMA_signal_22463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C ( clk ), .D ( new_AGEMA_signal_22468 ), .Q ( new_AGEMA_signal_22469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C ( clk ), .D ( new_AGEMA_signal_22474 ), .Q ( new_AGEMA_signal_22475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C ( clk ), .D ( new_AGEMA_signal_22480 ), .Q ( new_AGEMA_signal_22481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C ( clk ), .D ( new_AGEMA_signal_22482 ), .Q ( new_AGEMA_signal_22483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C ( clk ), .D ( new_AGEMA_signal_22484 ), .Q ( new_AGEMA_signal_22485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C ( clk ), .D ( new_AGEMA_signal_22486 ), .Q ( new_AGEMA_signal_22487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C ( clk ), .D ( new_AGEMA_signal_22488 ), .Q ( new_AGEMA_signal_22489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C ( clk ), .D ( new_AGEMA_signal_22490 ), .Q ( new_AGEMA_signal_22491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C ( clk ), .D ( new_AGEMA_signal_22494 ), .Q ( new_AGEMA_signal_22495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C ( clk ), .D ( new_AGEMA_signal_22498 ), .Q ( new_AGEMA_signal_22499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C ( clk ), .D ( new_AGEMA_signal_22502 ), .Q ( new_AGEMA_signal_22503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C ( clk ), .D ( new_AGEMA_signal_22506 ), .Q ( new_AGEMA_signal_22507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C ( clk ), .D ( new_AGEMA_signal_22510 ), .Q ( new_AGEMA_signal_22511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C ( clk ), .D ( new_AGEMA_signal_22518 ), .Q ( new_AGEMA_signal_22519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C ( clk ), .D ( new_AGEMA_signal_22526 ), .Q ( new_AGEMA_signal_22527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C ( clk ), .D ( new_AGEMA_signal_22534 ), .Q ( new_AGEMA_signal_22535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C ( clk ), .D ( new_AGEMA_signal_22542 ), .Q ( new_AGEMA_signal_22543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C ( clk ), .D ( new_AGEMA_signal_22550 ), .Q ( new_AGEMA_signal_22551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C ( clk ), .D ( new_AGEMA_signal_22558 ), .Q ( new_AGEMA_signal_22559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C ( clk ), .D ( new_AGEMA_signal_22566 ), .Q ( new_AGEMA_signal_22567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C ( clk ), .D ( new_AGEMA_signal_22574 ), .Q ( new_AGEMA_signal_22575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C ( clk ), .D ( new_AGEMA_signal_22582 ), .Q ( new_AGEMA_signal_22583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C ( clk ), .D ( new_AGEMA_signal_22590 ), .Q ( new_AGEMA_signal_22591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C ( clk ), .D ( new_AGEMA_signal_22598 ), .Q ( new_AGEMA_signal_22599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C ( clk ), .D ( new_AGEMA_signal_22606 ), .Q ( new_AGEMA_signal_22607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C ( clk ), .D ( new_AGEMA_signal_22614 ), .Q ( new_AGEMA_signal_22615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C ( clk ), .D ( new_AGEMA_signal_22622 ), .Q ( new_AGEMA_signal_22623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C ( clk ), .D ( new_AGEMA_signal_22630 ), .Q ( new_AGEMA_signal_22631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C ( clk ), .D ( new_AGEMA_signal_22638 ), .Q ( new_AGEMA_signal_22639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C ( clk ), .D ( new_AGEMA_signal_22646 ), .Q ( new_AGEMA_signal_22647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C ( clk ), .D ( new_AGEMA_signal_22654 ), .Q ( new_AGEMA_signal_22655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C ( clk ), .D ( new_AGEMA_signal_22662 ), .Q ( new_AGEMA_signal_22663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C ( clk ), .D ( new_AGEMA_signal_22670 ), .Q ( new_AGEMA_signal_22671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C ( clk ), .D ( new_AGEMA_signal_22676 ), .Q ( new_AGEMA_signal_22677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C ( clk ), .D ( new_AGEMA_signal_22682 ), .Q ( new_AGEMA_signal_22683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C ( clk ), .D ( new_AGEMA_signal_22688 ), .Q ( new_AGEMA_signal_22689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C ( clk ), .D ( new_AGEMA_signal_22694 ), .Q ( new_AGEMA_signal_22695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C ( clk ), .D ( new_AGEMA_signal_22700 ), .Q ( new_AGEMA_signal_22701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C ( clk ), .D ( new_AGEMA_signal_22710 ), .Q ( new_AGEMA_signal_22711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C ( clk ), .D ( new_AGEMA_signal_22720 ), .Q ( new_AGEMA_signal_22721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C ( clk ), .D ( new_AGEMA_signal_22730 ), .Q ( new_AGEMA_signal_22731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C ( clk ), .D ( new_AGEMA_signal_22740 ), .Q ( new_AGEMA_signal_22741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C ( clk ), .D ( new_AGEMA_signal_22750 ), .Q ( new_AGEMA_signal_22751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C ( clk ), .D ( new_AGEMA_signal_22758 ), .Q ( new_AGEMA_signal_22759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C ( clk ), .D ( new_AGEMA_signal_22766 ), .Q ( new_AGEMA_signal_22767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C ( clk ), .D ( new_AGEMA_signal_22774 ), .Q ( new_AGEMA_signal_22775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C ( clk ), .D ( new_AGEMA_signal_22782 ), .Q ( new_AGEMA_signal_22783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C ( clk ), .D ( new_AGEMA_signal_22790 ), .Q ( new_AGEMA_signal_22791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C ( clk ), .D ( new_AGEMA_signal_22798 ), .Q ( new_AGEMA_signal_22799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C ( clk ), .D ( new_AGEMA_signal_22806 ), .Q ( new_AGEMA_signal_22807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C ( clk ), .D ( new_AGEMA_signal_22814 ), .Q ( new_AGEMA_signal_22815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C ( clk ), .D ( new_AGEMA_signal_22822 ), .Q ( new_AGEMA_signal_22823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C ( clk ), .D ( new_AGEMA_signal_22830 ), .Q ( new_AGEMA_signal_22831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C ( clk ), .D ( new_AGEMA_signal_22838 ), .Q ( new_AGEMA_signal_22839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C ( clk ), .D ( new_AGEMA_signal_22846 ), .Q ( new_AGEMA_signal_22847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C ( clk ), .D ( new_AGEMA_signal_22854 ), .Q ( new_AGEMA_signal_22855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C ( clk ), .D ( new_AGEMA_signal_22862 ), .Q ( new_AGEMA_signal_22863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C ( clk ), .D ( new_AGEMA_signal_22870 ), .Q ( new_AGEMA_signal_22871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C ( clk ), .D ( new_AGEMA_signal_22872 ), .Q ( new_AGEMA_signal_22873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C ( clk ), .D ( new_AGEMA_signal_22874 ), .Q ( new_AGEMA_signal_22875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C ( clk ), .D ( new_AGEMA_signal_22876 ), .Q ( new_AGEMA_signal_22877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C ( clk ), .D ( new_AGEMA_signal_22878 ), .Q ( new_AGEMA_signal_22879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C ( clk ), .D ( new_AGEMA_signal_22880 ), .Q ( new_AGEMA_signal_22881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C ( clk ), .D ( new_AGEMA_signal_22884 ), .Q ( new_AGEMA_signal_22885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C ( clk ), .D ( new_AGEMA_signal_22888 ), .Q ( new_AGEMA_signal_22889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C ( clk ), .D ( new_AGEMA_signal_22892 ), .Q ( new_AGEMA_signal_22893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C ( clk ), .D ( new_AGEMA_signal_22896 ), .Q ( new_AGEMA_signal_22897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C ( clk ), .D ( new_AGEMA_signal_22900 ), .Q ( new_AGEMA_signal_22901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C ( clk ), .D ( new_AGEMA_signal_22906 ), .Q ( new_AGEMA_signal_22907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C ( clk ), .D ( new_AGEMA_signal_22912 ), .Q ( new_AGEMA_signal_22913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C ( clk ), .D ( new_AGEMA_signal_22918 ), .Q ( new_AGEMA_signal_22919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C ( clk ), .D ( new_AGEMA_signal_22924 ), .Q ( new_AGEMA_signal_22925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C ( clk ), .D ( new_AGEMA_signal_22930 ), .Q ( new_AGEMA_signal_22931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C ( clk ), .D ( new_AGEMA_signal_22934 ), .Q ( new_AGEMA_signal_22935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C ( clk ), .D ( new_AGEMA_signal_22938 ), .Q ( new_AGEMA_signal_22939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C ( clk ), .D ( new_AGEMA_signal_22942 ), .Q ( new_AGEMA_signal_22943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C ( clk ), .D ( new_AGEMA_signal_22946 ), .Q ( new_AGEMA_signal_22947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C ( clk ), .D ( new_AGEMA_signal_22950 ), .Q ( new_AGEMA_signal_22951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C ( clk ), .D ( new_AGEMA_signal_22960 ), .Q ( new_AGEMA_signal_22961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C ( clk ), .D ( new_AGEMA_signal_22970 ), .Q ( new_AGEMA_signal_22971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C ( clk ), .D ( new_AGEMA_signal_22980 ), .Q ( new_AGEMA_signal_22981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C ( clk ), .D ( new_AGEMA_signal_22990 ), .Q ( new_AGEMA_signal_22991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C ( clk ), .D ( new_AGEMA_signal_23000 ), .Q ( new_AGEMA_signal_23001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C ( clk ), .D ( new_AGEMA_signal_23008 ), .Q ( new_AGEMA_signal_23009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C ( clk ), .D ( new_AGEMA_signal_23016 ), .Q ( new_AGEMA_signal_23017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C ( clk ), .D ( new_AGEMA_signal_23024 ), .Q ( new_AGEMA_signal_23025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C ( clk ), .D ( new_AGEMA_signal_23032 ), .Q ( new_AGEMA_signal_23033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C ( clk ), .D ( new_AGEMA_signal_23040 ), .Q ( new_AGEMA_signal_23041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C ( clk ), .D ( new_AGEMA_signal_23044 ), .Q ( new_AGEMA_signal_23045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C ( clk ), .D ( new_AGEMA_signal_23048 ), .Q ( new_AGEMA_signal_23049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C ( clk ), .D ( new_AGEMA_signal_23052 ), .Q ( new_AGEMA_signal_23053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C ( clk ), .D ( new_AGEMA_signal_23056 ), .Q ( new_AGEMA_signal_23057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C ( clk ), .D ( new_AGEMA_signal_23060 ), .Q ( new_AGEMA_signal_23061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C ( clk ), .D ( new_AGEMA_signal_23062 ), .Q ( new_AGEMA_signal_23063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C ( clk ), .D ( new_AGEMA_signal_23064 ), .Q ( new_AGEMA_signal_23065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C ( clk ), .D ( new_AGEMA_signal_23066 ), .Q ( new_AGEMA_signal_23067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C ( clk ), .D ( new_AGEMA_signal_23068 ), .Q ( new_AGEMA_signal_23069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C ( clk ), .D ( new_AGEMA_signal_23070 ), .Q ( new_AGEMA_signal_23071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C ( clk ), .D ( new_AGEMA_signal_23078 ), .Q ( new_AGEMA_signal_23079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C ( clk ), .D ( new_AGEMA_signal_23086 ), .Q ( new_AGEMA_signal_23087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C ( clk ), .D ( new_AGEMA_signal_23094 ), .Q ( new_AGEMA_signal_23095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C ( clk ), .D ( new_AGEMA_signal_23102 ), .Q ( new_AGEMA_signal_23103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C ( clk ), .D ( new_AGEMA_signal_23110 ), .Q ( new_AGEMA_signal_23111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C ( clk ), .D ( new_AGEMA_signal_23118 ), .Q ( new_AGEMA_signal_23119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C ( clk ), .D ( new_AGEMA_signal_23126 ), .Q ( new_AGEMA_signal_23127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C ( clk ), .D ( new_AGEMA_signal_23134 ), .Q ( new_AGEMA_signal_23135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C ( clk ), .D ( new_AGEMA_signal_23142 ), .Q ( new_AGEMA_signal_23143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C ( clk ), .D ( new_AGEMA_signal_23150 ), .Q ( new_AGEMA_signal_23151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C ( clk ), .D ( new_AGEMA_signal_23156 ), .Q ( new_AGEMA_signal_23157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C ( clk ), .D ( new_AGEMA_signal_23162 ), .Q ( new_AGEMA_signal_23163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C ( clk ), .D ( new_AGEMA_signal_23168 ), .Q ( new_AGEMA_signal_23169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C ( clk ), .D ( new_AGEMA_signal_23174 ), .Q ( new_AGEMA_signal_23175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C ( clk ), .D ( new_AGEMA_signal_23180 ), .Q ( new_AGEMA_signal_23181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C ( clk ), .D ( new_AGEMA_signal_23184 ), .Q ( new_AGEMA_signal_23185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C ( clk ), .D ( new_AGEMA_signal_23188 ), .Q ( new_AGEMA_signal_23189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C ( clk ), .D ( new_AGEMA_signal_23192 ), .Q ( new_AGEMA_signal_23193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C ( clk ), .D ( new_AGEMA_signal_23196 ), .Q ( new_AGEMA_signal_23197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C ( clk ), .D ( new_AGEMA_signal_23200 ), .Q ( new_AGEMA_signal_23201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C ( clk ), .D ( new_AGEMA_signal_23208 ), .Q ( new_AGEMA_signal_23209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C ( clk ), .D ( new_AGEMA_signal_23216 ), .Q ( new_AGEMA_signal_23217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C ( clk ), .D ( new_AGEMA_signal_23224 ), .Q ( new_AGEMA_signal_23225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C ( clk ), .D ( new_AGEMA_signal_23232 ), .Q ( new_AGEMA_signal_23233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C ( clk ), .D ( new_AGEMA_signal_23240 ), .Q ( new_AGEMA_signal_23241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C ( clk ), .D ( new_AGEMA_signal_23242 ), .Q ( new_AGEMA_signal_23243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C ( clk ), .D ( new_AGEMA_signal_23244 ), .Q ( new_AGEMA_signal_23245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C ( clk ), .D ( new_AGEMA_signal_23246 ), .Q ( new_AGEMA_signal_23247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C ( clk ), .D ( new_AGEMA_signal_23248 ), .Q ( new_AGEMA_signal_23249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C ( clk ), .D ( new_AGEMA_signal_23250 ), .Q ( new_AGEMA_signal_23251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C ( clk ), .D ( new_AGEMA_signal_23254 ), .Q ( new_AGEMA_signal_23255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C ( clk ), .D ( new_AGEMA_signal_23260 ), .Q ( new_AGEMA_signal_23261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C ( clk ), .D ( new_AGEMA_signal_23266 ), .Q ( new_AGEMA_signal_23267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C ( clk ), .D ( new_AGEMA_signal_23272 ), .Q ( new_AGEMA_signal_23273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C ( clk ), .D ( new_AGEMA_signal_23278 ), .Q ( new_AGEMA_signal_23279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C ( clk ), .D ( new_AGEMA_signal_23284 ), .Q ( new_AGEMA_signal_23285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C ( clk ), .D ( new_AGEMA_signal_23290 ), .Q ( new_AGEMA_signal_23291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C ( clk ), .D ( new_AGEMA_signal_23296 ), .Q ( new_AGEMA_signal_23297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C ( clk ), .D ( new_AGEMA_signal_23302 ), .Q ( new_AGEMA_signal_23303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C ( clk ), .D ( new_AGEMA_signal_23308 ), .Q ( new_AGEMA_signal_23309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C ( clk ), .D ( new_AGEMA_signal_23314 ), .Q ( new_AGEMA_signal_23315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C ( clk ), .D ( new_AGEMA_signal_23320 ), .Q ( new_AGEMA_signal_23321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C ( clk ), .D ( new_AGEMA_signal_23326 ), .Q ( new_AGEMA_signal_23327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C ( clk ), .D ( new_AGEMA_signal_23332 ), .Q ( new_AGEMA_signal_23333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C ( clk ), .D ( new_AGEMA_signal_23338 ), .Q ( new_AGEMA_signal_23339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C ( clk ), .D ( new_AGEMA_signal_23342 ), .Q ( new_AGEMA_signal_23343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C ( clk ), .D ( new_AGEMA_signal_23346 ), .Q ( new_AGEMA_signal_23347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C ( clk ), .D ( new_AGEMA_signal_23350 ), .Q ( new_AGEMA_signal_23351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C ( clk ), .D ( new_AGEMA_signal_23354 ), .Q ( new_AGEMA_signal_23355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C ( clk ), .D ( new_AGEMA_signal_23358 ), .Q ( new_AGEMA_signal_23359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C ( clk ), .D ( new_AGEMA_signal_23366 ), .Q ( new_AGEMA_signal_23367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C ( clk ), .D ( new_AGEMA_signal_23374 ), .Q ( new_AGEMA_signal_23375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C ( clk ), .D ( new_AGEMA_signal_23382 ), .Q ( new_AGEMA_signal_23383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C ( clk ), .D ( new_AGEMA_signal_23390 ), .Q ( new_AGEMA_signal_23391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C ( clk ), .D ( new_AGEMA_signal_23398 ), .Q ( new_AGEMA_signal_23399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C ( clk ), .D ( new_AGEMA_signal_23404 ), .Q ( new_AGEMA_signal_23405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C ( clk ), .D ( new_AGEMA_signal_23410 ), .Q ( new_AGEMA_signal_23411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C ( clk ), .D ( new_AGEMA_signal_23416 ), .Q ( new_AGEMA_signal_23417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C ( clk ), .D ( new_AGEMA_signal_23422 ), .Q ( new_AGEMA_signal_23423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C ( clk ), .D ( new_AGEMA_signal_23428 ), .Q ( new_AGEMA_signal_23429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C ( clk ), .D ( new_AGEMA_signal_23432 ), .Q ( new_AGEMA_signal_23433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C ( clk ), .D ( new_AGEMA_signal_23436 ), .Q ( new_AGEMA_signal_23437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C ( clk ), .D ( new_AGEMA_signal_23440 ), .Q ( new_AGEMA_signal_23441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C ( clk ), .D ( new_AGEMA_signal_23444 ), .Q ( new_AGEMA_signal_23445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C ( clk ), .D ( new_AGEMA_signal_23448 ), .Q ( new_AGEMA_signal_23449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C ( clk ), .D ( new_AGEMA_signal_23456 ), .Q ( new_AGEMA_signal_23457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C ( clk ), .D ( new_AGEMA_signal_23464 ), .Q ( new_AGEMA_signal_23465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C ( clk ), .D ( new_AGEMA_signal_23472 ), .Q ( new_AGEMA_signal_23473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C ( clk ), .D ( new_AGEMA_signal_23480 ), .Q ( new_AGEMA_signal_23481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C ( clk ), .D ( new_AGEMA_signal_23488 ), .Q ( new_AGEMA_signal_23489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C ( clk ), .D ( new_AGEMA_signal_23496 ), .Q ( new_AGEMA_signal_23497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C ( clk ), .D ( new_AGEMA_signal_23504 ), .Q ( new_AGEMA_signal_23505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C ( clk ), .D ( new_AGEMA_signal_23512 ), .Q ( new_AGEMA_signal_23513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C ( clk ), .D ( new_AGEMA_signal_23520 ), .Q ( new_AGEMA_signal_23521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C ( clk ), .D ( new_AGEMA_signal_23528 ), .Q ( new_AGEMA_signal_23529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C ( clk ), .D ( new_AGEMA_signal_23538 ), .Q ( new_AGEMA_signal_23539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C ( clk ), .D ( new_AGEMA_signal_23548 ), .Q ( new_AGEMA_signal_23549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C ( clk ), .D ( new_AGEMA_signal_23558 ), .Q ( new_AGEMA_signal_23559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C ( clk ), .D ( new_AGEMA_signal_23568 ), .Q ( new_AGEMA_signal_23569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C ( clk ), .D ( new_AGEMA_signal_23578 ), .Q ( new_AGEMA_signal_23579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C ( clk ), .D ( new_AGEMA_signal_23586 ), .Q ( new_AGEMA_signal_23587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C ( clk ), .D ( new_AGEMA_signal_23594 ), .Q ( new_AGEMA_signal_23595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C ( clk ), .D ( new_AGEMA_signal_23602 ), .Q ( new_AGEMA_signal_23603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C ( clk ), .D ( new_AGEMA_signal_23610 ), .Q ( new_AGEMA_signal_23611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C ( clk ), .D ( new_AGEMA_signal_23618 ), .Q ( new_AGEMA_signal_23619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C ( clk ), .D ( new_AGEMA_signal_23624 ), .Q ( new_AGEMA_signal_23625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C ( clk ), .D ( new_AGEMA_signal_23630 ), .Q ( new_AGEMA_signal_23631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C ( clk ), .D ( new_AGEMA_signal_23636 ), .Q ( new_AGEMA_signal_23637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C ( clk ), .D ( new_AGEMA_signal_23642 ), .Q ( new_AGEMA_signal_23643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C ( clk ), .D ( new_AGEMA_signal_23648 ), .Q ( new_AGEMA_signal_23649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C ( clk ), .D ( new_AGEMA_signal_23652 ), .Q ( new_AGEMA_signal_23653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C ( clk ), .D ( new_AGEMA_signal_23656 ), .Q ( new_AGEMA_signal_23657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C ( clk ), .D ( new_AGEMA_signal_23660 ), .Q ( new_AGEMA_signal_23661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C ( clk ), .D ( new_AGEMA_signal_23664 ), .Q ( new_AGEMA_signal_23665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C ( clk ), .D ( new_AGEMA_signal_23668 ), .Q ( new_AGEMA_signal_23669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C ( clk ), .D ( new_AGEMA_signal_23674 ), .Q ( new_AGEMA_signal_23675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C ( clk ), .D ( new_AGEMA_signal_23680 ), .Q ( new_AGEMA_signal_23681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C ( clk ), .D ( new_AGEMA_signal_23686 ), .Q ( new_AGEMA_signal_23687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C ( clk ), .D ( new_AGEMA_signal_23692 ), .Q ( new_AGEMA_signal_23693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C ( clk ), .D ( new_AGEMA_signal_23698 ), .Q ( new_AGEMA_signal_23699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C ( clk ), .D ( new_AGEMA_signal_23706 ), .Q ( new_AGEMA_signal_23707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C ( clk ), .D ( new_AGEMA_signal_23714 ), .Q ( new_AGEMA_signal_23715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C ( clk ), .D ( new_AGEMA_signal_23722 ), .Q ( new_AGEMA_signal_23723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C ( clk ), .D ( new_AGEMA_signal_23730 ), .Q ( new_AGEMA_signal_23731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C ( clk ), .D ( new_AGEMA_signal_23738 ), .Q ( new_AGEMA_signal_23739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C ( clk ), .D ( new_AGEMA_signal_23744 ), .Q ( new_AGEMA_signal_23745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C ( clk ), .D ( new_AGEMA_signal_23750 ), .Q ( new_AGEMA_signal_23751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C ( clk ), .D ( new_AGEMA_signal_23756 ), .Q ( new_AGEMA_signal_23757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C ( clk ), .D ( new_AGEMA_signal_23762 ), .Q ( new_AGEMA_signal_23763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C ( clk ), .D ( new_AGEMA_signal_23768 ), .Q ( new_AGEMA_signal_23769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C ( clk ), .D ( new_AGEMA_signal_23786 ), .Q ( new_AGEMA_signal_23787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C ( clk ), .D ( new_AGEMA_signal_23794 ), .Q ( new_AGEMA_signal_23795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C ( clk ), .D ( new_AGEMA_signal_23802 ), .Q ( new_AGEMA_signal_23803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C ( clk ), .D ( new_AGEMA_signal_23810 ), .Q ( new_AGEMA_signal_23811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C ( clk ), .D ( new_AGEMA_signal_23818 ), .Q ( new_AGEMA_signal_23819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C ( clk ), .D ( new_AGEMA_signal_23822 ), .Q ( new_AGEMA_signal_23823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C ( clk ), .D ( new_AGEMA_signal_23826 ), .Q ( new_AGEMA_signal_23827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C ( clk ), .D ( new_AGEMA_signal_23830 ), .Q ( new_AGEMA_signal_23831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C ( clk ), .D ( new_AGEMA_signal_23834 ), .Q ( new_AGEMA_signal_23835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C ( clk ), .D ( new_AGEMA_signal_23838 ), .Q ( new_AGEMA_signal_23839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C ( clk ), .D ( new_AGEMA_signal_23844 ), .Q ( new_AGEMA_signal_23845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C ( clk ), .D ( new_AGEMA_signal_23850 ), .Q ( new_AGEMA_signal_23851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C ( clk ), .D ( new_AGEMA_signal_23856 ), .Q ( new_AGEMA_signal_23857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C ( clk ), .D ( new_AGEMA_signal_23862 ), .Q ( new_AGEMA_signal_23863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C ( clk ), .D ( new_AGEMA_signal_23868 ), .Q ( new_AGEMA_signal_23869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C ( clk ), .D ( new_AGEMA_signal_23874 ), .Q ( new_AGEMA_signal_23875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C ( clk ), .D ( new_AGEMA_signal_23880 ), .Q ( new_AGEMA_signal_23881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C ( clk ), .D ( new_AGEMA_signal_23886 ), .Q ( new_AGEMA_signal_23887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C ( clk ), .D ( new_AGEMA_signal_23892 ), .Q ( new_AGEMA_signal_23893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C ( clk ), .D ( new_AGEMA_signal_23898 ), .Q ( new_AGEMA_signal_23899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C ( clk ), .D ( new_AGEMA_signal_23902 ), .Q ( new_AGEMA_signal_23903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C ( clk ), .D ( new_AGEMA_signal_23906 ), .Q ( new_AGEMA_signal_23907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C ( clk ), .D ( new_AGEMA_signal_23910 ), .Q ( new_AGEMA_signal_23911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C ( clk ), .D ( new_AGEMA_signal_23914 ), .Q ( new_AGEMA_signal_23915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C ( clk ), .D ( new_AGEMA_signal_23918 ), .Q ( new_AGEMA_signal_23919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C ( clk ), .D ( new_AGEMA_signal_23922 ), .Q ( new_AGEMA_signal_23923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C ( clk ), .D ( new_AGEMA_signal_23928 ), .Q ( new_AGEMA_signal_23929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C ( clk ), .D ( new_AGEMA_signal_23934 ), .Q ( new_AGEMA_signal_23935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C ( clk ), .D ( new_AGEMA_signal_23940 ), .Q ( new_AGEMA_signal_23941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C ( clk ), .D ( new_AGEMA_signal_23946 ), .Q ( new_AGEMA_signal_23947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C ( clk ), .D ( new_AGEMA_signal_23972 ), .Q ( new_AGEMA_signal_23973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C ( clk ), .D ( new_AGEMA_signal_23978 ), .Q ( new_AGEMA_signal_23979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C ( clk ), .D ( new_AGEMA_signal_23984 ), .Q ( new_AGEMA_signal_23985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C ( clk ), .D ( new_AGEMA_signal_23990 ), .Q ( new_AGEMA_signal_23991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C ( clk ), .D ( new_AGEMA_signal_23996 ), .Q ( new_AGEMA_signal_23997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C ( clk ), .D ( new_AGEMA_signal_24006 ), .Q ( new_AGEMA_signal_24007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C ( clk ), .D ( new_AGEMA_signal_24016 ), .Q ( new_AGEMA_signal_24017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C ( clk ), .D ( new_AGEMA_signal_24026 ), .Q ( new_AGEMA_signal_24027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C ( clk ), .D ( new_AGEMA_signal_24036 ), .Q ( new_AGEMA_signal_24037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C ( clk ), .D ( new_AGEMA_signal_24046 ), .Q ( new_AGEMA_signal_24047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C ( clk ), .D ( new_AGEMA_signal_24052 ), .Q ( new_AGEMA_signal_24053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C ( clk ), .D ( new_AGEMA_signal_24058 ), .Q ( new_AGEMA_signal_24059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C ( clk ), .D ( new_AGEMA_signal_24064 ), .Q ( new_AGEMA_signal_24065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C ( clk ), .D ( new_AGEMA_signal_24070 ), .Q ( new_AGEMA_signal_24071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C ( clk ), .D ( new_AGEMA_signal_24076 ), .Q ( new_AGEMA_signal_24077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C ( clk ), .D ( new_AGEMA_signal_24082 ), .Q ( new_AGEMA_signal_24083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C ( clk ), .D ( new_AGEMA_signal_24088 ), .Q ( new_AGEMA_signal_24089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C ( clk ), .D ( new_AGEMA_signal_24094 ), .Q ( new_AGEMA_signal_24095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C ( clk ), .D ( new_AGEMA_signal_24100 ), .Q ( new_AGEMA_signal_24101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C ( clk ), .D ( new_AGEMA_signal_24106 ), .Q ( new_AGEMA_signal_24107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C ( clk ), .D ( new_AGEMA_signal_24154 ), .Q ( new_AGEMA_signal_24155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C ( clk ), .D ( new_AGEMA_signal_24162 ), .Q ( new_AGEMA_signal_24163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C ( clk ), .D ( new_AGEMA_signal_24170 ), .Q ( new_AGEMA_signal_24171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C ( clk ), .D ( new_AGEMA_signal_24178 ), .Q ( new_AGEMA_signal_24179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C ( clk ), .D ( new_AGEMA_signal_24186 ), .Q ( new_AGEMA_signal_24187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C ( clk ), .D ( new_AGEMA_signal_24192 ), .Q ( new_AGEMA_signal_24193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C ( clk ), .D ( new_AGEMA_signal_24198 ), .Q ( new_AGEMA_signal_24199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C ( clk ), .D ( new_AGEMA_signal_24204 ), .Q ( new_AGEMA_signal_24205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C ( clk ), .D ( new_AGEMA_signal_24210 ), .Q ( new_AGEMA_signal_24211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C ( clk ), .D ( new_AGEMA_signal_24216 ), .Q ( new_AGEMA_signal_24217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C ( clk ), .D ( new_AGEMA_signal_24224 ), .Q ( new_AGEMA_signal_24225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C ( clk ), .D ( new_AGEMA_signal_24232 ), .Q ( new_AGEMA_signal_24233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C ( clk ), .D ( new_AGEMA_signal_24240 ), .Q ( new_AGEMA_signal_24241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C ( clk ), .D ( new_AGEMA_signal_24248 ), .Q ( new_AGEMA_signal_24249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C ( clk ), .D ( new_AGEMA_signal_24256 ), .Q ( new_AGEMA_signal_24257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C ( clk ), .D ( new_AGEMA_signal_24264 ), .Q ( new_AGEMA_signal_24265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C ( clk ), .D ( new_AGEMA_signal_24272 ), .Q ( new_AGEMA_signal_24273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C ( clk ), .D ( new_AGEMA_signal_24280 ), .Q ( new_AGEMA_signal_24281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C ( clk ), .D ( new_AGEMA_signal_24288 ), .Q ( new_AGEMA_signal_24289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C ( clk ), .D ( new_AGEMA_signal_24296 ), .Q ( new_AGEMA_signal_24297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C ( clk ), .D ( new_AGEMA_signal_24354 ), .Q ( new_AGEMA_signal_24355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C ( clk ), .D ( new_AGEMA_signal_24362 ), .Q ( new_AGEMA_signal_24363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C ( clk ), .D ( new_AGEMA_signal_24370 ), .Q ( new_AGEMA_signal_24371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C ( clk ), .D ( new_AGEMA_signal_24378 ), .Q ( new_AGEMA_signal_24379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C ( clk ), .D ( new_AGEMA_signal_24386 ), .Q ( new_AGEMA_signal_24387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C ( clk ), .D ( new_AGEMA_signal_24412 ), .Q ( new_AGEMA_signal_24413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C ( clk ), .D ( new_AGEMA_signal_24420 ), .Q ( new_AGEMA_signal_24421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C ( clk ), .D ( new_AGEMA_signal_24428 ), .Q ( new_AGEMA_signal_24429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C ( clk ), .D ( new_AGEMA_signal_24436 ), .Q ( new_AGEMA_signal_24437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7670 ( .C ( clk ), .D ( new_AGEMA_signal_24444 ), .Q ( new_AGEMA_signal_24445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7682 ( .C ( clk ), .D ( new_AGEMA_signal_24456 ), .Q ( new_AGEMA_signal_24457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7694 ( .C ( clk ), .D ( new_AGEMA_signal_24468 ), .Q ( new_AGEMA_signal_24469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7706 ( .C ( clk ), .D ( new_AGEMA_signal_24480 ), .Q ( new_AGEMA_signal_24481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7718 ( .C ( clk ), .D ( new_AGEMA_signal_24492 ), .Q ( new_AGEMA_signal_24493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7730 ( .C ( clk ), .D ( new_AGEMA_signal_24504 ), .Q ( new_AGEMA_signal_24505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7744 ( .C ( clk ), .D ( new_AGEMA_signal_24518 ), .Q ( new_AGEMA_signal_24519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7758 ( .C ( clk ), .D ( new_AGEMA_signal_24532 ), .Q ( new_AGEMA_signal_24533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7772 ( .C ( clk ), .D ( new_AGEMA_signal_24546 ), .Q ( new_AGEMA_signal_24547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7786 ( .C ( clk ), .D ( new_AGEMA_signal_24560 ), .Q ( new_AGEMA_signal_24561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7800 ( .C ( clk ), .D ( new_AGEMA_signal_24574 ), .Q ( new_AGEMA_signal_24575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7808 ( .C ( clk ), .D ( new_AGEMA_signal_24582 ), .Q ( new_AGEMA_signal_24583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7816 ( .C ( clk ), .D ( new_AGEMA_signal_24590 ), .Q ( new_AGEMA_signal_24591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7824 ( .C ( clk ), .D ( new_AGEMA_signal_24598 ), .Q ( new_AGEMA_signal_24599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7832 ( .C ( clk ), .D ( new_AGEMA_signal_24606 ), .Q ( new_AGEMA_signal_24607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7840 ( .C ( clk ), .D ( new_AGEMA_signal_24614 ), .Q ( new_AGEMA_signal_24615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7854 ( .C ( clk ), .D ( new_AGEMA_signal_24628 ), .Q ( new_AGEMA_signal_24629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7868 ( .C ( clk ), .D ( new_AGEMA_signal_24642 ), .Q ( new_AGEMA_signal_24643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7882 ( .C ( clk ), .D ( new_AGEMA_signal_24656 ), .Q ( new_AGEMA_signal_24657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7896 ( .C ( clk ), .D ( new_AGEMA_signal_24670 ), .Q ( new_AGEMA_signal_24671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7910 ( .C ( clk ), .D ( new_AGEMA_signal_24684 ), .Q ( new_AGEMA_signal_24685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7918 ( .C ( clk ), .D ( new_AGEMA_signal_24692 ), .Q ( new_AGEMA_signal_24693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7926 ( .C ( clk ), .D ( new_AGEMA_signal_24700 ), .Q ( new_AGEMA_signal_24701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7934 ( .C ( clk ), .D ( new_AGEMA_signal_24708 ), .Q ( new_AGEMA_signal_24709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7942 ( .C ( clk ), .D ( new_AGEMA_signal_24716 ), .Q ( new_AGEMA_signal_24717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7950 ( .C ( clk ), .D ( new_AGEMA_signal_24724 ), .Q ( new_AGEMA_signal_24725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7958 ( .C ( clk ), .D ( new_AGEMA_signal_24732 ), .Q ( new_AGEMA_signal_24733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7966 ( .C ( clk ), .D ( new_AGEMA_signal_24740 ), .Q ( new_AGEMA_signal_24741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7974 ( .C ( clk ), .D ( new_AGEMA_signal_24748 ), .Q ( new_AGEMA_signal_24749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7982 ( .C ( clk ), .D ( new_AGEMA_signal_24756 ), .Q ( new_AGEMA_signal_24757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7990 ( .C ( clk ), .D ( new_AGEMA_signal_24764 ), .Q ( new_AGEMA_signal_24765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8034 ( .C ( clk ), .D ( new_AGEMA_signal_24808 ), .Q ( new_AGEMA_signal_24809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8050 ( .C ( clk ), .D ( new_AGEMA_signal_24824 ), .Q ( new_AGEMA_signal_24825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8066 ( .C ( clk ), .D ( new_AGEMA_signal_24840 ), .Q ( new_AGEMA_signal_24841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8082 ( .C ( clk ), .D ( new_AGEMA_signal_24856 ), .Q ( new_AGEMA_signal_24857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8098 ( .C ( clk ), .D ( new_AGEMA_signal_24872 ), .Q ( new_AGEMA_signal_24873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8144 ( .C ( clk ), .D ( new_AGEMA_signal_24918 ), .Q ( new_AGEMA_signal_24919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8160 ( .C ( clk ), .D ( new_AGEMA_signal_24934 ), .Q ( new_AGEMA_signal_24935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8176 ( .C ( clk ), .D ( new_AGEMA_signal_24950 ), .Q ( new_AGEMA_signal_24951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8192 ( .C ( clk ), .D ( new_AGEMA_signal_24966 ), .Q ( new_AGEMA_signal_24967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8208 ( .C ( clk ), .D ( new_AGEMA_signal_24982 ), .Q ( new_AGEMA_signal_24983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8218 ( .C ( clk ), .D ( new_AGEMA_signal_24992 ), .Q ( new_AGEMA_signal_24993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8228 ( .C ( clk ), .D ( new_AGEMA_signal_25002 ), .Q ( new_AGEMA_signal_25003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8238 ( .C ( clk ), .D ( new_AGEMA_signal_25012 ), .Q ( new_AGEMA_signal_25013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8248 ( .C ( clk ), .D ( new_AGEMA_signal_25022 ), .Q ( new_AGEMA_signal_25023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8258 ( .C ( clk ), .D ( new_AGEMA_signal_25032 ), .Q ( new_AGEMA_signal_25033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8392 ( .C ( clk ), .D ( new_AGEMA_signal_25166 ), .Q ( new_AGEMA_signal_25167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8408 ( .C ( clk ), .D ( new_AGEMA_signal_25182 ), .Q ( new_AGEMA_signal_25183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8424 ( .C ( clk ), .D ( new_AGEMA_signal_25198 ), .Q ( new_AGEMA_signal_25199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8440 ( .C ( clk ), .D ( new_AGEMA_signal_25214 ), .Q ( new_AGEMA_signal_25215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8456 ( .C ( clk ), .D ( new_AGEMA_signal_25230 ), .Q ( new_AGEMA_signal_25231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8524 ( .C ( clk ), .D ( new_AGEMA_signal_25298 ), .Q ( new_AGEMA_signal_25299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8542 ( .C ( clk ), .D ( new_AGEMA_signal_25316 ), .Q ( new_AGEMA_signal_25317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8560 ( .C ( clk ), .D ( new_AGEMA_signal_25334 ), .Q ( new_AGEMA_signal_25335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8578 ( .C ( clk ), .D ( new_AGEMA_signal_25352 ), .Q ( new_AGEMA_signal_25353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8596 ( .C ( clk ), .D ( new_AGEMA_signal_25370 ), .Q ( new_AGEMA_signal_25371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8774 ( .C ( clk ), .D ( new_AGEMA_signal_25548 ), .Q ( new_AGEMA_signal_25549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8794 ( .C ( clk ), .D ( new_AGEMA_signal_25568 ), .Q ( new_AGEMA_signal_25569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8814 ( .C ( clk ), .D ( new_AGEMA_signal_25588 ), .Q ( new_AGEMA_signal_25589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8834 ( .C ( clk ), .D ( new_AGEMA_signal_25608 ), .Q ( new_AGEMA_signal_25609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8854 ( .C ( clk ), .D ( new_AGEMA_signal_25628 ), .Q ( new_AGEMA_signal_25629 ) ) ;

    /* cells in depth 15 */
    buf_clk new_AGEMA_reg_buffer_6481 ( .C ( clk ), .D ( new_AGEMA_signal_23255 ), .Q ( new_AGEMA_signal_23256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C ( clk ), .D ( new_AGEMA_signal_23261 ), .Q ( new_AGEMA_signal_23262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C ( clk ), .D ( new_AGEMA_signal_23267 ), .Q ( new_AGEMA_signal_23268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C ( clk ), .D ( new_AGEMA_signal_23273 ), .Q ( new_AGEMA_signal_23274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C ( clk ), .D ( new_AGEMA_signal_23279 ), .Q ( new_AGEMA_signal_23280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C ( clk ), .D ( new_AGEMA_signal_23285 ), .Q ( new_AGEMA_signal_23286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C ( clk ), .D ( new_AGEMA_signal_23291 ), .Q ( new_AGEMA_signal_23292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C ( clk ), .D ( new_AGEMA_signal_23297 ), .Q ( new_AGEMA_signal_23298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C ( clk ), .D ( new_AGEMA_signal_23303 ), .Q ( new_AGEMA_signal_23304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C ( clk ), .D ( new_AGEMA_signal_23309 ), .Q ( new_AGEMA_signal_23310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C ( clk ), .D ( new_AGEMA_signal_23315 ), .Q ( new_AGEMA_signal_23316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C ( clk ), .D ( new_AGEMA_signal_23321 ), .Q ( new_AGEMA_signal_23322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C ( clk ), .D ( new_AGEMA_signal_23327 ), .Q ( new_AGEMA_signal_23328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C ( clk ), .D ( new_AGEMA_signal_23333 ), .Q ( new_AGEMA_signal_23334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C ( clk ), .D ( new_AGEMA_signal_23339 ), .Q ( new_AGEMA_signal_23340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C ( clk ), .D ( new_AGEMA_signal_23343 ), .Q ( new_AGEMA_signal_23344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C ( clk ), .D ( new_AGEMA_signal_23347 ), .Q ( new_AGEMA_signal_23348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C ( clk ), .D ( new_AGEMA_signal_23351 ), .Q ( new_AGEMA_signal_23352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C ( clk ), .D ( new_AGEMA_signal_23355 ), .Q ( new_AGEMA_signal_23356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6585 ( .C ( clk ), .D ( new_AGEMA_signal_23359 ), .Q ( new_AGEMA_signal_23360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C ( clk ), .D ( new_AGEMA_signal_23367 ), .Q ( new_AGEMA_signal_23368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C ( clk ), .D ( new_AGEMA_signal_23375 ), .Q ( new_AGEMA_signal_23376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C ( clk ), .D ( new_AGEMA_signal_23383 ), .Q ( new_AGEMA_signal_23384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C ( clk ), .D ( new_AGEMA_signal_23391 ), .Q ( new_AGEMA_signal_23392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C ( clk ), .D ( new_AGEMA_signal_23399 ), .Q ( new_AGEMA_signal_23400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C ( clk ), .D ( new_AGEMA_signal_23405 ), .Q ( new_AGEMA_signal_23406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C ( clk ), .D ( new_AGEMA_signal_23411 ), .Q ( new_AGEMA_signal_23412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C ( clk ), .D ( new_AGEMA_signal_23417 ), .Q ( new_AGEMA_signal_23418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C ( clk ), .D ( new_AGEMA_signal_23423 ), .Q ( new_AGEMA_signal_23424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C ( clk ), .D ( new_AGEMA_signal_23429 ), .Q ( new_AGEMA_signal_23430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C ( clk ), .D ( new_AGEMA_signal_23433 ), .Q ( new_AGEMA_signal_23434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C ( clk ), .D ( new_AGEMA_signal_23437 ), .Q ( new_AGEMA_signal_23438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C ( clk ), .D ( new_AGEMA_signal_23441 ), .Q ( new_AGEMA_signal_23442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C ( clk ), .D ( new_AGEMA_signal_23445 ), .Q ( new_AGEMA_signal_23446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C ( clk ), .D ( new_AGEMA_signal_23449 ), .Q ( new_AGEMA_signal_23450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C ( clk ), .D ( new_AGEMA_signal_23457 ), .Q ( new_AGEMA_signal_23458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C ( clk ), .D ( new_AGEMA_signal_23465 ), .Q ( new_AGEMA_signal_23466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C ( clk ), .D ( new_AGEMA_signal_23473 ), .Q ( new_AGEMA_signal_23474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C ( clk ), .D ( new_AGEMA_signal_23481 ), .Q ( new_AGEMA_signal_23482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C ( clk ), .D ( new_AGEMA_signal_23489 ), .Q ( new_AGEMA_signal_23490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C ( clk ), .D ( new_AGEMA_signal_23497 ), .Q ( new_AGEMA_signal_23498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C ( clk ), .D ( new_AGEMA_signal_23505 ), .Q ( new_AGEMA_signal_23506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C ( clk ), .D ( new_AGEMA_signal_23513 ), .Q ( new_AGEMA_signal_23514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C ( clk ), .D ( new_AGEMA_signal_23521 ), .Q ( new_AGEMA_signal_23522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C ( clk ), .D ( new_AGEMA_signal_23529 ), .Q ( new_AGEMA_signal_23530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C ( clk ), .D ( new_AGEMA_signal_23539 ), .Q ( new_AGEMA_signal_23540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C ( clk ), .D ( new_AGEMA_signal_23549 ), .Q ( new_AGEMA_signal_23550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C ( clk ), .D ( new_AGEMA_signal_23559 ), .Q ( new_AGEMA_signal_23560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C ( clk ), .D ( new_AGEMA_signal_23569 ), .Q ( new_AGEMA_signal_23570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C ( clk ), .D ( new_AGEMA_signal_23579 ), .Q ( new_AGEMA_signal_23580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C ( clk ), .D ( new_AGEMA_signal_23587 ), .Q ( new_AGEMA_signal_23588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C ( clk ), .D ( new_AGEMA_signal_23595 ), .Q ( new_AGEMA_signal_23596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C ( clk ), .D ( new_AGEMA_signal_23603 ), .Q ( new_AGEMA_signal_23604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C ( clk ), .D ( new_AGEMA_signal_23611 ), .Q ( new_AGEMA_signal_23612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C ( clk ), .D ( new_AGEMA_signal_23619 ), .Q ( new_AGEMA_signal_23620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6851 ( .C ( clk ), .D ( new_AGEMA_signal_23625 ), .Q ( new_AGEMA_signal_23626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C ( clk ), .D ( new_AGEMA_signal_23631 ), .Q ( new_AGEMA_signal_23632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C ( clk ), .D ( new_AGEMA_signal_23637 ), .Q ( new_AGEMA_signal_23638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C ( clk ), .D ( new_AGEMA_signal_23643 ), .Q ( new_AGEMA_signal_23644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C ( clk ), .D ( new_AGEMA_signal_23649 ), .Q ( new_AGEMA_signal_23650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C ( clk ), .D ( new_AGEMA_signal_23653 ), .Q ( new_AGEMA_signal_23654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C ( clk ), .D ( new_AGEMA_signal_23657 ), .Q ( new_AGEMA_signal_23658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C ( clk ), .D ( new_AGEMA_signal_23661 ), .Q ( new_AGEMA_signal_23662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C ( clk ), .D ( new_AGEMA_signal_23665 ), .Q ( new_AGEMA_signal_23666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C ( clk ), .D ( new_AGEMA_signal_23669 ), .Q ( new_AGEMA_signal_23670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C ( clk ), .D ( new_AGEMA_signal_23675 ), .Q ( new_AGEMA_signal_23676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C ( clk ), .D ( new_AGEMA_signal_23681 ), .Q ( new_AGEMA_signal_23682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C ( clk ), .D ( new_AGEMA_signal_23687 ), .Q ( new_AGEMA_signal_23688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C ( clk ), .D ( new_AGEMA_signal_23693 ), .Q ( new_AGEMA_signal_23694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C ( clk ), .D ( new_AGEMA_signal_23699 ), .Q ( new_AGEMA_signal_23700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C ( clk ), .D ( new_AGEMA_signal_23707 ), .Q ( new_AGEMA_signal_23708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C ( clk ), .D ( new_AGEMA_signal_23715 ), .Q ( new_AGEMA_signal_23716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C ( clk ), .D ( new_AGEMA_signal_23723 ), .Q ( new_AGEMA_signal_23724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C ( clk ), .D ( new_AGEMA_signal_23731 ), .Q ( new_AGEMA_signal_23732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C ( clk ), .D ( new_AGEMA_signal_23739 ), .Q ( new_AGEMA_signal_23740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C ( clk ), .D ( new_AGEMA_signal_23745 ), .Q ( new_AGEMA_signal_23746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C ( clk ), .D ( new_AGEMA_signal_23751 ), .Q ( new_AGEMA_signal_23752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C ( clk ), .D ( new_AGEMA_signal_23757 ), .Q ( new_AGEMA_signal_23758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C ( clk ), .D ( new_AGEMA_signal_23763 ), .Q ( new_AGEMA_signal_23764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C ( clk ), .D ( new_AGEMA_signal_23769 ), .Q ( new_AGEMA_signal_23770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_23772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C ( clk ), .D ( new_AGEMA_signal_4194 ), .Q ( new_AGEMA_signal_23774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C ( clk ), .D ( new_AGEMA_signal_4195 ), .Q ( new_AGEMA_signal_23776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C ( clk ), .D ( new_AGEMA_signal_4196 ), .Q ( new_AGEMA_signal_23778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C ( clk ), .D ( new_AGEMA_signal_4197 ), .Q ( new_AGEMA_signal_23780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C ( clk ), .D ( new_AGEMA_signal_23787 ), .Q ( new_AGEMA_signal_23788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C ( clk ), .D ( new_AGEMA_signal_23795 ), .Q ( new_AGEMA_signal_23796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C ( clk ), .D ( new_AGEMA_signal_23803 ), .Q ( new_AGEMA_signal_23804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C ( clk ), .D ( new_AGEMA_signal_23811 ), .Q ( new_AGEMA_signal_23812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C ( clk ), .D ( new_AGEMA_signal_23819 ), .Q ( new_AGEMA_signal_23820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C ( clk ), .D ( new_AGEMA_signal_23823 ), .Q ( new_AGEMA_signal_23824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C ( clk ), .D ( new_AGEMA_signal_23827 ), .Q ( new_AGEMA_signal_23828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C ( clk ), .D ( new_AGEMA_signal_23831 ), .Q ( new_AGEMA_signal_23832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C ( clk ), .D ( new_AGEMA_signal_23835 ), .Q ( new_AGEMA_signal_23836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C ( clk ), .D ( new_AGEMA_signal_23839 ), .Q ( new_AGEMA_signal_23840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C ( clk ), .D ( new_AGEMA_signal_23845 ), .Q ( new_AGEMA_signal_23846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C ( clk ), .D ( new_AGEMA_signal_23851 ), .Q ( new_AGEMA_signal_23852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C ( clk ), .D ( new_AGEMA_signal_23857 ), .Q ( new_AGEMA_signal_23858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C ( clk ), .D ( new_AGEMA_signal_23863 ), .Q ( new_AGEMA_signal_23864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C ( clk ), .D ( new_AGEMA_signal_23869 ), .Q ( new_AGEMA_signal_23870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C ( clk ), .D ( new_AGEMA_signal_23875 ), .Q ( new_AGEMA_signal_23876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C ( clk ), .D ( new_AGEMA_signal_23881 ), .Q ( new_AGEMA_signal_23882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C ( clk ), .D ( new_AGEMA_signal_23887 ), .Q ( new_AGEMA_signal_23888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C ( clk ), .D ( new_AGEMA_signal_23893 ), .Q ( new_AGEMA_signal_23894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C ( clk ), .D ( new_AGEMA_signal_23899 ), .Q ( new_AGEMA_signal_23900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C ( clk ), .D ( new_AGEMA_signal_23903 ), .Q ( new_AGEMA_signal_23904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C ( clk ), .D ( new_AGEMA_signal_23907 ), .Q ( new_AGEMA_signal_23908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C ( clk ), .D ( new_AGEMA_signal_23911 ), .Q ( new_AGEMA_signal_23912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7141 ( .C ( clk ), .D ( new_AGEMA_signal_23915 ), .Q ( new_AGEMA_signal_23916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C ( clk ), .D ( new_AGEMA_signal_23919 ), .Q ( new_AGEMA_signal_23920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C ( clk ), .D ( new_AGEMA_signal_23923 ), .Q ( new_AGEMA_signal_23924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C ( clk ), .D ( new_AGEMA_signal_23929 ), .Q ( new_AGEMA_signal_23930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C ( clk ), .D ( new_AGEMA_signal_23935 ), .Q ( new_AGEMA_signal_23936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C ( clk ), .D ( new_AGEMA_signal_23941 ), .Q ( new_AGEMA_signal_23942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C ( clk ), .D ( new_AGEMA_signal_23947 ), .Q ( new_AGEMA_signal_23948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_23952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C ( clk ), .D ( new_AGEMA_signal_4098 ), .Q ( new_AGEMA_signal_23956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C ( clk ), .D ( new_AGEMA_signal_4099 ), .Q ( new_AGEMA_signal_23960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C ( clk ), .D ( new_AGEMA_signal_4100 ), .Q ( new_AGEMA_signal_23964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C ( clk ), .D ( new_AGEMA_signal_4101 ), .Q ( new_AGEMA_signal_23968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C ( clk ), .D ( new_AGEMA_signal_23973 ), .Q ( new_AGEMA_signal_23974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C ( clk ), .D ( new_AGEMA_signal_23979 ), .Q ( new_AGEMA_signal_23980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C ( clk ), .D ( new_AGEMA_signal_23985 ), .Q ( new_AGEMA_signal_23986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C ( clk ), .D ( new_AGEMA_signal_23991 ), .Q ( new_AGEMA_signal_23992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C ( clk ), .D ( new_AGEMA_signal_23997 ), .Q ( new_AGEMA_signal_23998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C ( clk ), .D ( new_AGEMA_signal_24007 ), .Q ( new_AGEMA_signal_24008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C ( clk ), .D ( new_AGEMA_signal_24017 ), .Q ( new_AGEMA_signal_24018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C ( clk ), .D ( new_AGEMA_signal_24027 ), .Q ( new_AGEMA_signal_24028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C ( clk ), .D ( new_AGEMA_signal_24037 ), .Q ( new_AGEMA_signal_24038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C ( clk ), .D ( new_AGEMA_signal_24047 ), .Q ( new_AGEMA_signal_24048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C ( clk ), .D ( new_AGEMA_signal_24053 ), .Q ( new_AGEMA_signal_24054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7285 ( .C ( clk ), .D ( new_AGEMA_signal_24059 ), .Q ( new_AGEMA_signal_24060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C ( clk ), .D ( new_AGEMA_signal_24065 ), .Q ( new_AGEMA_signal_24066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C ( clk ), .D ( new_AGEMA_signal_24071 ), .Q ( new_AGEMA_signal_24072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C ( clk ), .D ( new_AGEMA_signal_24077 ), .Q ( new_AGEMA_signal_24078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C ( clk ), .D ( new_AGEMA_signal_24083 ), .Q ( new_AGEMA_signal_24084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C ( clk ), .D ( new_AGEMA_signal_24089 ), .Q ( new_AGEMA_signal_24090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C ( clk ), .D ( new_AGEMA_signal_24095 ), .Q ( new_AGEMA_signal_24096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C ( clk ), .D ( new_AGEMA_signal_24101 ), .Q ( new_AGEMA_signal_24102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C ( clk ), .D ( new_AGEMA_signal_24107 ), .Q ( new_AGEMA_signal_24108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_24112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C ( clk ), .D ( new_AGEMA_signal_4134 ), .Q ( new_AGEMA_signal_24116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C ( clk ), .D ( new_AGEMA_signal_4135 ), .Q ( new_AGEMA_signal_24120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C ( clk ), .D ( new_AGEMA_signal_4136 ), .Q ( new_AGEMA_signal_24124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C ( clk ), .D ( new_AGEMA_signal_4137 ), .Q ( new_AGEMA_signal_24128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_24132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C ( clk ), .D ( new_AGEMA_signal_4298 ), .Q ( new_AGEMA_signal_24136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C ( clk ), .D ( new_AGEMA_signal_4299 ), .Q ( new_AGEMA_signal_24140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C ( clk ), .D ( new_AGEMA_signal_4300 ), .Q ( new_AGEMA_signal_24144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C ( clk ), .D ( new_AGEMA_signal_4301 ), .Q ( new_AGEMA_signal_24148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C ( clk ), .D ( new_AGEMA_signal_24155 ), .Q ( new_AGEMA_signal_24156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C ( clk ), .D ( new_AGEMA_signal_24163 ), .Q ( new_AGEMA_signal_24164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C ( clk ), .D ( new_AGEMA_signal_24171 ), .Q ( new_AGEMA_signal_24172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C ( clk ), .D ( new_AGEMA_signal_24179 ), .Q ( new_AGEMA_signal_24180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C ( clk ), .D ( new_AGEMA_signal_24187 ), .Q ( new_AGEMA_signal_24188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C ( clk ), .D ( new_AGEMA_signal_24193 ), .Q ( new_AGEMA_signal_24194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C ( clk ), .D ( new_AGEMA_signal_24199 ), .Q ( new_AGEMA_signal_24200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C ( clk ), .D ( new_AGEMA_signal_24205 ), .Q ( new_AGEMA_signal_24206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C ( clk ), .D ( new_AGEMA_signal_24211 ), .Q ( new_AGEMA_signal_24212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C ( clk ), .D ( new_AGEMA_signal_24217 ), .Q ( new_AGEMA_signal_24218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C ( clk ), .D ( new_AGEMA_signal_24225 ), .Q ( new_AGEMA_signal_24226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C ( clk ), .D ( new_AGEMA_signal_24233 ), .Q ( new_AGEMA_signal_24234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C ( clk ), .D ( new_AGEMA_signal_24241 ), .Q ( new_AGEMA_signal_24242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7475 ( .C ( clk ), .D ( new_AGEMA_signal_24249 ), .Q ( new_AGEMA_signal_24250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C ( clk ), .D ( new_AGEMA_signal_24257 ), .Q ( new_AGEMA_signal_24258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C ( clk ), .D ( new_AGEMA_signal_24265 ), .Q ( new_AGEMA_signal_24266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C ( clk ), .D ( new_AGEMA_signal_24273 ), .Q ( new_AGEMA_signal_24274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C ( clk ), .D ( new_AGEMA_signal_24281 ), .Q ( new_AGEMA_signal_24282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C ( clk ), .D ( new_AGEMA_signal_24289 ), .Q ( new_AGEMA_signal_24290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C ( clk ), .D ( new_AGEMA_signal_24297 ), .Q ( new_AGEMA_signal_24298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_24312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C ( clk ), .D ( new_AGEMA_signal_4214 ), .Q ( new_AGEMA_signal_24316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C ( clk ), .D ( new_AGEMA_signal_4215 ), .Q ( new_AGEMA_signal_24320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C ( clk ), .D ( new_AGEMA_signal_4216 ), .Q ( new_AGEMA_signal_24324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C ( clk ), .D ( new_AGEMA_signal_4217 ), .Q ( new_AGEMA_signal_24328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_24332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C ( clk ), .D ( new_AGEMA_signal_4226 ), .Q ( new_AGEMA_signal_24336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C ( clk ), .D ( new_AGEMA_signal_4227 ), .Q ( new_AGEMA_signal_24340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C ( clk ), .D ( new_AGEMA_signal_4228 ), .Q ( new_AGEMA_signal_24344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C ( clk ), .D ( new_AGEMA_signal_4229 ), .Q ( new_AGEMA_signal_24348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C ( clk ), .D ( new_AGEMA_signal_24355 ), .Q ( new_AGEMA_signal_24356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C ( clk ), .D ( new_AGEMA_signal_24363 ), .Q ( new_AGEMA_signal_24364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C ( clk ), .D ( new_AGEMA_signal_24371 ), .Q ( new_AGEMA_signal_24372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C ( clk ), .D ( new_AGEMA_signal_24379 ), .Q ( new_AGEMA_signal_24380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C ( clk ), .D ( new_AGEMA_signal_24387 ), .Q ( new_AGEMA_signal_24388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_24392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C ( clk ), .D ( new_AGEMA_signal_4238 ), .Q ( new_AGEMA_signal_24396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C ( clk ), .D ( new_AGEMA_signal_4239 ), .Q ( new_AGEMA_signal_24400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C ( clk ), .D ( new_AGEMA_signal_4240 ), .Q ( new_AGEMA_signal_24404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C ( clk ), .D ( new_AGEMA_signal_4241 ), .Q ( new_AGEMA_signal_24408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C ( clk ), .D ( new_AGEMA_signal_24413 ), .Q ( new_AGEMA_signal_24414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C ( clk ), .D ( new_AGEMA_signal_24421 ), .Q ( new_AGEMA_signal_24422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C ( clk ), .D ( new_AGEMA_signal_24429 ), .Q ( new_AGEMA_signal_24430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7663 ( .C ( clk ), .D ( new_AGEMA_signal_24437 ), .Q ( new_AGEMA_signal_24438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7671 ( .C ( clk ), .D ( new_AGEMA_signal_24445 ), .Q ( new_AGEMA_signal_24446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7683 ( .C ( clk ), .D ( new_AGEMA_signal_24457 ), .Q ( new_AGEMA_signal_24458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7695 ( .C ( clk ), .D ( new_AGEMA_signal_24469 ), .Q ( new_AGEMA_signal_24470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7707 ( .C ( clk ), .D ( new_AGEMA_signal_24481 ), .Q ( new_AGEMA_signal_24482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7719 ( .C ( clk ), .D ( new_AGEMA_signal_24493 ), .Q ( new_AGEMA_signal_24494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7731 ( .C ( clk ), .D ( new_AGEMA_signal_24505 ), .Q ( new_AGEMA_signal_24506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7745 ( .C ( clk ), .D ( new_AGEMA_signal_24519 ), .Q ( new_AGEMA_signal_24520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7759 ( .C ( clk ), .D ( new_AGEMA_signal_24533 ), .Q ( new_AGEMA_signal_24534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7773 ( .C ( clk ), .D ( new_AGEMA_signal_24547 ), .Q ( new_AGEMA_signal_24548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7787 ( .C ( clk ), .D ( new_AGEMA_signal_24561 ), .Q ( new_AGEMA_signal_24562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7801 ( .C ( clk ), .D ( new_AGEMA_signal_24575 ), .Q ( new_AGEMA_signal_24576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7809 ( .C ( clk ), .D ( new_AGEMA_signal_24583 ), .Q ( new_AGEMA_signal_24584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7817 ( .C ( clk ), .D ( new_AGEMA_signal_24591 ), .Q ( new_AGEMA_signal_24592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7825 ( .C ( clk ), .D ( new_AGEMA_signal_24599 ), .Q ( new_AGEMA_signal_24600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7833 ( .C ( clk ), .D ( new_AGEMA_signal_24607 ), .Q ( new_AGEMA_signal_24608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7841 ( .C ( clk ), .D ( new_AGEMA_signal_24615 ), .Q ( new_AGEMA_signal_24616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7855 ( .C ( clk ), .D ( new_AGEMA_signal_24629 ), .Q ( new_AGEMA_signal_24630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7869 ( .C ( clk ), .D ( new_AGEMA_signal_24643 ), .Q ( new_AGEMA_signal_24644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7883 ( .C ( clk ), .D ( new_AGEMA_signal_24657 ), .Q ( new_AGEMA_signal_24658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7897 ( .C ( clk ), .D ( new_AGEMA_signal_24671 ), .Q ( new_AGEMA_signal_24672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7911 ( .C ( clk ), .D ( new_AGEMA_signal_24685 ), .Q ( new_AGEMA_signal_24686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7919 ( .C ( clk ), .D ( new_AGEMA_signal_24693 ), .Q ( new_AGEMA_signal_24694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7927 ( .C ( clk ), .D ( new_AGEMA_signal_24701 ), .Q ( new_AGEMA_signal_24702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7935 ( .C ( clk ), .D ( new_AGEMA_signal_24709 ), .Q ( new_AGEMA_signal_24710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7943 ( .C ( clk ), .D ( new_AGEMA_signal_24717 ), .Q ( new_AGEMA_signal_24718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7951 ( .C ( clk ), .D ( new_AGEMA_signal_24725 ), .Q ( new_AGEMA_signal_24726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7959 ( .C ( clk ), .D ( new_AGEMA_signal_24733 ), .Q ( new_AGEMA_signal_24734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7967 ( .C ( clk ), .D ( new_AGEMA_signal_24741 ), .Q ( new_AGEMA_signal_24742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7975 ( .C ( clk ), .D ( new_AGEMA_signal_24749 ), .Q ( new_AGEMA_signal_24750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7983 ( .C ( clk ), .D ( new_AGEMA_signal_24757 ), .Q ( new_AGEMA_signal_24758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7991 ( .C ( clk ), .D ( new_AGEMA_signal_24765 ), .Q ( new_AGEMA_signal_24766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8035 ( .C ( clk ), .D ( new_AGEMA_signal_24809 ), .Q ( new_AGEMA_signal_24810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8051 ( .C ( clk ), .D ( new_AGEMA_signal_24825 ), .Q ( new_AGEMA_signal_24826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8067 ( .C ( clk ), .D ( new_AGEMA_signal_24841 ), .Q ( new_AGEMA_signal_24842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8083 ( .C ( clk ), .D ( new_AGEMA_signal_24857 ), .Q ( new_AGEMA_signal_24858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8099 ( .C ( clk ), .D ( new_AGEMA_signal_24873 ), .Q ( new_AGEMA_signal_24874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8145 ( .C ( clk ), .D ( new_AGEMA_signal_24919 ), .Q ( new_AGEMA_signal_24920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8161 ( .C ( clk ), .D ( new_AGEMA_signal_24935 ), .Q ( new_AGEMA_signal_24936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8177 ( .C ( clk ), .D ( new_AGEMA_signal_24951 ), .Q ( new_AGEMA_signal_24952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8193 ( .C ( clk ), .D ( new_AGEMA_signal_24967 ), .Q ( new_AGEMA_signal_24968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8209 ( .C ( clk ), .D ( new_AGEMA_signal_24983 ), .Q ( new_AGEMA_signal_24984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8219 ( .C ( clk ), .D ( new_AGEMA_signal_24993 ), .Q ( new_AGEMA_signal_24994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8229 ( .C ( clk ), .D ( new_AGEMA_signal_25003 ), .Q ( new_AGEMA_signal_25004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8239 ( .C ( clk ), .D ( new_AGEMA_signal_25013 ), .Q ( new_AGEMA_signal_25014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8249 ( .C ( clk ), .D ( new_AGEMA_signal_25023 ), .Q ( new_AGEMA_signal_25024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8259 ( .C ( clk ), .D ( new_AGEMA_signal_25033 ), .Q ( new_AGEMA_signal_25034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8287 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_25062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8295 ( .C ( clk ), .D ( new_AGEMA_signal_4246 ), .Q ( new_AGEMA_signal_25070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8303 ( .C ( clk ), .D ( new_AGEMA_signal_4247 ), .Q ( new_AGEMA_signal_25078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8311 ( .C ( clk ), .D ( new_AGEMA_signal_4248 ), .Q ( new_AGEMA_signal_25086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8319 ( .C ( clk ), .D ( new_AGEMA_signal_4249 ), .Q ( new_AGEMA_signal_25094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8393 ( .C ( clk ), .D ( new_AGEMA_signal_25167 ), .Q ( new_AGEMA_signal_25168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8409 ( .C ( clk ), .D ( new_AGEMA_signal_25183 ), .Q ( new_AGEMA_signal_25184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8425 ( .C ( clk ), .D ( new_AGEMA_signal_25199 ), .Q ( new_AGEMA_signal_25200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8441 ( .C ( clk ), .D ( new_AGEMA_signal_25215 ), .Q ( new_AGEMA_signal_25216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8457 ( .C ( clk ), .D ( new_AGEMA_signal_25231 ), .Q ( new_AGEMA_signal_25232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8467 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_25242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8477 ( .C ( clk ), .D ( new_AGEMA_signal_4142 ), .Q ( new_AGEMA_signal_25252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8487 ( .C ( clk ), .D ( new_AGEMA_signal_4143 ), .Q ( new_AGEMA_signal_25262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8497 ( .C ( clk ), .D ( new_AGEMA_signal_4144 ), .Q ( new_AGEMA_signal_25272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8507 ( .C ( clk ), .D ( new_AGEMA_signal_4145 ), .Q ( new_AGEMA_signal_25282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8525 ( .C ( clk ), .D ( new_AGEMA_signal_25299 ), .Q ( new_AGEMA_signal_25300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8543 ( .C ( clk ), .D ( new_AGEMA_signal_25317 ), .Q ( new_AGEMA_signal_25318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8561 ( .C ( clk ), .D ( new_AGEMA_signal_25335 ), .Q ( new_AGEMA_signal_25336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8579 ( .C ( clk ), .D ( new_AGEMA_signal_25353 ), .Q ( new_AGEMA_signal_25354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8597 ( .C ( clk ), .D ( new_AGEMA_signal_25371 ), .Q ( new_AGEMA_signal_25372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8775 ( .C ( clk ), .D ( new_AGEMA_signal_25549 ), .Q ( new_AGEMA_signal_25550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8795 ( .C ( clk ), .D ( new_AGEMA_signal_25569 ), .Q ( new_AGEMA_signal_25570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8815 ( .C ( clk ), .D ( new_AGEMA_signal_25589 ), .Q ( new_AGEMA_signal_25590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8835 ( .C ( clk ), .D ( new_AGEMA_signal_25609 ), .Q ( new_AGEMA_signal_25610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8855 ( .C ( clk ), .D ( new_AGEMA_signal_25629 ), .Q ( new_AGEMA_signal_25630 ) ) ;

    /* cells in depth 16 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2003 ( .ina ({new_AGEMA_signal_22481, new_AGEMA_signal_22475, new_AGEMA_signal_22469, new_AGEMA_signal_22463, new_AGEMA_signal_22457}), .inb ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, new_AGEMA_signal_4079, new_AGEMA_signal_4078, n1935}), .clk ( clk ), .rnd ({Fresh[11474], Fresh[11473], Fresh[11472], Fresh[11471], Fresh[11470], Fresh[11469], Fresh[11468], Fresh[11467], Fresh[11466], Fresh[11465], Fresh[11464], Fresh[11463], Fresh[11462], Fresh[11461], Fresh[11460]}), .outt ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, new_AGEMA_signal_4251, new_AGEMA_signal_4250, n1941}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2059 ( .ina ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, new_AGEMA_signal_4083, new_AGEMA_signal_4082, n1959}), .inb ({new_AGEMA_signal_22491, new_AGEMA_signal_22489, new_AGEMA_signal_22487, new_AGEMA_signal_22485, new_AGEMA_signal_22483}), .clk ( clk ), .rnd ({Fresh[11489], Fresh[11488], Fresh[11487], Fresh[11486], Fresh[11485], Fresh[11484], Fresh[11483], Fresh[11482], Fresh[11481], Fresh[11480], Fresh[11479], Fresh[11478], Fresh[11477], Fresh[11476], Fresh[11475]}), .outt ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, new_AGEMA_signal_4254, n1960}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2110 ( .ina ({new_AGEMA_signal_22511, new_AGEMA_signal_22507, new_AGEMA_signal_22503, new_AGEMA_signal_22499, new_AGEMA_signal_22495}), .inb ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, new_AGEMA_signal_4086, n1983}), .clk ( clk ), .rnd ({Fresh[11504], Fresh[11503], Fresh[11502], Fresh[11501], Fresh[11500], Fresh[11499], Fresh[11498], Fresh[11497], Fresh[11496], Fresh[11495], Fresh[11494], Fresh[11493], Fresh[11492], Fresh[11491], Fresh[11490]}), .outt ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, new_AGEMA_signal_4259, new_AGEMA_signal_4258, n1988}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2153 ( .ina ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, new_AGEMA_signal_4091, new_AGEMA_signal_4090, n2014}), .inb ({new_AGEMA_signal_22551, new_AGEMA_signal_22543, new_AGEMA_signal_22535, new_AGEMA_signal_22527, new_AGEMA_signal_22519}), .clk ( clk ), .rnd ({Fresh[11519], Fresh[11518], Fresh[11517], Fresh[11516], Fresh[11515], Fresh[11514], Fresh[11513], Fresh[11512], Fresh[11511], Fresh[11510], Fresh[11509], Fresh[11508], Fresh[11507], Fresh[11506], Fresh[11505]}), .outt ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, new_AGEMA_signal_4263, new_AGEMA_signal_4262, n2015}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2169 ( .ina ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, new_AGEMA_signal_3866, n2029}), .inb ({new_AGEMA_signal_22591, new_AGEMA_signal_22583, new_AGEMA_signal_22575, new_AGEMA_signal_22567, new_AGEMA_signal_22559}), .clk ( clk ), .rnd ({Fresh[11534], Fresh[11533], Fresh[11532], Fresh[11531], Fresh[11530], Fresh[11529], Fresh[11528], Fresh[11527], Fresh[11526], Fresh[11525], Fresh[11524], Fresh[11523], Fresh[11522], Fresh[11521], Fresh[11520]}), .outt ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, n2030}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2200 ( .ina ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, new_AGEMA_signal_4103, new_AGEMA_signal_4102, n2052}), .inb ({new_AGEMA_signal_22631, new_AGEMA_signal_22623, new_AGEMA_signal_22615, new_AGEMA_signal_22607, new_AGEMA_signal_22599}), .clk ( clk ), .rnd ({Fresh[11549], Fresh[11548], Fresh[11547], Fresh[11546], Fresh[11545], Fresh[11544], Fresh[11543], Fresh[11542], Fresh[11541], Fresh[11540], Fresh[11539], Fresh[11538], Fresh[11537], Fresh[11536], Fresh[11535]}), .outt ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, new_AGEMA_signal_4271, new_AGEMA_signal_4270, n2053}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2222 ( .ina ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, new_AGEMA_signal_4107, new_AGEMA_signal_4106, n2070}), .inb ({new_AGEMA_signal_22671, new_AGEMA_signal_22663, new_AGEMA_signal_22655, new_AGEMA_signal_22647, new_AGEMA_signal_22639}), .clk ( clk ), .rnd ({Fresh[11564], Fresh[11563], Fresh[11562], Fresh[11561], Fresh[11560], Fresh[11559], Fresh[11558], Fresh[11557], Fresh[11556], Fresh[11555], Fresh[11554], Fresh[11553], Fresh[11552], Fresh[11551], Fresh[11550]}), .outt ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, n2071}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2259 ( .ina ({new_AGEMA_signal_22701, new_AGEMA_signal_22695, new_AGEMA_signal_22689, new_AGEMA_signal_22683, new_AGEMA_signal_22677}), .inb ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, new_AGEMA_signal_4110, n2098}), .clk ( clk ), .rnd ({Fresh[11579], Fresh[11578], Fresh[11577], Fresh[11576], Fresh[11575], Fresh[11574], Fresh[11573], Fresh[11572], Fresh[11571], Fresh[11570], Fresh[11569], Fresh[11568], Fresh[11567], Fresh[11566], Fresh[11565]}), .outt ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, new_AGEMA_signal_4278, n2103}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2288 ( .ina ({new_AGEMA_signal_22751, new_AGEMA_signal_22741, new_AGEMA_signal_22731, new_AGEMA_signal_22721, new_AGEMA_signal_22711}), .inb ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, new_AGEMA_signal_4119, new_AGEMA_signal_4118, n2125}), .clk ( clk ), .rnd ({Fresh[11594], Fresh[11593], Fresh[11592], Fresh[11591], Fresh[11590], Fresh[11589], Fresh[11588], Fresh[11587], Fresh[11586], Fresh[11585], Fresh[11584], Fresh[11583], Fresh[11582], Fresh[11581], Fresh[11580]}), .outt ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, new_AGEMA_signal_4282, n2126}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2314 ( .ina ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, new_AGEMA_signal_4122, n2145}), .inb ({new_AGEMA_signal_22791, new_AGEMA_signal_22783, new_AGEMA_signal_22775, new_AGEMA_signal_22767, new_AGEMA_signal_22759}), .clk ( clk ), .rnd ({Fresh[11609], Fresh[11608], Fresh[11607], Fresh[11606], Fresh[11605], Fresh[11604], Fresh[11603], Fresh[11602], Fresh[11601], Fresh[11600], Fresh[11599], Fresh[11598], Fresh[11597], Fresh[11596], Fresh[11595]}), .outt ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, new_AGEMA_signal_4287, new_AGEMA_signal_4286, n2146}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2334 ( .ina ({new_AGEMA_signal_22831, new_AGEMA_signal_22823, new_AGEMA_signal_22815, new_AGEMA_signal_22807, new_AGEMA_signal_22799}), .inb ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, new_AGEMA_signal_4127, new_AGEMA_signal_4126, n2169}), .clk ( clk ), .rnd ({Fresh[11624], Fresh[11623], Fresh[11622], Fresh[11621], Fresh[11620], Fresh[11619], Fresh[11618], Fresh[11617], Fresh[11616], Fresh[11615], Fresh[11614], Fresh[11613], Fresh[11612], Fresh[11611], Fresh[11610]}), .outt ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, new_AGEMA_signal_4290, n2173}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2351 ( .ina ({new_AGEMA_signal_22871, new_AGEMA_signal_22863, new_AGEMA_signal_22855, new_AGEMA_signal_22847, new_AGEMA_signal_22839}), .inb ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, new_AGEMA_signal_4131, new_AGEMA_signal_4130, n2185}), .clk ( clk ), .rnd ({Fresh[11639], Fresh[11638], Fresh[11637], Fresh[11636], Fresh[11635], Fresh[11634], Fresh[11633], Fresh[11632], Fresh[11631], Fresh[11630], Fresh[11629], Fresh[11628], Fresh[11627], Fresh[11626], Fresh[11625]}), .outt ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, new_AGEMA_signal_4295, new_AGEMA_signal_4294, n2187}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2416 ( .ina ({new_AGEMA_signal_22881, new_AGEMA_signal_22879, new_AGEMA_signal_22877, new_AGEMA_signal_22875, new_AGEMA_signal_22873}), .inb ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, new_AGEMA_signal_4151, new_AGEMA_signal_4150, n2251}), .clk ( clk ), .rnd ({Fresh[11654], Fresh[11653], Fresh[11652], Fresh[11651], Fresh[11650], Fresh[11649], Fresh[11648], Fresh[11647], Fresh[11646], Fresh[11645], Fresh[11644], Fresh[11643], Fresh[11642], Fresh[11641], Fresh[11640]}), .outt ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, new_AGEMA_signal_4302, n2256}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2441 ( .ina ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, new_AGEMA_signal_4155, new_AGEMA_signal_4154, n2274}), .inb ({new_AGEMA_signal_22901, new_AGEMA_signal_22897, new_AGEMA_signal_22893, new_AGEMA_signal_22889, new_AGEMA_signal_22885}), .clk ( clk ), .rnd ({Fresh[11669], Fresh[11668], Fresh[11667], Fresh[11666], Fresh[11665], Fresh[11664], Fresh[11663], Fresh[11662], Fresh[11661], Fresh[11660], Fresh[11659], Fresh[11658], Fresh[11657], Fresh[11656], Fresh[11655]}), .outt ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, new_AGEMA_signal_4307, new_AGEMA_signal_4306, n2275}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2474 ( .ina ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, new_AGEMA_signal_4158, n2302}), .inb ({new_AGEMA_signal_22931, new_AGEMA_signal_22925, new_AGEMA_signal_22919, new_AGEMA_signal_22913, new_AGEMA_signal_22907}), .clk ( clk ), .rnd ({Fresh[11684], Fresh[11683], Fresh[11682], Fresh[11681], Fresh[11680], Fresh[11679], Fresh[11678], Fresh[11677], Fresh[11676], Fresh[11675], Fresh[11674], Fresh[11673], Fresh[11672], Fresh[11671], Fresh[11670]}), .outt ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, n2303}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2504 ( .ina ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, new_AGEMA_signal_4163, new_AGEMA_signal_4162, n2339}), .inb ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, new_AGEMA_signal_4167, new_AGEMA_signal_4166, n2338}), .clk ( clk ), .rnd ({Fresh[11699], Fresh[11698], Fresh[11697], Fresh[11696], Fresh[11695], Fresh[11694], Fresh[11693], Fresh[11692], Fresh[11691], Fresh[11690], Fresh[11689], Fresh[11688], Fresh[11687], Fresh[11686], Fresh[11685]}), .outt ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, new_AGEMA_signal_4315, new_AGEMA_signal_4314, n2382}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2516 ( .ina ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, new_AGEMA_signal_4170, n2351}), .inb ({new_AGEMA_signal_22951, new_AGEMA_signal_22947, new_AGEMA_signal_22943, new_AGEMA_signal_22939, new_AGEMA_signal_22935}), .clk ( clk ), .rnd ({Fresh[11714], Fresh[11713], Fresh[11712], Fresh[11711], Fresh[11710], Fresh[11709], Fresh[11708], Fresh[11707], Fresh[11706], Fresh[11705], Fresh[11704], Fresh[11703], Fresh[11702], Fresh[11701], Fresh[11700]}), .outt ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, new_AGEMA_signal_4319, new_AGEMA_signal_4318, n2380}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2531 ( .ina ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, new_AGEMA_signal_4175, new_AGEMA_signal_4174, n2365}), .inb ({new_AGEMA_signal_23001, new_AGEMA_signal_22991, new_AGEMA_signal_22981, new_AGEMA_signal_22971, new_AGEMA_signal_22961}), .clk ( clk ), .rnd ({Fresh[11729], Fresh[11728], Fresh[11727], Fresh[11726], Fresh[11725], Fresh[11724], Fresh[11723], Fresh[11722], Fresh[11721], Fresh[11720], Fresh[11719], Fresh[11718], Fresh[11717], Fresh[11716], Fresh[11715]}), .outt ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, new_AGEMA_signal_4323, new_AGEMA_signal_4322, n2366}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2561 ( .ina ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, new_AGEMA_signal_3971, new_AGEMA_signal_3970, n2399}), .inb ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, new_AGEMA_signal_4179, new_AGEMA_signal_4178, n2398}), .clk ( clk ), .rnd ({Fresh[11744], Fresh[11743], Fresh[11742], Fresh[11741], Fresh[11740], Fresh[11739], Fresh[11738], Fresh[11737], Fresh[11736], Fresh[11735], Fresh[11734], Fresh[11733], Fresh[11732], Fresh[11731], Fresh[11730]}), .outt ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, new_AGEMA_signal_4326, n2425}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2582 ( .ina ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, new_AGEMA_signal_3979, new_AGEMA_signal_3978, n2423}), .inb ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, new_AGEMA_signal_3983, new_AGEMA_signal_3982, n2422}), .clk ( clk ), .rnd ({Fresh[11759], Fresh[11758], Fresh[11757], Fresh[11756], Fresh[11755], Fresh[11754], Fresh[11753], Fresh[11752], Fresh[11751], Fresh[11750], Fresh[11749], Fresh[11748], Fresh[11747], Fresh[11746], Fresh[11745]}), .outt ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, new_AGEMA_signal_4182, n2424}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2597 ( .ina ({new_AGEMA_signal_23041, new_AGEMA_signal_23033, new_AGEMA_signal_23025, new_AGEMA_signal_23017, new_AGEMA_signal_23009}), .inb ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, new_AGEMA_signal_4187, new_AGEMA_signal_4186, n2441}), .clk ( clk ), .rnd ({Fresh[11774], Fresh[11773], Fresh[11772], Fresh[11771], Fresh[11770], Fresh[11769], Fresh[11768], Fresh[11767], Fresh[11766], Fresh[11765], Fresh[11764], Fresh[11763], Fresh[11762], Fresh[11761], Fresh[11760]}), .outt ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, new_AGEMA_signal_4331, new_AGEMA_signal_4330, n2451}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2631 ( .ina ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_3995, new_AGEMA_signal_3994, n2479}), .inb ({new_AGEMA_signal_23061, new_AGEMA_signal_23057, new_AGEMA_signal_23053, new_AGEMA_signal_23049, new_AGEMA_signal_23045}), .clk ( clk ), .rnd ({Fresh[11789], Fresh[11788], Fresh[11787], Fresh[11786], Fresh[11785], Fresh[11784], Fresh[11783], Fresh[11782], Fresh[11781], Fresh[11780], Fresh[11779], Fresh[11778], Fresh[11777], Fresh[11776], Fresh[11775]}), .outt ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, new_AGEMA_signal_4191, new_AGEMA_signal_4190, n2514}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2658 ( .ina ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, new_AGEMA_signal_4199, new_AGEMA_signal_4198, n2510}), .inb ({new_AGEMA_signal_23071, new_AGEMA_signal_23069, new_AGEMA_signal_23067, new_AGEMA_signal_23065, new_AGEMA_signal_23063}), .clk ( clk ), .rnd ({Fresh[11804], Fresh[11803], Fresh[11802], Fresh[11801], Fresh[11800], Fresh[11799], Fresh[11798], Fresh[11797], Fresh[11796], Fresh[11795], Fresh[11794], Fresh[11793], Fresh[11792], Fresh[11791], Fresh[11790]}), .outt ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, new_AGEMA_signal_4335, new_AGEMA_signal_4334, n2511}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2688 ( .ina ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, new_AGEMA_signal_4211, new_AGEMA_signal_4210, n2552}), .inb ({new_AGEMA_signal_23111, new_AGEMA_signal_23103, new_AGEMA_signal_23095, new_AGEMA_signal_23087, new_AGEMA_signal_23079}), .clk ( clk ), .rnd ({Fresh[11819], Fresh[11818], Fresh[11817], Fresh[11816], Fresh[11815], Fresh[11814], Fresh[11813], Fresh[11812], Fresh[11811], Fresh[11810], Fresh[11809], Fresh[11808], Fresh[11807], Fresh[11806], Fresh[11805]}), .outt ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, new_AGEMA_signal_4339, new_AGEMA_signal_4338, n2671}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2716 ( .ina ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, new_AGEMA_signal_4218, n2589}), .inb ({new_AGEMA_signal_23151, new_AGEMA_signal_23143, new_AGEMA_signal_23135, new_AGEMA_signal_23127, new_AGEMA_signal_23119}), .clk ( clk ), .rnd ({Fresh[11834], Fresh[11833], Fresh[11832], Fresh[11831], Fresh[11830], Fresh[11829], Fresh[11828], Fresh[11827], Fresh[11826], Fresh[11825], Fresh[11824], Fresh[11823], Fresh[11822], Fresh[11821], Fresh[11820]}), .outt ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, new_AGEMA_signal_4343, new_AGEMA_signal_4342, n2590}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2731 ( .ina ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_4031, new_AGEMA_signal_4030, n2608}), .inb ({new_AGEMA_signal_23181, new_AGEMA_signal_23175, new_AGEMA_signal_23169, new_AGEMA_signal_23163, new_AGEMA_signal_23157}), .clk ( clk ), .rnd ({Fresh[11849], Fresh[11848], Fresh[11847], Fresh[11846], Fresh[11845], Fresh[11844], Fresh[11843], Fresh[11842], Fresh[11841], Fresh[11840], Fresh[11839], Fresh[11838], Fresh[11837], Fresh[11836], Fresh[11835]}), .outt ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, new_AGEMA_signal_4223, new_AGEMA_signal_4222, n2623}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2763 ( .ina ({new_AGEMA_signal_23201, new_AGEMA_signal_23197, new_AGEMA_signal_23193, new_AGEMA_signal_23189, new_AGEMA_signal_23185}), .inb ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, new_AGEMA_signal_4230, n2659}), .clk ( clk ), .rnd ({Fresh[11864], Fresh[11863], Fresh[11862], Fresh[11861], Fresh[11860], Fresh[11859], Fresh[11858], Fresh[11857], Fresh[11856], Fresh[11855], Fresh[11854], Fresh[11853], Fresh[11852], Fresh[11851], Fresh[11850]}), .outt ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, new_AGEMA_signal_4350, n2667}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2786 ( .ina ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, new_AGEMA_signal_4235, new_AGEMA_signal_4234, n2702}), .inb ({new_AGEMA_signal_23241, new_AGEMA_signal_23233, new_AGEMA_signal_23225, new_AGEMA_signal_23217, new_AGEMA_signal_23209}), .clk ( clk ), .rnd ({Fresh[11879], Fresh[11878], Fresh[11877], Fresh[11876], Fresh[11875], Fresh[11874], Fresh[11873], Fresh[11872], Fresh[11871], Fresh[11870], Fresh[11869], Fresh[11868], Fresh[11867], Fresh[11866], Fresh[11865]}), .outt ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, new_AGEMA_signal_4354, n2703}) ) ;
    mux2_HPC1 #(.security_order(4), .pipeline(1)) U2840 ( .ins ({new_AGEMA_signal_22901, new_AGEMA_signal_22897, new_AGEMA_signal_22893, new_AGEMA_signal_22889, new_AGEMA_signal_22885}), .inb ({new_AGEMA_signal_23251, new_AGEMA_signal_23249, new_AGEMA_signal_23247, new_AGEMA_signal_23245, new_AGEMA_signal_23243}), .ina ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, new_AGEMA_signal_4071, new_AGEMA_signal_4070, n2801}), .clk ( clk ), .rnd ({Fresh[11894], Fresh[11893], Fresh[11892], Fresh[11891], Fresh[11890], Fresh[11889], Fresh[11888], Fresh[11887], Fresh[11886], Fresh[11885], Fresh[11884], Fresh[11883], Fresh[11882], Fresh[11881], Fresh[11880]}), .outt ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, new_AGEMA_signal_4242, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C ( clk ), .D ( new_AGEMA_signal_23256 ), .Q ( new_AGEMA_signal_23257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C ( clk ), .D ( new_AGEMA_signal_23262 ), .Q ( new_AGEMA_signal_23263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C ( clk ), .D ( new_AGEMA_signal_23268 ), .Q ( new_AGEMA_signal_23269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C ( clk ), .D ( new_AGEMA_signal_23274 ), .Q ( new_AGEMA_signal_23275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C ( clk ), .D ( new_AGEMA_signal_23280 ), .Q ( new_AGEMA_signal_23281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C ( clk ), .D ( new_AGEMA_signal_23286 ), .Q ( new_AGEMA_signal_23287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C ( clk ), .D ( new_AGEMA_signal_23292 ), .Q ( new_AGEMA_signal_23293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C ( clk ), .D ( new_AGEMA_signal_23298 ), .Q ( new_AGEMA_signal_23299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C ( clk ), .D ( new_AGEMA_signal_23304 ), .Q ( new_AGEMA_signal_23305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C ( clk ), .D ( new_AGEMA_signal_23310 ), .Q ( new_AGEMA_signal_23311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C ( clk ), .D ( new_AGEMA_signal_23316 ), .Q ( new_AGEMA_signal_23317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C ( clk ), .D ( new_AGEMA_signal_23322 ), .Q ( new_AGEMA_signal_23323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C ( clk ), .D ( new_AGEMA_signal_23328 ), .Q ( new_AGEMA_signal_23329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C ( clk ), .D ( new_AGEMA_signal_23334 ), .Q ( new_AGEMA_signal_23335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C ( clk ), .D ( new_AGEMA_signal_23340 ), .Q ( new_AGEMA_signal_23341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C ( clk ), .D ( new_AGEMA_signal_23344 ), .Q ( new_AGEMA_signal_23345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C ( clk ), .D ( new_AGEMA_signal_23348 ), .Q ( new_AGEMA_signal_23349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C ( clk ), .D ( new_AGEMA_signal_23352 ), .Q ( new_AGEMA_signal_23353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C ( clk ), .D ( new_AGEMA_signal_23356 ), .Q ( new_AGEMA_signal_23357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C ( clk ), .D ( new_AGEMA_signal_23360 ), .Q ( new_AGEMA_signal_23361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C ( clk ), .D ( new_AGEMA_signal_23368 ), .Q ( new_AGEMA_signal_23369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C ( clk ), .D ( new_AGEMA_signal_23376 ), .Q ( new_AGEMA_signal_23377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C ( clk ), .D ( new_AGEMA_signal_23384 ), .Q ( new_AGEMA_signal_23385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C ( clk ), .D ( new_AGEMA_signal_23392 ), .Q ( new_AGEMA_signal_23393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C ( clk ), .D ( new_AGEMA_signal_23400 ), .Q ( new_AGEMA_signal_23401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C ( clk ), .D ( new_AGEMA_signal_23406 ), .Q ( new_AGEMA_signal_23407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C ( clk ), .D ( new_AGEMA_signal_23412 ), .Q ( new_AGEMA_signal_23413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C ( clk ), .D ( new_AGEMA_signal_23418 ), .Q ( new_AGEMA_signal_23419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C ( clk ), .D ( new_AGEMA_signal_23424 ), .Q ( new_AGEMA_signal_23425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C ( clk ), .D ( new_AGEMA_signal_23430 ), .Q ( new_AGEMA_signal_23431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C ( clk ), .D ( new_AGEMA_signal_23434 ), .Q ( new_AGEMA_signal_23435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C ( clk ), .D ( new_AGEMA_signal_23438 ), .Q ( new_AGEMA_signal_23439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C ( clk ), .D ( new_AGEMA_signal_23442 ), .Q ( new_AGEMA_signal_23443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C ( clk ), .D ( new_AGEMA_signal_23446 ), .Q ( new_AGEMA_signal_23447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C ( clk ), .D ( new_AGEMA_signal_23450 ), .Q ( new_AGEMA_signal_23451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C ( clk ), .D ( new_AGEMA_signal_23458 ), .Q ( new_AGEMA_signal_23459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C ( clk ), .D ( new_AGEMA_signal_23466 ), .Q ( new_AGEMA_signal_23467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C ( clk ), .D ( new_AGEMA_signal_23474 ), .Q ( new_AGEMA_signal_23475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C ( clk ), .D ( new_AGEMA_signal_23482 ), .Q ( new_AGEMA_signal_23483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C ( clk ), .D ( new_AGEMA_signal_23490 ), .Q ( new_AGEMA_signal_23491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C ( clk ), .D ( new_AGEMA_signal_23498 ), .Q ( new_AGEMA_signal_23499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C ( clk ), .D ( new_AGEMA_signal_23506 ), .Q ( new_AGEMA_signal_23507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C ( clk ), .D ( new_AGEMA_signal_23514 ), .Q ( new_AGEMA_signal_23515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C ( clk ), .D ( new_AGEMA_signal_23522 ), .Q ( new_AGEMA_signal_23523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C ( clk ), .D ( new_AGEMA_signal_23530 ), .Q ( new_AGEMA_signal_23531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C ( clk ), .D ( new_AGEMA_signal_23540 ), .Q ( new_AGEMA_signal_23541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C ( clk ), .D ( new_AGEMA_signal_23550 ), .Q ( new_AGEMA_signal_23551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C ( clk ), .D ( new_AGEMA_signal_23560 ), .Q ( new_AGEMA_signal_23561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C ( clk ), .D ( new_AGEMA_signal_23570 ), .Q ( new_AGEMA_signal_23571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C ( clk ), .D ( new_AGEMA_signal_23580 ), .Q ( new_AGEMA_signal_23581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C ( clk ), .D ( new_AGEMA_signal_23588 ), .Q ( new_AGEMA_signal_23589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C ( clk ), .D ( new_AGEMA_signal_23596 ), .Q ( new_AGEMA_signal_23597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C ( clk ), .D ( new_AGEMA_signal_23604 ), .Q ( new_AGEMA_signal_23605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C ( clk ), .D ( new_AGEMA_signal_23612 ), .Q ( new_AGEMA_signal_23613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C ( clk ), .D ( new_AGEMA_signal_23620 ), .Q ( new_AGEMA_signal_23621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C ( clk ), .D ( new_AGEMA_signal_23626 ), .Q ( new_AGEMA_signal_23627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C ( clk ), .D ( new_AGEMA_signal_23632 ), .Q ( new_AGEMA_signal_23633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C ( clk ), .D ( new_AGEMA_signal_23638 ), .Q ( new_AGEMA_signal_23639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C ( clk ), .D ( new_AGEMA_signal_23644 ), .Q ( new_AGEMA_signal_23645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C ( clk ), .D ( new_AGEMA_signal_23650 ), .Q ( new_AGEMA_signal_23651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C ( clk ), .D ( new_AGEMA_signal_23654 ), .Q ( new_AGEMA_signal_23655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C ( clk ), .D ( new_AGEMA_signal_23658 ), .Q ( new_AGEMA_signal_23659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C ( clk ), .D ( new_AGEMA_signal_23662 ), .Q ( new_AGEMA_signal_23663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C ( clk ), .D ( new_AGEMA_signal_23666 ), .Q ( new_AGEMA_signal_23667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C ( clk ), .D ( new_AGEMA_signal_23670 ), .Q ( new_AGEMA_signal_23671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C ( clk ), .D ( new_AGEMA_signal_23676 ), .Q ( new_AGEMA_signal_23677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C ( clk ), .D ( new_AGEMA_signal_23682 ), .Q ( new_AGEMA_signal_23683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C ( clk ), .D ( new_AGEMA_signal_23688 ), .Q ( new_AGEMA_signal_23689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C ( clk ), .D ( new_AGEMA_signal_23694 ), .Q ( new_AGEMA_signal_23695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C ( clk ), .D ( new_AGEMA_signal_23700 ), .Q ( new_AGEMA_signal_23701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C ( clk ), .D ( new_AGEMA_signal_23708 ), .Q ( new_AGEMA_signal_23709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C ( clk ), .D ( new_AGEMA_signal_23716 ), .Q ( new_AGEMA_signal_23717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C ( clk ), .D ( new_AGEMA_signal_23724 ), .Q ( new_AGEMA_signal_23725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C ( clk ), .D ( new_AGEMA_signal_23732 ), .Q ( new_AGEMA_signal_23733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C ( clk ), .D ( new_AGEMA_signal_23740 ), .Q ( new_AGEMA_signal_23741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C ( clk ), .D ( new_AGEMA_signal_23746 ), .Q ( new_AGEMA_signal_23747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C ( clk ), .D ( new_AGEMA_signal_23752 ), .Q ( new_AGEMA_signal_23753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C ( clk ), .D ( new_AGEMA_signal_23758 ), .Q ( new_AGEMA_signal_23759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C ( clk ), .D ( new_AGEMA_signal_23764 ), .Q ( new_AGEMA_signal_23765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C ( clk ), .D ( new_AGEMA_signal_23770 ), .Q ( new_AGEMA_signal_23771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C ( clk ), .D ( new_AGEMA_signal_23772 ), .Q ( new_AGEMA_signal_23773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C ( clk ), .D ( new_AGEMA_signal_23774 ), .Q ( new_AGEMA_signal_23775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C ( clk ), .D ( new_AGEMA_signal_23776 ), .Q ( new_AGEMA_signal_23777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C ( clk ), .D ( new_AGEMA_signal_23778 ), .Q ( new_AGEMA_signal_23779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C ( clk ), .D ( new_AGEMA_signal_23780 ), .Q ( new_AGEMA_signal_23781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C ( clk ), .D ( new_AGEMA_signal_23788 ), .Q ( new_AGEMA_signal_23789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C ( clk ), .D ( new_AGEMA_signal_23796 ), .Q ( new_AGEMA_signal_23797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C ( clk ), .D ( new_AGEMA_signal_23804 ), .Q ( new_AGEMA_signal_23805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C ( clk ), .D ( new_AGEMA_signal_23812 ), .Q ( new_AGEMA_signal_23813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C ( clk ), .D ( new_AGEMA_signal_23820 ), .Q ( new_AGEMA_signal_23821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C ( clk ), .D ( new_AGEMA_signal_23824 ), .Q ( new_AGEMA_signal_23825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C ( clk ), .D ( new_AGEMA_signal_23828 ), .Q ( new_AGEMA_signal_23829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C ( clk ), .D ( new_AGEMA_signal_23832 ), .Q ( new_AGEMA_signal_23833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C ( clk ), .D ( new_AGEMA_signal_23836 ), .Q ( new_AGEMA_signal_23837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C ( clk ), .D ( new_AGEMA_signal_23840 ), .Q ( new_AGEMA_signal_23841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C ( clk ), .D ( new_AGEMA_signal_23846 ), .Q ( new_AGEMA_signal_23847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C ( clk ), .D ( new_AGEMA_signal_23852 ), .Q ( new_AGEMA_signal_23853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C ( clk ), .D ( new_AGEMA_signal_23858 ), .Q ( new_AGEMA_signal_23859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C ( clk ), .D ( new_AGEMA_signal_23864 ), .Q ( new_AGEMA_signal_23865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C ( clk ), .D ( new_AGEMA_signal_23870 ), .Q ( new_AGEMA_signal_23871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C ( clk ), .D ( new_AGEMA_signal_23876 ), .Q ( new_AGEMA_signal_23877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C ( clk ), .D ( new_AGEMA_signal_23882 ), .Q ( new_AGEMA_signal_23883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C ( clk ), .D ( new_AGEMA_signal_23888 ), .Q ( new_AGEMA_signal_23889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C ( clk ), .D ( new_AGEMA_signal_23894 ), .Q ( new_AGEMA_signal_23895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C ( clk ), .D ( new_AGEMA_signal_23900 ), .Q ( new_AGEMA_signal_23901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C ( clk ), .D ( new_AGEMA_signal_23904 ), .Q ( new_AGEMA_signal_23905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C ( clk ), .D ( new_AGEMA_signal_23908 ), .Q ( new_AGEMA_signal_23909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C ( clk ), .D ( new_AGEMA_signal_23912 ), .Q ( new_AGEMA_signal_23913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C ( clk ), .D ( new_AGEMA_signal_23916 ), .Q ( new_AGEMA_signal_23917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C ( clk ), .D ( new_AGEMA_signal_23920 ), .Q ( new_AGEMA_signal_23921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C ( clk ), .D ( new_AGEMA_signal_23924 ), .Q ( new_AGEMA_signal_23925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C ( clk ), .D ( new_AGEMA_signal_23930 ), .Q ( new_AGEMA_signal_23931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C ( clk ), .D ( new_AGEMA_signal_23936 ), .Q ( new_AGEMA_signal_23937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C ( clk ), .D ( new_AGEMA_signal_23942 ), .Q ( new_AGEMA_signal_23943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C ( clk ), .D ( new_AGEMA_signal_23948 ), .Q ( new_AGEMA_signal_23949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C ( clk ), .D ( new_AGEMA_signal_23952 ), .Q ( new_AGEMA_signal_23953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C ( clk ), .D ( new_AGEMA_signal_23956 ), .Q ( new_AGEMA_signal_23957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C ( clk ), .D ( new_AGEMA_signal_23960 ), .Q ( new_AGEMA_signal_23961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C ( clk ), .D ( new_AGEMA_signal_23964 ), .Q ( new_AGEMA_signal_23965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C ( clk ), .D ( new_AGEMA_signal_23968 ), .Q ( new_AGEMA_signal_23969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C ( clk ), .D ( new_AGEMA_signal_23974 ), .Q ( new_AGEMA_signal_23975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C ( clk ), .D ( new_AGEMA_signal_23980 ), .Q ( new_AGEMA_signal_23981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C ( clk ), .D ( new_AGEMA_signal_23986 ), .Q ( new_AGEMA_signal_23987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C ( clk ), .D ( new_AGEMA_signal_23992 ), .Q ( new_AGEMA_signal_23993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C ( clk ), .D ( new_AGEMA_signal_23998 ), .Q ( new_AGEMA_signal_23999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C ( clk ), .D ( new_AGEMA_signal_24008 ), .Q ( new_AGEMA_signal_24009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C ( clk ), .D ( new_AGEMA_signal_24018 ), .Q ( new_AGEMA_signal_24019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C ( clk ), .D ( new_AGEMA_signal_24028 ), .Q ( new_AGEMA_signal_24029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C ( clk ), .D ( new_AGEMA_signal_24038 ), .Q ( new_AGEMA_signal_24039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C ( clk ), .D ( new_AGEMA_signal_24048 ), .Q ( new_AGEMA_signal_24049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C ( clk ), .D ( new_AGEMA_signal_24054 ), .Q ( new_AGEMA_signal_24055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C ( clk ), .D ( new_AGEMA_signal_24060 ), .Q ( new_AGEMA_signal_24061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C ( clk ), .D ( new_AGEMA_signal_24066 ), .Q ( new_AGEMA_signal_24067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C ( clk ), .D ( new_AGEMA_signal_24072 ), .Q ( new_AGEMA_signal_24073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C ( clk ), .D ( new_AGEMA_signal_24078 ), .Q ( new_AGEMA_signal_24079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C ( clk ), .D ( new_AGEMA_signal_24084 ), .Q ( new_AGEMA_signal_24085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C ( clk ), .D ( new_AGEMA_signal_24090 ), .Q ( new_AGEMA_signal_24091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C ( clk ), .D ( new_AGEMA_signal_24096 ), .Q ( new_AGEMA_signal_24097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C ( clk ), .D ( new_AGEMA_signal_24102 ), .Q ( new_AGEMA_signal_24103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C ( clk ), .D ( new_AGEMA_signal_24108 ), .Q ( new_AGEMA_signal_24109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C ( clk ), .D ( new_AGEMA_signal_24112 ), .Q ( new_AGEMA_signal_24113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C ( clk ), .D ( new_AGEMA_signal_24116 ), .Q ( new_AGEMA_signal_24117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C ( clk ), .D ( new_AGEMA_signal_24120 ), .Q ( new_AGEMA_signal_24121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C ( clk ), .D ( new_AGEMA_signal_24124 ), .Q ( new_AGEMA_signal_24125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C ( clk ), .D ( new_AGEMA_signal_24128 ), .Q ( new_AGEMA_signal_24129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C ( clk ), .D ( new_AGEMA_signal_24132 ), .Q ( new_AGEMA_signal_24133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C ( clk ), .D ( new_AGEMA_signal_24136 ), .Q ( new_AGEMA_signal_24137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C ( clk ), .D ( new_AGEMA_signal_24140 ), .Q ( new_AGEMA_signal_24141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C ( clk ), .D ( new_AGEMA_signal_24144 ), .Q ( new_AGEMA_signal_24145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C ( clk ), .D ( new_AGEMA_signal_24148 ), .Q ( new_AGEMA_signal_24149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C ( clk ), .D ( new_AGEMA_signal_24156 ), .Q ( new_AGEMA_signal_24157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C ( clk ), .D ( new_AGEMA_signal_24164 ), .Q ( new_AGEMA_signal_24165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C ( clk ), .D ( new_AGEMA_signal_24172 ), .Q ( new_AGEMA_signal_24173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C ( clk ), .D ( new_AGEMA_signal_24180 ), .Q ( new_AGEMA_signal_24181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C ( clk ), .D ( new_AGEMA_signal_24188 ), .Q ( new_AGEMA_signal_24189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C ( clk ), .D ( new_AGEMA_signal_24194 ), .Q ( new_AGEMA_signal_24195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C ( clk ), .D ( new_AGEMA_signal_24200 ), .Q ( new_AGEMA_signal_24201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C ( clk ), .D ( new_AGEMA_signal_24206 ), .Q ( new_AGEMA_signal_24207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C ( clk ), .D ( new_AGEMA_signal_24212 ), .Q ( new_AGEMA_signal_24213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C ( clk ), .D ( new_AGEMA_signal_24218 ), .Q ( new_AGEMA_signal_24219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C ( clk ), .D ( new_AGEMA_signal_24226 ), .Q ( new_AGEMA_signal_24227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C ( clk ), .D ( new_AGEMA_signal_24234 ), .Q ( new_AGEMA_signal_24235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C ( clk ), .D ( new_AGEMA_signal_24242 ), .Q ( new_AGEMA_signal_24243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C ( clk ), .D ( new_AGEMA_signal_24250 ), .Q ( new_AGEMA_signal_24251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C ( clk ), .D ( new_AGEMA_signal_24258 ), .Q ( new_AGEMA_signal_24259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C ( clk ), .D ( new_AGEMA_signal_24266 ), .Q ( new_AGEMA_signal_24267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C ( clk ), .D ( new_AGEMA_signal_24274 ), .Q ( new_AGEMA_signal_24275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C ( clk ), .D ( new_AGEMA_signal_24282 ), .Q ( new_AGEMA_signal_24283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C ( clk ), .D ( new_AGEMA_signal_24290 ), .Q ( new_AGEMA_signal_24291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C ( clk ), .D ( new_AGEMA_signal_24298 ), .Q ( new_AGEMA_signal_24299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C ( clk ), .D ( new_AGEMA_signal_24312 ), .Q ( new_AGEMA_signal_24313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C ( clk ), .D ( new_AGEMA_signal_24316 ), .Q ( new_AGEMA_signal_24317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C ( clk ), .D ( new_AGEMA_signal_24320 ), .Q ( new_AGEMA_signal_24321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C ( clk ), .D ( new_AGEMA_signal_24324 ), .Q ( new_AGEMA_signal_24325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C ( clk ), .D ( new_AGEMA_signal_24328 ), .Q ( new_AGEMA_signal_24329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C ( clk ), .D ( new_AGEMA_signal_24332 ), .Q ( new_AGEMA_signal_24333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C ( clk ), .D ( new_AGEMA_signal_24336 ), .Q ( new_AGEMA_signal_24337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C ( clk ), .D ( new_AGEMA_signal_24340 ), .Q ( new_AGEMA_signal_24341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C ( clk ), .D ( new_AGEMA_signal_24344 ), .Q ( new_AGEMA_signal_24345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C ( clk ), .D ( new_AGEMA_signal_24348 ), .Q ( new_AGEMA_signal_24349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C ( clk ), .D ( new_AGEMA_signal_24356 ), .Q ( new_AGEMA_signal_24357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C ( clk ), .D ( new_AGEMA_signal_24364 ), .Q ( new_AGEMA_signal_24365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C ( clk ), .D ( new_AGEMA_signal_24372 ), .Q ( new_AGEMA_signal_24373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C ( clk ), .D ( new_AGEMA_signal_24380 ), .Q ( new_AGEMA_signal_24381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C ( clk ), .D ( new_AGEMA_signal_24388 ), .Q ( new_AGEMA_signal_24389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C ( clk ), .D ( new_AGEMA_signal_24392 ), .Q ( new_AGEMA_signal_24393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C ( clk ), .D ( new_AGEMA_signal_24396 ), .Q ( new_AGEMA_signal_24397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C ( clk ), .D ( new_AGEMA_signal_24400 ), .Q ( new_AGEMA_signal_24401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C ( clk ), .D ( new_AGEMA_signal_24404 ), .Q ( new_AGEMA_signal_24405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C ( clk ), .D ( new_AGEMA_signal_24408 ), .Q ( new_AGEMA_signal_24409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C ( clk ), .D ( new_AGEMA_signal_24414 ), .Q ( new_AGEMA_signal_24415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C ( clk ), .D ( new_AGEMA_signal_24422 ), .Q ( new_AGEMA_signal_24423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C ( clk ), .D ( new_AGEMA_signal_24430 ), .Q ( new_AGEMA_signal_24431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7664 ( .C ( clk ), .D ( new_AGEMA_signal_24438 ), .Q ( new_AGEMA_signal_24439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7672 ( .C ( clk ), .D ( new_AGEMA_signal_24446 ), .Q ( new_AGEMA_signal_24447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7684 ( .C ( clk ), .D ( new_AGEMA_signal_24458 ), .Q ( new_AGEMA_signal_24459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7696 ( .C ( clk ), .D ( new_AGEMA_signal_24470 ), .Q ( new_AGEMA_signal_24471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7708 ( .C ( clk ), .D ( new_AGEMA_signal_24482 ), .Q ( new_AGEMA_signal_24483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7720 ( .C ( clk ), .D ( new_AGEMA_signal_24494 ), .Q ( new_AGEMA_signal_24495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7732 ( .C ( clk ), .D ( new_AGEMA_signal_24506 ), .Q ( new_AGEMA_signal_24507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7746 ( .C ( clk ), .D ( new_AGEMA_signal_24520 ), .Q ( new_AGEMA_signal_24521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7760 ( .C ( clk ), .D ( new_AGEMA_signal_24534 ), .Q ( new_AGEMA_signal_24535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7774 ( .C ( clk ), .D ( new_AGEMA_signal_24548 ), .Q ( new_AGEMA_signal_24549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7788 ( .C ( clk ), .D ( new_AGEMA_signal_24562 ), .Q ( new_AGEMA_signal_24563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7802 ( .C ( clk ), .D ( new_AGEMA_signal_24576 ), .Q ( new_AGEMA_signal_24577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7810 ( .C ( clk ), .D ( new_AGEMA_signal_24584 ), .Q ( new_AGEMA_signal_24585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7818 ( .C ( clk ), .D ( new_AGEMA_signal_24592 ), .Q ( new_AGEMA_signal_24593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7826 ( .C ( clk ), .D ( new_AGEMA_signal_24600 ), .Q ( new_AGEMA_signal_24601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7834 ( .C ( clk ), .D ( new_AGEMA_signal_24608 ), .Q ( new_AGEMA_signal_24609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7842 ( .C ( clk ), .D ( new_AGEMA_signal_24616 ), .Q ( new_AGEMA_signal_24617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7856 ( .C ( clk ), .D ( new_AGEMA_signal_24630 ), .Q ( new_AGEMA_signal_24631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7870 ( .C ( clk ), .D ( new_AGEMA_signal_24644 ), .Q ( new_AGEMA_signal_24645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7884 ( .C ( clk ), .D ( new_AGEMA_signal_24658 ), .Q ( new_AGEMA_signal_24659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7898 ( .C ( clk ), .D ( new_AGEMA_signal_24672 ), .Q ( new_AGEMA_signal_24673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7912 ( .C ( clk ), .D ( new_AGEMA_signal_24686 ), .Q ( new_AGEMA_signal_24687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7920 ( .C ( clk ), .D ( new_AGEMA_signal_24694 ), .Q ( new_AGEMA_signal_24695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7928 ( .C ( clk ), .D ( new_AGEMA_signal_24702 ), .Q ( new_AGEMA_signal_24703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7936 ( .C ( clk ), .D ( new_AGEMA_signal_24710 ), .Q ( new_AGEMA_signal_24711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7944 ( .C ( clk ), .D ( new_AGEMA_signal_24718 ), .Q ( new_AGEMA_signal_24719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7952 ( .C ( clk ), .D ( new_AGEMA_signal_24726 ), .Q ( new_AGEMA_signal_24727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7960 ( .C ( clk ), .D ( new_AGEMA_signal_24734 ), .Q ( new_AGEMA_signal_24735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7968 ( .C ( clk ), .D ( new_AGEMA_signal_24742 ), .Q ( new_AGEMA_signal_24743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7976 ( .C ( clk ), .D ( new_AGEMA_signal_24750 ), .Q ( new_AGEMA_signal_24751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7984 ( .C ( clk ), .D ( new_AGEMA_signal_24758 ), .Q ( new_AGEMA_signal_24759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7992 ( .C ( clk ), .D ( new_AGEMA_signal_24766 ), .Q ( new_AGEMA_signal_24767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8036 ( .C ( clk ), .D ( new_AGEMA_signal_24810 ), .Q ( new_AGEMA_signal_24811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8052 ( .C ( clk ), .D ( new_AGEMA_signal_24826 ), .Q ( new_AGEMA_signal_24827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8068 ( .C ( clk ), .D ( new_AGEMA_signal_24842 ), .Q ( new_AGEMA_signal_24843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8084 ( .C ( clk ), .D ( new_AGEMA_signal_24858 ), .Q ( new_AGEMA_signal_24859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8100 ( .C ( clk ), .D ( new_AGEMA_signal_24874 ), .Q ( new_AGEMA_signal_24875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8146 ( .C ( clk ), .D ( new_AGEMA_signal_24920 ), .Q ( new_AGEMA_signal_24921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8162 ( .C ( clk ), .D ( new_AGEMA_signal_24936 ), .Q ( new_AGEMA_signal_24937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8178 ( .C ( clk ), .D ( new_AGEMA_signal_24952 ), .Q ( new_AGEMA_signal_24953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8194 ( .C ( clk ), .D ( new_AGEMA_signal_24968 ), .Q ( new_AGEMA_signal_24969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8210 ( .C ( clk ), .D ( new_AGEMA_signal_24984 ), .Q ( new_AGEMA_signal_24985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8220 ( .C ( clk ), .D ( new_AGEMA_signal_24994 ), .Q ( new_AGEMA_signal_24995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8230 ( .C ( clk ), .D ( new_AGEMA_signal_25004 ), .Q ( new_AGEMA_signal_25005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8240 ( .C ( clk ), .D ( new_AGEMA_signal_25014 ), .Q ( new_AGEMA_signal_25015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8250 ( .C ( clk ), .D ( new_AGEMA_signal_25024 ), .Q ( new_AGEMA_signal_25025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8260 ( .C ( clk ), .D ( new_AGEMA_signal_25034 ), .Q ( new_AGEMA_signal_25035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8288 ( .C ( clk ), .D ( new_AGEMA_signal_25062 ), .Q ( new_AGEMA_signal_25063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8296 ( .C ( clk ), .D ( new_AGEMA_signal_25070 ), .Q ( new_AGEMA_signal_25071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8304 ( .C ( clk ), .D ( new_AGEMA_signal_25078 ), .Q ( new_AGEMA_signal_25079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8312 ( .C ( clk ), .D ( new_AGEMA_signal_25086 ), .Q ( new_AGEMA_signal_25087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8320 ( .C ( clk ), .D ( new_AGEMA_signal_25094 ), .Q ( new_AGEMA_signal_25095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8394 ( .C ( clk ), .D ( new_AGEMA_signal_25168 ), .Q ( new_AGEMA_signal_25169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8410 ( .C ( clk ), .D ( new_AGEMA_signal_25184 ), .Q ( new_AGEMA_signal_25185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8426 ( .C ( clk ), .D ( new_AGEMA_signal_25200 ), .Q ( new_AGEMA_signal_25201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8442 ( .C ( clk ), .D ( new_AGEMA_signal_25216 ), .Q ( new_AGEMA_signal_25217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8458 ( .C ( clk ), .D ( new_AGEMA_signal_25232 ), .Q ( new_AGEMA_signal_25233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8468 ( .C ( clk ), .D ( new_AGEMA_signal_25242 ), .Q ( new_AGEMA_signal_25243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8478 ( .C ( clk ), .D ( new_AGEMA_signal_25252 ), .Q ( new_AGEMA_signal_25253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8488 ( .C ( clk ), .D ( new_AGEMA_signal_25262 ), .Q ( new_AGEMA_signal_25263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8498 ( .C ( clk ), .D ( new_AGEMA_signal_25272 ), .Q ( new_AGEMA_signal_25273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8508 ( .C ( clk ), .D ( new_AGEMA_signal_25282 ), .Q ( new_AGEMA_signal_25283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8526 ( .C ( clk ), .D ( new_AGEMA_signal_25300 ), .Q ( new_AGEMA_signal_25301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8544 ( .C ( clk ), .D ( new_AGEMA_signal_25318 ), .Q ( new_AGEMA_signal_25319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8562 ( .C ( clk ), .D ( new_AGEMA_signal_25336 ), .Q ( new_AGEMA_signal_25337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8580 ( .C ( clk ), .D ( new_AGEMA_signal_25354 ), .Q ( new_AGEMA_signal_25355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8598 ( .C ( clk ), .D ( new_AGEMA_signal_25372 ), .Q ( new_AGEMA_signal_25373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8776 ( .C ( clk ), .D ( new_AGEMA_signal_25550 ), .Q ( new_AGEMA_signal_25551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8796 ( .C ( clk ), .D ( new_AGEMA_signal_25570 ), .Q ( new_AGEMA_signal_25571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8816 ( .C ( clk ), .D ( new_AGEMA_signal_25590 ), .Q ( new_AGEMA_signal_25591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8836 ( .C ( clk ), .D ( new_AGEMA_signal_25610 ), .Q ( new_AGEMA_signal_25611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8856 ( .C ( clk ), .D ( new_AGEMA_signal_25630 ), .Q ( new_AGEMA_signal_25631 ) ) ;

    /* cells in depth 17 */
    buf_clk new_AGEMA_reg_buffer_7151 ( .C ( clk ), .D ( new_AGEMA_signal_23925 ), .Q ( new_AGEMA_signal_23926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C ( clk ), .D ( new_AGEMA_signal_23931 ), .Q ( new_AGEMA_signal_23932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C ( clk ), .D ( new_AGEMA_signal_23937 ), .Q ( new_AGEMA_signal_23938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C ( clk ), .D ( new_AGEMA_signal_23943 ), .Q ( new_AGEMA_signal_23944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C ( clk ), .D ( new_AGEMA_signal_23949 ), .Q ( new_AGEMA_signal_23950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C ( clk ), .D ( new_AGEMA_signal_23953 ), .Q ( new_AGEMA_signal_23954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C ( clk ), .D ( new_AGEMA_signal_23957 ), .Q ( new_AGEMA_signal_23958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C ( clk ), .D ( new_AGEMA_signal_23961 ), .Q ( new_AGEMA_signal_23962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C ( clk ), .D ( new_AGEMA_signal_23965 ), .Q ( new_AGEMA_signal_23966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C ( clk ), .D ( new_AGEMA_signal_23969 ), .Q ( new_AGEMA_signal_23970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C ( clk ), .D ( new_AGEMA_signal_23975 ), .Q ( new_AGEMA_signal_23976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C ( clk ), .D ( new_AGEMA_signal_23981 ), .Q ( new_AGEMA_signal_23982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C ( clk ), .D ( new_AGEMA_signal_23987 ), .Q ( new_AGEMA_signal_23988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C ( clk ), .D ( new_AGEMA_signal_23993 ), .Q ( new_AGEMA_signal_23994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C ( clk ), .D ( new_AGEMA_signal_23999 ), .Q ( new_AGEMA_signal_24000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C ( clk ), .D ( new_AGEMA_signal_24009 ), .Q ( new_AGEMA_signal_24010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C ( clk ), .D ( new_AGEMA_signal_24019 ), .Q ( new_AGEMA_signal_24020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C ( clk ), .D ( new_AGEMA_signal_24029 ), .Q ( new_AGEMA_signal_24030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C ( clk ), .D ( new_AGEMA_signal_24039 ), .Q ( new_AGEMA_signal_24040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C ( clk ), .D ( new_AGEMA_signal_24049 ), .Q ( new_AGEMA_signal_24050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C ( clk ), .D ( new_AGEMA_signal_24055 ), .Q ( new_AGEMA_signal_24056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C ( clk ), .D ( new_AGEMA_signal_24061 ), .Q ( new_AGEMA_signal_24062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C ( clk ), .D ( new_AGEMA_signal_24067 ), .Q ( new_AGEMA_signal_24068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C ( clk ), .D ( new_AGEMA_signal_24073 ), .Q ( new_AGEMA_signal_24074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C ( clk ), .D ( new_AGEMA_signal_24079 ), .Q ( new_AGEMA_signal_24080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C ( clk ), .D ( new_AGEMA_signal_24085 ), .Q ( new_AGEMA_signal_24086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C ( clk ), .D ( new_AGEMA_signal_24091 ), .Q ( new_AGEMA_signal_24092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C ( clk ), .D ( new_AGEMA_signal_24097 ), .Q ( new_AGEMA_signal_24098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C ( clk ), .D ( new_AGEMA_signal_24103 ), .Q ( new_AGEMA_signal_24104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C ( clk ), .D ( new_AGEMA_signal_24109 ), .Q ( new_AGEMA_signal_24110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C ( clk ), .D ( new_AGEMA_signal_24113 ), .Q ( new_AGEMA_signal_24114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C ( clk ), .D ( new_AGEMA_signal_24117 ), .Q ( new_AGEMA_signal_24118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C ( clk ), .D ( new_AGEMA_signal_24121 ), .Q ( new_AGEMA_signal_24122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C ( clk ), .D ( new_AGEMA_signal_24125 ), .Q ( new_AGEMA_signal_24126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C ( clk ), .D ( new_AGEMA_signal_24129 ), .Q ( new_AGEMA_signal_24130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C ( clk ), .D ( new_AGEMA_signal_24133 ), .Q ( new_AGEMA_signal_24134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C ( clk ), .D ( new_AGEMA_signal_24137 ), .Q ( new_AGEMA_signal_24138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C ( clk ), .D ( new_AGEMA_signal_24141 ), .Q ( new_AGEMA_signal_24142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7371 ( .C ( clk ), .D ( new_AGEMA_signal_24145 ), .Q ( new_AGEMA_signal_24146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C ( clk ), .D ( new_AGEMA_signal_24149 ), .Q ( new_AGEMA_signal_24150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C ( clk ), .D ( new_AGEMA_signal_24157 ), .Q ( new_AGEMA_signal_24158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C ( clk ), .D ( new_AGEMA_signal_24165 ), .Q ( new_AGEMA_signal_24166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C ( clk ), .D ( new_AGEMA_signal_24173 ), .Q ( new_AGEMA_signal_24174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C ( clk ), .D ( new_AGEMA_signal_24181 ), .Q ( new_AGEMA_signal_24182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C ( clk ), .D ( new_AGEMA_signal_24189 ), .Q ( new_AGEMA_signal_24190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C ( clk ), .D ( new_AGEMA_signal_24195 ), .Q ( new_AGEMA_signal_24196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7427 ( .C ( clk ), .D ( new_AGEMA_signal_24201 ), .Q ( new_AGEMA_signal_24202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C ( clk ), .D ( new_AGEMA_signal_24207 ), .Q ( new_AGEMA_signal_24208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C ( clk ), .D ( new_AGEMA_signal_24213 ), .Q ( new_AGEMA_signal_24214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C ( clk ), .D ( new_AGEMA_signal_24219 ), .Q ( new_AGEMA_signal_24220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C ( clk ), .D ( new_AGEMA_signal_24227 ), .Q ( new_AGEMA_signal_24228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C ( clk ), .D ( new_AGEMA_signal_24235 ), .Q ( new_AGEMA_signal_24236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C ( clk ), .D ( new_AGEMA_signal_24243 ), .Q ( new_AGEMA_signal_24244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C ( clk ), .D ( new_AGEMA_signal_24251 ), .Q ( new_AGEMA_signal_24252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C ( clk ), .D ( new_AGEMA_signal_24259 ), .Q ( new_AGEMA_signal_24260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C ( clk ), .D ( new_AGEMA_signal_24267 ), .Q ( new_AGEMA_signal_24268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C ( clk ), .D ( new_AGEMA_signal_24275 ), .Q ( new_AGEMA_signal_24276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C ( clk ), .D ( new_AGEMA_signal_24283 ), .Q ( new_AGEMA_signal_24284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C ( clk ), .D ( new_AGEMA_signal_24291 ), .Q ( new_AGEMA_signal_24292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C ( clk ), .D ( new_AGEMA_signal_24299 ), .Q ( new_AGEMA_signal_24300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_24302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C ( clk ), .D ( new_AGEMA_signal_4190 ), .Q ( new_AGEMA_signal_24304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C ( clk ), .D ( new_AGEMA_signal_4191 ), .Q ( new_AGEMA_signal_24306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C ( clk ), .D ( new_AGEMA_signal_4192 ), .Q ( new_AGEMA_signal_24308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C ( clk ), .D ( new_AGEMA_signal_4193 ), .Q ( new_AGEMA_signal_24310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C ( clk ), .D ( new_AGEMA_signal_24313 ), .Q ( new_AGEMA_signal_24314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C ( clk ), .D ( new_AGEMA_signal_24317 ), .Q ( new_AGEMA_signal_24318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C ( clk ), .D ( new_AGEMA_signal_24321 ), .Q ( new_AGEMA_signal_24322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C ( clk ), .D ( new_AGEMA_signal_24325 ), .Q ( new_AGEMA_signal_24326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C ( clk ), .D ( new_AGEMA_signal_24329 ), .Q ( new_AGEMA_signal_24330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C ( clk ), .D ( new_AGEMA_signal_24333 ), .Q ( new_AGEMA_signal_24334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C ( clk ), .D ( new_AGEMA_signal_24337 ), .Q ( new_AGEMA_signal_24338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C ( clk ), .D ( new_AGEMA_signal_24341 ), .Q ( new_AGEMA_signal_24342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C ( clk ), .D ( new_AGEMA_signal_24345 ), .Q ( new_AGEMA_signal_24346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C ( clk ), .D ( new_AGEMA_signal_24349 ), .Q ( new_AGEMA_signal_24350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C ( clk ), .D ( new_AGEMA_signal_24357 ), .Q ( new_AGEMA_signal_24358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C ( clk ), .D ( new_AGEMA_signal_24365 ), .Q ( new_AGEMA_signal_24366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C ( clk ), .D ( new_AGEMA_signal_24373 ), .Q ( new_AGEMA_signal_24374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C ( clk ), .D ( new_AGEMA_signal_24381 ), .Q ( new_AGEMA_signal_24382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C ( clk ), .D ( new_AGEMA_signal_24389 ), .Q ( new_AGEMA_signal_24390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C ( clk ), .D ( new_AGEMA_signal_24393 ), .Q ( new_AGEMA_signal_24394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C ( clk ), .D ( new_AGEMA_signal_24397 ), .Q ( new_AGEMA_signal_24398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C ( clk ), .D ( new_AGEMA_signal_24401 ), .Q ( new_AGEMA_signal_24402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C ( clk ), .D ( new_AGEMA_signal_24405 ), .Q ( new_AGEMA_signal_24406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C ( clk ), .D ( new_AGEMA_signal_24409 ), .Q ( new_AGEMA_signal_24410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C ( clk ), .D ( new_AGEMA_signal_24415 ), .Q ( new_AGEMA_signal_24416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C ( clk ), .D ( new_AGEMA_signal_24423 ), .Q ( new_AGEMA_signal_24424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C ( clk ), .D ( new_AGEMA_signal_24431 ), .Q ( new_AGEMA_signal_24432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7665 ( .C ( clk ), .D ( new_AGEMA_signal_24439 ), .Q ( new_AGEMA_signal_24440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7673 ( .C ( clk ), .D ( new_AGEMA_signal_24447 ), .Q ( new_AGEMA_signal_24448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7685 ( .C ( clk ), .D ( new_AGEMA_signal_24459 ), .Q ( new_AGEMA_signal_24460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7697 ( .C ( clk ), .D ( new_AGEMA_signal_24471 ), .Q ( new_AGEMA_signal_24472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7709 ( .C ( clk ), .D ( new_AGEMA_signal_24483 ), .Q ( new_AGEMA_signal_24484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7721 ( .C ( clk ), .D ( new_AGEMA_signal_24495 ), .Q ( new_AGEMA_signal_24496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7733 ( .C ( clk ), .D ( new_AGEMA_signal_24507 ), .Q ( new_AGEMA_signal_24508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7747 ( .C ( clk ), .D ( new_AGEMA_signal_24521 ), .Q ( new_AGEMA_signal_24522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7761 ( .C ( clk ), .D ( new_AGEMA_signal_24535 ), .Q ( new_AGEMA_signal_24536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7775 ( .C ( clk ), .D ( new_AGEMA_signal_24549 ), .Q ( new_AGEMA_signal_24550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7789 ( .C ( clk ), .D ( new_AGEMA_signal_24563 ), .Q ( new_AGEMA_signal_24564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7803 ( .C ( clk ), .D ( new_AGEMA_signal_24577 ), .Q ( new_AGEMA_signal_24578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7811 ( .C ( clk ), .D ( new_AGEMA_signal_24585 ), .Q ( new_AGEMA_signal_24586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7819 ( .C ( clk ), .D ( new_AGEMA_signal_24593 ), .Q ( new_AGEMA_signal_24594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7827 ( .C ( clk ), .D ( new_AGEMA_signal_24601 ), .Q ( new_AGEMA_signal_24602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7835 ( .C ( clk ), .D ( new_AGEMA_signal_24609 ), .Q ( new_AGEMA_signal_24610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7843 ( .C ( clk ), .D ( new_AGEMA_signal_24617 ), .Q ( new_AGEMA_signal_24618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7857 ( .C ( clk ), .D ( new_AGEMA_signal_24631 ), .Q ( new_AGEMA_signal_24632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7871 ( .C ( clk ), .D ( new_AGEMA_signal_24645 ), .Q ( new_AGEMA_signal_24646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7885 ( .C ( clk ), .D ( new_AGEMA_signal_24659 ), .Q ( new_AGEMA_signal_24660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7899 ( .C ( clk ), .D ( new_AGEMA_signal_24673 ), .Q ( new_AGEMA_signal_24674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7913 ( .C ( clk ), .D ( new_AGEMA_signal_24687 ), .Q ( new_AGEMA_signal_24688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7921 ( .C ( clk ), .D ( new_AGEMA_signal_24695 ), .Q ( new_AGEMA_signal_24696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7929 ( .C ( clk ), .D ( new_AGEMA_signal_24703 ), .Q ( new_AGEMA_signal_24704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7937 ( .C ( clk ), .D ( new_AGEMA_signal_24711 ), .Q ( new_AGEMA_signal_24712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7945 ( .C ( clk ), .D ( new_AGEMA_signal_24719 ), .Q ( new_AGEMA_signal_24720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7953 ( .C ( clk ), .D ( new_AGEMA_signal_24727 ), .Q ( new_AGEMA_signal_24728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7961 ( .C ( clk ), .D ( new_AGEMA_signal_24735 ), .Q ( new_AGEMA_signal_24736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7969 ( .C ( clk ), .D ( new_AGEMA_signal_24743 ), .Q ( new_AGEMA_signal_24744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7977 ( .C ( clk ), .D ( new_AGEMA_signal_24751 ), .Q ( new_AGEMA_signal_24752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7985 ( .C ( clk ), .D ( new_AGEMA_signal_24759 ), .Q ( new_AGEMA_signal_24760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7993 ( .C ( clk ), .D ( new_AGEMA_signal_24767 ), .Q ( new_AGEMA_signal_24768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8037 ( .C ( clk ), .D ( new_AGEMA_signal_24811 ), .Q ( new_AGEMA_signal_24812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8053 ( .C ( clk ), .D ( new_AGEMA_signal_24827 ), .Q ( new_AGEMA_signal_24828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8069 ( .C ( clk ), .D ( new_AGEMA_signal_24843 ), .Q ( new_AGEMA_signal_24844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8085 ( .C ( clk ), .D ( new_AGEMA_signal_24859 ), .Q ( new_AGEMA_signal_24860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8101 ( .C ( clk ), .D ( new_AGEMA_signal_24875 ), .Q ( new_AGEMA_signal_24876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8147 ( .C ( clk ), .D ( new_AGEMA_signal_24921 ), .Q ( new_AGEMA_signal_24922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8163 ( .C ( clk ), .D ( new_AGEMA_signal_24937 ), .Q ( new_AGEMA_signal_24938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8179 ( .C ( clk ), .D ( new_AGEMA_signal_24953 ), .Q ( new_AGEMA_signal_24954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8195 ( .C ( clk ), .D ( new_AGEMA_signal_24969 ), .Q ( new_AGEMA_signal_24970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8211 ( .C ( clk ), .D ( new_AGEMA_signal_24985 ), .Q ( new_AGEMA_signal_24986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8221 ( .C ( clk ), .D ( new_AGEMA_signal_24995 ), .Q ( new_AGEMA_signal_24996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8231 ( .C ( clk ), .D ( new_AGEMA_signal_25005 ), .Q ( new_AGEMA_signal_25006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8241 ( .C ( clk ), .D ( new_AGEMA_signal_25015 ), .Q ( new_AGEMA_signal_25016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8251 ( .C ( clk ), .D ( new_AGEMA_signal_25025 ), .Q ( new_AGEMA_signal_25026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8261 ( .C ( clk ), .D ( new_AGEMA_signal_25035 ), .Q ( new_AGEMA_signal_25036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8289 ( .C ( clk ), .D ( new_AGEMA_signal_25063 ), .Q ( new_AGEMA_signal_25064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8297 ( .C ( clk ), .D ( new_AGEMA_signal_25071 ), .Q ( new_AGEMA_signal_25072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8305 ( .C ( clk ), .D ( new_AGEMA_signal_25079 ), .Q ( new_AGEMA_signal_25080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8313 ( .C ( clk ), .D ( new_AGEMA_signal_25087 ), .Q ( new_AGEMA_signal_25088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8321 ( .C ( clk ), .D ( new_AGEMA_signal_25095 ), .Q ( new_AGEMA_signal_25096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8395 ( .C ( clk ), .D ( new_AGEMA_signal_25169 ), .Q ( new_AGEMA_signal_25170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8411 ( .C ( clk ), .D ( new_AGEMA_signal_25185 ), .Q ( new_AGEMA_signal_25186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8427 ( .C ( clk ), .D ( new_AGEMA_signal_25201 ), .Q ( new_AGEMA_signal_25202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8443 ( .C ( clk ), .D ( new_AGEMA_signal_25217 ), .Q ( new_AGEMA_signal_25218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8459 ( .C ( clk ), .D ( new_AGEMA_signal_25233 ), .Q ( new_AGEMA_signal_25234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8469 ( .C ( clk ), .D ( new_AGEMA_signal_25243 ), .Q ( new_AGEMA_signal_25244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8479 ( .C ( clk ), .D ( new_AGEMA_signal_25253 ), .Q ( new_AGEMA_signal_25254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8489 ( .C ( clk ), .D ( new_AGEMA_signal_25263 ), .Q ( new_AGEMA_signal_25264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8499 ( .C ( clk ), .D ( new_AGEMA_signal_25273 ), .Q ( new_AGEMA_signal_25274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8509 ( .C ( clk ), .D ( new_AGEMA_signal_25283 ), .Q ( new_AGEMA_signal_25284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8527 ( .C ( clk ), .D ( new_AGEMA_signal_25301 ), .Q ( new_AGEMA_signal_25302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8545 ( .C ( clk ), .D ( new_AGEMA_signal_25319 ), .Q ( new_AGEMA_signal_25320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8563 ( .C ( clk ), .D ( new_AGEMA_signal_25337 ), .Q ( new_AGEMA_signal_25338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8581 ( .C ( clk ), .D ( new_AGEMA_signal_25355 ), .Q ( new_AGEMA_signal_25356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8599 ( .C ( clk ), .D ( new_AGEMA_signal_25373 ), .Q ( new_AGEMA_signal_25374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8627 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_25402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8635 ( .C ( clk ), .D ( new_AGEMA_signal_4338 ), .Q ( new_AGEMA_signal_25410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8643 ( .C ( clk ), .D ( new_AGEMA_signal_4339 ), .Q ( new_AGEMA_signal_25418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8651 ( .C ( clk ), .D ( new_AGEMA_signal_4340 ), .Q ( new_AGEMA_signal_25426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8659 ( .C ( clk ), .D ( new_AGEMA_signal_4341 ), .Q ( new_AGEMA_signal_25434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8777 ( .C ( clk ), .D ( new_AGEMA_signal_25551 ), .Q ( new_AGEMA_signal_25552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8797 ( .C ( clk ), .D ( new_AGEMA_signal_25571 ), .Q ( new_AGEMA_signal_25572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8817 ( .C ( clk ), .D ( new_AGEMA_signal_25591 ), .Q ( new_AGEMA_signal_25592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8837 ( .C ( clk ), .D ( new_AGEMA_signal_25611 ), .Q ( new_AGEMA_signal_25612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8857 ( .C ( clk ), .D ( new_AGEMA_signal_25631 ), .Q ( new_AGEMA_signal_25632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8907 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_25682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8919 ( .C ( clk ), .D ( new_AGEMA_signal_4318 ), .Q ( new_AGEMA_signal_25694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8931 ( .C ( clk ), .D ( new_AGEMA_signal_4319 ), .Q ( new_AGEMA_signal_25706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8943 ( .C ( clk ), .D ( new_AGEMA_signal_4320 ), .Q ( new_AGEMA_signal_25718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8955 ( .C ( clk ), .D ( new_AGEMA_signal_4321 ), .Q ( new_AGEMA_signal_25730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8967 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_25742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8981 ( .C ( clk ), .D ( new_AGEMA_signal_4314 ), .Q ( new_AGEMA_signal_25756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8995 ( .C ( clk ), .D ( new_AGEMA_signal_4315 ), .Q ( new_AGEMA_signal_25770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9009 ( .C ( clk ), .D ( new_AGEMA_signal_4316 ), .Q ( new_AGEMA_signal_25784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9023 ( .C ( clk ), .D ( new_AGEMA_signal_4317 ), .Q ( new_AGEMA_signal_25798 ) ) ;

    /* cells in depth 18 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2016 ( .ina ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, new_AGEMA_signal_4251, new_AGEMA_signal_4250, n1941}), .inb ({new_AGEMA_signal_23281, new_AGEMA_signal_23275, new_AGEMA_signal_23269, new_AGEMA_signal_23263, new_AGEMA_signal_23257}), .clk ( clk ), .rnd ({Fresh[11909], Fresh[11908], Fresh[11907], Fresh[11906], Fresh[11905], Fresh[11904], Fresh[11903], Fresh[11902], Fresh[11901], Fresh[11900], Fresh[11899], Fresh[11898], Fresh[11897], Fresh[11896], Fresh[11895]}), .outt ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, new_AGEMA_signal_4363, new_AGEMA_signal_4362, n2019}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2060 ( .ina ({new_AGEMA_signal_23311, new_AGEMA_signal_23305, new_AGEMA_signal_23299, new_AGEMA_signal_23293, new_AGEMA_signal_23287}), .inb ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, new_AGEMA_signal_4254, n1960}), .clk ( clk ), .rnd ({Fresh[11924], Fresh[11923], Fresh[11922], Fresh[11921], Fresh[11920], Fresh[11919], Fresh[11918], Fresh[11917], Fresh[11916], Fresh[11915], Fresh[11914], Fresh[11913], Fresh[11912], Fresh[11911], Fresh[11910]}), .outt ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, new_AGEMA_signal_4367, new_AGEMA_signal_4366, n2002}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2116 ( .ina ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, new_AGEMA_signal_4259, new_AGEMA_signal_4258, n1988}), .inb ({new_AGEMA_signal_23341, new_AGEMA_signal_23335, new_AGEMA_signal_23329, new_AGEMA_signal_23323, new_AGEMA_signal_23317}), .clk ( clk ), .rnd ({Fresh[11939], Fresh[11938], Fresh[11937], Fresh[11936], Fresh[11935], Fresh[11934], Fresh[11933], Fresh[11932], Fresh[11931], Fresh[11930], Fresh[11929], Fresh[11928], Fresh[11927], Fresh[11926], Fresh[11925]}), .outt ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, new_AGEMA_signal_4371, new_AGEMA_signal_4370, n1989}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2154 ( .ina ({new_AGEMA_signal_23361, new_AGEMA_signal_23357, new_AGEMA_signal_23353, new_AGEMA_signal_23349, new_AGEMA_signal_23345}), .inb ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, new_AGEMA_signal_4263, new_AGEMA_signal_4262, n2015}), .clk ( clk ), .rnd ({Fresh[11954], Fresh[11953], Fresh[11952], Fresh[11951], Fresh[11950], Fresh[11949], Fresh[11948], Fresh[11947], Fresh[11946], Fresh[11945], Fresh[11944], Fresh[11943], Fresh[11942], Fresh[11941], Fresh[11940]}), .outt ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, new_AGEMA_signal_4375, new_AGEMA_signal_4374, n2016}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2170 ( .ina ({new_AGEMA_signal_23401, new_AGEMA_signal_23393, new_AGEMA_signal_23385, new_AGEMA_signal_23377, new_AGEMA_signal_23369}), .inb ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, new_AGEMA_signal_4095, new_AGEMA_signal_4094, n2030}), .clk ( clk ), .rnd ({Fresh[11969], Fresh[11968], Fresh[11967], Fresh[11966], Fresh[11965], Fresh[11964], Fresh[11963], Fresh[11962], Fresh[11961], Fresh[11960], Fresh[11959], Fresh[11958], Fresh[11957], Fresh[11956], Fresh[11955]}), .outt ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, new_AGEMA_signal_4266, n2038}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2201 ( .ina ({new_AGEMA_signal_23431, new_AGEMA_signal_23425, new_AGEMA_signal_23419, new_AGEMA_signal_23413, new_AGEMA_signal_23407}), .inb ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, new_AGEMA_signal_4271, new_AGEMA_signal_4270, n2053}), .clk ( clk ), .rnd ({Fresh[11984], Fresh[11983], Fresh[11982], Fresh[11981], Fresh[11980], Fresh[11979], Fresh[11978], Fresh[11977], Fresh[11976], Fresh[11975], Fresh[11974], Fresh[11973], Fresh[11972], Fresh[11971], Fresh[11970]}), .outt ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, new_AGEMA_signal_4383, new_AGEMA_signal_4382, n2111}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2223 ( .ina ({new_AGEMA_signal_23451, new_AGEMA_signal_23447, new_AGEMA_signal_23443, new_AGEMA_signal_23439, new_AGEMA_signal_23435}), .inb ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, new_AGEMA_signal_4275, new_AGEMA_signal_4274, n2071}), .clk ( clk ), .rnd ({Fresh[11999], Fresh[11998], Fresh[11997], Fresh[11996], Fresh[11995], Fresh[11994], Fresh[11993], Fresh[11992], Fresh[11991], Fresh[11990], Fresh[11989], Fresh[11988], Fresh[11987], Fresh[11986], Fresh[11985]}), .outt ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, new_AGEMA_signal_4386, n2079}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2263 ( .ina ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, new_AGEMA_signal_4278, n2103}), .inb ({new_AGEMA_signal_23491, new_AGEMA_signal_23483, new_AGEMA_signal_23475, new_AGEMA_signal_23467, new_AGEMA_signal_23459}), .clk ( clk ), .rnd ({Fresh[12014], Fresh[12013], Fresh[12012], Fresh[12011], Fresh[12010], Fresh[12009], Fresh[12008], Fresh[12007], Fresh[12006], Fresh[12005], Fresh[12004], Fresh[12003], Fresh[12002], Fresh[12001], Fresh[12000]}), .outt ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, new_AGEMA_signal_4391, new_AGEMA_signal_4390, n2104}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2289 ( .ina ({new_AGEMA_signal_23531, new_AGEMA_signal_23523, new_AGEMA_signal_23515, new_AGEMA_signal_23507, new_AGEMA_signal_23499}), .inb ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, new_AGEMA_signal_4283, new_AGEMA_signal_4282, n2126}), .clk ( clk ), .rnd ({Fresh[12029], Fresh[12028], Fresh[12027], Fresh[12026], Fresh[12025], Fresh[12024], Fresh[12023], Fresh[12022], Fresh[12021], Fresh[12020], Fresh[12019], Fresh[12018], Fresh[12017], Fresh[12016], Fresh[12015]}), .outt ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, new_AGEMA_signal_4395, new_AGEMA_signal_4394, n2127}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2315 ( .ina ({new_AGEMA_signal_23361, new_AGEMA_signal_23357, new_AGEMA_signal_23353, new_AGEMA_signal_23349, new_AGEMA_signal_23345}), .inb ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, new_AGEMA_signal_4287, new_AGEMA_signal_4286, n2146}), .clk ( clk ), .rnd ({Fresh[12044], Fresh[12043], Fresh[12042], Fresh[12041], Fresh[12040], Fresh[12039], Fresh[12038], Fresh[12037], Fresh[12036], Fresh[12035], Fresh[12034], Fresh[12033], Fresh[12032], Fresh[12031], Fresh[12030]}), .outt ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, new_AGEMA_signal_4398, n2147}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2336 ( .ina ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, new_AGEMA_signal_4290, n2173}), .inb ({new_AGEMA_signal_23581, new_AGEMA_signal_23571, new_AGEMA_signal_23561, new_AGEMA_signal_23551, new_AGEMA_signal_23541}), .clk ( clk ), .rnd ({Fresh[12059], Fresh[12058], Fresh[12057], Fresh[12056], Fresh[12055], Fresh[12054], Fresh[12053], Fresh[12052], Fresh[12051], Fresh[12050], Fresh[12049], Fresh[12048], Fresh[12047], Fresh[12046], Fresh[12045]}), .outt ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, new_AGEMA_signal_4403, new_AGEMA_signal_4402, n2208}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2352 ( .ina ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, new_AGEMA_signal_4295, new_AGEMA_signal_4294, n2187}), .inb ({new_AGEMA_signal_23621, new_AGEMA_signal_23613, new_AGEMA_signal_23605, new_AGEMA_signal_23597, new_AGEMA_signal_23589}), .clk ( clk ), .rnd ({Fresh[12074], Fresh[12073], Fresh[12072], Fresh[12071], Fresh[12070], Fresh[12069], Fresh[12068], Fresh[12067], Fresh[12066], Fresh[12065], Fresh[12064], Fresh[12063], Fresh[12062], Fresh[12061], Fresh[12060]}), .outt ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, new_AGEMA_signal_4407, new_AGEMA_signal_4406, n2199}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2420 ( .ina ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, new_AGEMA_signal_4302, n2256}), .inb ({new_AGEMA_signal_23651, new_AGEMA_signal_23645, new_AGEMA_signal_23639, new_AGEMA_signal_23633, new_AGEMA_signal_23627}), .clk ( clk ), .rnd ({Fresh[12089], Fresh[12088], Fresh[12087], Fresh[12086], Fresh[12085], Fresh[12084], Fresh[12083], Fresh[12082], Fresh[12081], Fresh[12080], Fresh[12079], Fresh[12078], Fresh[12077], Fresh[12076], Fresh[12075]}), .outt ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, new_AGEMA_signal_4410, n2257}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2442 ( .ina ({new_AGEMA_signal_23671, new_AGEMA_signal_23667, new_AGEMA_signal_23663, new_AGEMA_signal_23659, new_AGEMA_signal_23655}), .inb ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, new_AGEMA_signal_4307, new_AGEMA_signal_4306, n2275}), .clk ( clk ), .rnd ({Fresh[12104], Fresh[12103], Fresh[12102], Fresh[12101], Fresh[12100], Fresh[12099], Fresh[12098], Fresh[12097], Fresh[12096], Fresh[12095], Fresh[12094], Fresh[12093], Fresh[12092], Fresh[12091], Fresh[12090]}), .outt ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, new_AGEMA_signal_4415, new_AGEMA_signal_4414, n2281}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2475 ( .ina ({new_AGEMA_signal_23701, new_AGEMA_signal_23695, new_AGEMA_signal_23689, new_AGEMA_signal_23683, new_AGEMA_signal_23677}), .inb ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, new_AGEMA_signal_4311, new_AGEMA_signal_4310, n2303}), .clk ( clk ), .rnd ({Fresh[12119], Fresh[12118], Fresh[12117], Fresh[12116], Fresh[12115], Fresh[12114], Fresh[12113], Fresh[12112], Fresh[12111], Fresh[12110], Fresh[12109], Fresh[12108], Fresh[12107], Fresh[12106], Fresh[12105]}), .outt ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, new_AGEMA_signal_4419, new_AGEMA_signal_4418, n2305}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2532 ( .ina ({new_AGEMA_signal_23741, new_AGEMA_signal_23733, new_AGEMA_signal_23725, new_AGEMA_signal_23717, new_AGEMA_signal_23709}), .inb ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, new_AGEMA_signal_4323, new_AGEMA_signal_4322, n2366}), .clk ( clk ), .rnd ({Fresh[12134], Fresh[12133], Fresh[12132], Fresh[12131], Fresh[12130], Fresh[12129], Fresh[12128], Fresh[12127], Fresh[12126], Fresh[12125], Fresh[12124], Fresh[12123], Fresh[12122], Fresh[12121], Fresh[12120]}), .outt ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, new_AGEMA_signal_4423, new_AGEMA_signal_4422, n2368}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2583 ( .ina ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, new_AGEMA_signal_4326, n2425}), .inb ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, new_AGEMA_signal_4182, n2424}), .clk ( clk ), .rnd ({Fresh[12149], Fresh[12148], Fresh[12147], Fresh[12146], Fresh[12145], Fresh[12144], Fresh[12143], Fresh[12142], Fresh[12141], Fresh[12140], Fresh[12139], Fresh[12138], Fresh[12137], Fresh[12136], Fresh[12135]}), .outt ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, new_AGEMA_signal_4427, new_AGEMA_signal_4426, n2426}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2605 ( .ina ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, new_AGEMA_signal_4331, new_AGEMA_signal_4330, n2451}), .inb ({new_AGEMA_signal_23771, new_AGEMA_signal_23765, new_AGEMA_signal_23759, new_AGEMA_signal_23753, new_AGEMA_signal_23747}), .clk ( clk ), .rnd ({Fresh[12164], Fresh[12163], Fresh[12162], Fresh[12161], Fresh[12160], Fresh[12159], Fresh[12158], Fresh[12157], Fresh[12156], Fresh[12155], Fresh[12154], Fresh[12153], Fresh[12152], Fresh[12151], Fresh[12150]}), .outt ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, new_AGEMA_signal_4431, new_AGEMA_signal_4430, n2457}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2659 ( .ina ({new_AGEMA_signal_23781, new_AGEMA_signal_23779, new_AGEMA_signal_23777, new_AGEMA_signal_23775, new_AGEMA_signal_23773}), .inb ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, new_AGEMA_signal_4335, new_AGEMA_signal_4334, n2511}), .clk ( clk ), .rnd ({Fresh[12179], Fresh[12178], Fresh[12177], Fresh[12176], Fresh[12175], Fresh[12174], Fresh[12173], Fresh[12172], Fresh[12171], Fresh[12170], Fresh[12169], Fresh[12168], Fresh[12167], Fresh[12166], Fresh[12165]}), .outt ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, new_AGEMA_signal_4435, new_AGEMA_signal_4434, n2513}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2717 ( .ina ({new_AGEMA_signal_23821, new_AGEMA_signal_23813, new_AGEMA_signal_23805, new_AGEMA_signal_23797, new_AGEMA_signal_23789}), .inb ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, new_AGEMA_signal_4343, new_AGEMA_signal_4342, n2590}), .clk ( clk ), .rnd ({Fresh[12194], Fresh[12193], Fresh[12192], Fresh[12191], Fresh[12190], Fresh[12189], Fresh[12188], Fresh[12187], Fresh[12186], Fresh[12185], Fresh[12184], Fresh[12183], Fresh[12182], Fresh[12181], Fresh[12180]}), .outt ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, new_AGEMA_signal_4439, new_AGEMA_signal_4438, n2592}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2741 ( .ina ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, new_AGEMA_signal_4223, new_AGEMA_signal_4222, n2623}), .inb ({new_AGEMA_signal_23841, new_AGEMA_signal_23837, new_AGEMA_signal_23833, new_AGEMA_signal_23829, new_AGEMA_signal_23825}), .clk ( clk ), .rnd ({Fresh[12209], Fresh[12208], Fresh[12207], Fresh[12206], Fresh[12205], Fresh[12204], Fresh[12203], Fresh[12202], Fresh[12201], Fresh[12200], Fresh[12199], Fresh[12198], Fresh[12197], Fresh[12196], Fresh[12195]}), .outt ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, n2637}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2767 ( .ina ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, new_AGEMA_signal_4350, n2667}), .inb ({new_AGEMA_signal_23871, new_AGEMA_signal_23865, new_AGEMA_signal_23859, new_AGEMA_signal_23853, new_AGEMA_signal_23847}), .clk ( clk ), .rnd ({Fresh[12224], Fresh[12223], Fresh[12222], Fresh[12221], Fresh[12220], Fresh[12219], Fresh[12218], Fresh[12217], Fresh[12216], Fresh[12215], Fresh[12214], Fresh[12213], Fresh[12212], Fresh[12211], Fresh[12210]}), .outt ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, new_AGEMA_signal_4447, new_AGEMA_signal_4446, n2668}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2787 ( .ina ({new_AGEMA_signal_23901, new_AGEMA_signal_23895, new_AGEMA_signal_23889, new_AGEMA_signal_23883, new_AGEMA_signal_23877}), .inb ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, new_AGEMA_signal_4355, new_AGEMA_signal_4354, n2703}), .clk ( clk ), .rnd ({Fresh[12239], Fresh[12238], Fresh[12237], Fresh[12236], Fresh[12235], Fresh[12234], Fresh[12233], Fresh[12232], Fresh[12231], Fresh[12230], Fresh[12229], Fresh[12228], Fresh[12227], Fresh[12226], Fresh[12225]}), .outt ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, n2705}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2841 ( .ina ({new_AGEMA_signal_23921, new_AGEMA_signal_23917, new_AGEMA_signal_23913, new_AGEMA_signal_23909, new_AGEMA_signal_23905}), .inb ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, new_AGEMA_signal_4242, n2803}), .clk ( clk ), .rnd ({Fresh[12254], Fresh[12253], Fresh[12252], Fresh[12251], Fresh[12250], Fresh[12249], Fresh[12248], Fresh[12247], Fresh[12246], Fresh[12245], Fresh[12244], Fresh[12243], Fresh[12242], Fresh[12241], Fresh[12240]}), .outt ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, new_AGEMA_signal_4359, new_AGEMA_signal_4358, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C ( clk ), .D ( new_AGEMA_signal_23926 ), .Q ( new_AGEMA_signal_23927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C ( clk ), .D ( new_AGEMA_signal_23932 ), .Q ( new_AGEMA_signal_23933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C ( clk ), .D ( new_AGEMA_signal_23938 ), .Q ( new_AGEMA_signal_23939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C ( clk ), .D ( new_AGEMA_signal_23944 ), .Q ( new_AGEMA_signal_23945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C ( clk ), .D ( new_AGEMA_signal_23950 ), .Q ( new_AGEMA_signal_23951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C ( clk ), .D ( new_AGEMA_signal_23954 ), .Q ( new_AGEMA_signal_23955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C ( clk ), .D ( new_AGEMA_signal_23958 ), .Q ( new_AGEMA_signal_23959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C ( clk ), .D ( new_AGEMA_signal_23962 ), .Q ( new_AGEMA_signal_23963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C ( clk ), .D ( new_AGEMA_signal_23966 ), .Q ( new_AGEMA_signal_23967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C ( clk ), .D ( new_AGEMA_signal_23970 ), .Q ( new_AGEMA_signal_23971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C ( clk ), .D ( new_AGEMA_signal_23976 ), .Q ( new_AGEMA_signal_23977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C ( clk ), .D ( new_AGEMA_signal_23982 ), .Q ( new_AGEMA_signal_23983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C ( clk ), .D ( new_AGEMA_signal_23988 ), .Q ( new_AGEMA_signal_23989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C ( clk ), .D ( new_AGEMA_signal_23994 ), .Q ( new_AGEMA_signal_23995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C ( clk ), .D ( new_AGEMA_signal_24000 ), .Q ( new_AGEMA_signal_24001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C ( clk ), .D ( new_AGEMA_signal_24010 ), .Q ( new_AGEMA_signal_24011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C ( clk ), .D ( new_AGEMA_signal_24020 ), .Q ( new_AGEMA_signal_24021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C ( clk ), .D ( new_AGEMA_signal_24030 ), .Q ( new_AGEMA_signal_24031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C ( clk ), .D ( new_AGEMA_signal_24040 ), .Q ( new_AGEMA_signal_24041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C ( clk ), .D ( new_AGEMA_signal_24050 ), .Q ( new_AGEMA_signal_24051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C ( clk ), .D ( new_AGEMA_signal_24056 ), .Q ( new_AGEMA_signal_24057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C ( clk ), .D ( new_AGEMA_signal_24062 ), .Q ( new_AGEMA_signal_24063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C ( clk ), .D ( new_AGEMA_signal_24068 ), .Q ( new_AGEMA_signal_24069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C ( clk ), .D ( new_AGEMA_signal_24074 ), .Q ( new_AGEMA_signal_24075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C ( clk ), .D ( new_AGEMA_signal_24080 ), .Q ( new_AGEMA_signal_24081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C ( clk ), .D ( new_AGEMA_signal_24086 ), .Q ( new_AGEMA_signal_24087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C ( clk ), .D ( new_AGEMA_signal_24092 ), .Q ( new_AGEMA_signal_24093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C ( clk ), .D ( new_AGEMA_signal_24098 ), .Q ( new_AGEMA_signal_24099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C ( clk ), .D ( new_AGEMA_signal_24104 ), .Q ( new_AGEMA_signal_24105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C ( clk ), .D ( new_AGEMA_signal_24110 ), .Q ( new_AGEMA_signal_24111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C ( clk ), .D ( new_AGEMA_signal_24114 ), .Q ( new_AGEMA_signal_24115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C ( clk ), .D ( new_AGEMA_signal_24118 ), .Q ( new_AGEMA_signal_24119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C ( clk ), .D ( new_AGEMA_signal_24122 ), .Q ( new_AGEMA_signal_24123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C ( clk ), .D ( new_AGEMA_signal_24126 ), .Q ( new_AGEMA_signal_24127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C ( clk ), .D ( new_AGEMA_signal_24130 ), .Q ( new_AGEMA_signal_24131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C ( clk ), .D ( new_AGEMA_signal_24134 ), .Q ( new_AGEMA_signal_24135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C ( clk ), .D ( new_AGEMA_signal_24138 ), .Q ( new_AGEMA_signal_24139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C ( clk ), .D ( new_AGEMA_signal_24142 ), .Q ( new_AGEMA_signal_24143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C ( clk ), .D ( new_AGEMA_signal_24146 ), .Q ( new_AGEMA_signal_24147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C ( clk ), .D ( new_AGEMA_signal_24150 ), .Q ( new_AGEMA_signal_24151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C ( clk ), .D ( new_AGEMA_signal_24158 ), .Q ( new_AGEMA_signal_24159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C ( clk ), .D ( new_AGEMA_signal_24166 ), .Q ( new_AGEMA_signal_24167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C ( clk ), .D ( new_AGEMA_signal_24174 ), .Q ( new_AGEMA_signal_24175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C ( clk ), .D ( new_AGEMA_signal_24182 ), .Q ( new_AGEMA_signal_24183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C ( clk ), .D ( new_AGEMA_signal_24190 ), .Q ( new_AGEMA_signal_24191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C ( clk ), .D ( new_AGEMA_signal_24196 ), .Q ( new_AGEMA_signal_24197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C ( clk ), .D ( new_AGEMA_signal_24202 ), .Q ( new_AGEMA_signal_24203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C ( clk ), .D ( new_AGEMA_signal_24208 ), .Q ( new_AGEMA_signal_24209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C ( clk ), .D ( new_AGEMA_signal_24214 ), .Q ( new_AGEMA_signal_24215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C ( clk ), .D ( new_AGEMA_signal_24220 ), .Q ( new_AGEMA_signal_24221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C ( clk ), .D ( new_AGEMA_signal_24228 ), .Q ( new_AGEMA_signal_24229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C ( clk ), .D ( new_AGEMA_signal_24236 ), .Q ( new_AGEMA_signal_24237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C ( clk ), .D ( new_AGEMA_signal_24244 ), .Q ( new_AGEMA_signal_24245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C ( clk ), .D ( new_AGEMA_signal_24252 ), .Q ( new_AGEMA_signal_24253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C ( clk ), .D ( new_AGEMA_signal_24260 ), .Q ( new_AGEMA_signal_24261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C ( clk ), .D ( new_AGEMA_signal_24268 ), .Q ( new_AGEMA_signal_24269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C ( clk ), .D ( new_AGEMA_signal_24276 ), .Q ( new_AGEMA_signal_24277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C ( clk ), .D ( new_AGEMA_signal_24284 ), .Q ( new_AGEMA_signal_24285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C ( clk ), .D ( new_AGEMA_signal_24292 ), .Q ( new_AGEMA_signal_24293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C ( clk ), .D ( new_AGEMA_signal_24300 ), .Q ( new_AGEMA_signal_24301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C ( clk ), .D ( new_AGEMA_signal_24302 ), .Q ( new_AGEMA_signal_24303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C ( clk ), .D ( new_AGEMA_signal_24304 ), .Q ( new_AGEMA_signal_24305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C ( clk ), .D ( new_AGEMA_signal_24306 ), .Q ( new_AGEMA_signal_24307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C ( clk ), .D ( new_AGEMA_signal_24308 ), .Q ( new_AGEMA_signal_24309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C ( clk ), .D ( new_AGEMA_signal_24310 ), .Q ( new_AGEMA_signal_24311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C ( clk ), .D ( new_AGEMA_signal_24314 ), .Q ( new_AGEMA_signal_24315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C ( clk ), .D ( new_AGEMA_signal_24318 ), .Q ( new_AGEMA_signal_24319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C ( clk ), .D ( new_AGEMA_signal_24322 ), .Q ( new_AGEMA_signal_24323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C ( clk ), .D ( new_AGEMA_signal_24326 ), .Q ( new_AGEMA_signal_24327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C ( clk ), .D ( new_AGEMA_signal_24330 ), .Q ( new_AGEMA_signal_24331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C ( clk ), .D ( new_AGEMA_signal_24334 ), .Q ( new_AGEMA_signal_24335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C ( clk ), .D ( new_AGEMA_signal_24338 ), .Q ( new_AGEMA_signal_24339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C ( clk ), .D ( new_AGEMA_signal_24342 ), .Q ( new_AGEMA_signal_24343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C ( clk ), .D ( new_AGEMA_signal_24346 ), .Q ( new_AGEMA_signal_24347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C ( clk ), .D ( new_AGEMA_signal_24350 ), .Q ( new_AGEMA_signal_24351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C ( clk ), .D ( new_AGEMA_signal_24358 ), .Q ( new_AGEMA_signal_24359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C ( clk ), .D ( new_AGEMA_signal_24366 ), .Q ( new_AGEMA_signal_24367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C ( clk ), .D ( new_AGEMA_signal_24374 ), .Q ( new_AGEMA_signal_24375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C ( clk ), .D ( new_AGEMA_signal_24382 ), .Q ( new_AGEMA_signal_24383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C ( clk ), .D ( new_AGEMA_signal_24390 ), .Q ( new_AGEMA_signal_24391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C ( clk ), .D ( new_AGEMA_signal_24394 ), .Q ( new_AGEMA_signal_24395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C ( clk ), .D ( new_AGEMA_signal_24398 ), .Q ( new_AGEMA_signal_24399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C ( clk ), .D ( new_AGEMA_signal_24402 ), .Q ( new_AGEMA_signal_24403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C ( clk ), .D ( new_AGEMA_signal_24406 ), .Q ( new_AGEMA_signal_24407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C ( clk ), .D ( new_AGEMA_signal_24410 ), .Q ( new_AGEMA_signal_24411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C ( clk ), .D ( new_AGEMA_signal_24416 ), .Q ( new_AGEMA_signal_24417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C ( clk ), .D ( new_AGEMA_signal_24424 ), .Q ( new_AGEMA_signal_24425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C ( clk ), .D ( new_AGEMA_signal_24432 ), .Q ( new_AGEMA_signal_24433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7666 ( .C ( clk ), .D ( new_AGEMA_signal_24440 ), .Q ( new_AGEMA_signal_24441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7674 ( .C ( clk ), .D ( new_AGEMA_signal_24448 ), .Q ( new_AGEMA_signal_24449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7686 ( .C ( clk ), .D ( new_AGEMA_signal_24460 ), .Q ( new_AGEMA_signal_24461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7698 ( .C ( clk ), .D ( new_AGEMA_signal_24472 ), .Q ( new_AGEMA_signal_24473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7710 ( .C ( clk ), .D ( new_AGEMA_signal_24484 ), .Q ( new_AGEMA_signal_24485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7722 ( .C ( clk ), .D ( new_AGEMA_signal_24496 ), .Q ( new_AGEMA_signal_24497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7734 ( .C ( clk ), .D ( new_AGEMA_signal_24508 ), .Q ( new_AGEMA_signal_24509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7748 ( .C ( clk ), .D ( new_AGEMA_signal_24522 ), .Q ( new_AGEMA_signal_24523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7762 ( .C ( clk ), .D ( new_AGEMA_signal_24536 ), .Q ( new_AGEMA_signal_24537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7776 ( .C ( clk ), .D ( new_AGEMA_signal_24550 ), .Q ( new_AGEMA_signal_24551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7790 ( .C ( clk ), .D ( new_AGEMA_signal_24564 ), .Q ( new_AGEMA_signal_24565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7804 ( .C ( clk ), .D ( new_AGEMA_signal_24578 ), .Q ( new_AGEMA_signal_24579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7812 ( .C ( clk ), .D ( new_AGEMA_signal_24586 ), .Q ( new_AGEMA_signal_24587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7820 ( .C ( clk ), .D ( new_AGEMA_signal_24594 ), .Q ( new_AGEMA_signal_24595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7828 ( .C ( clk ), .D ( new_AGEMA_signal_24602 ), .Q ( new_AGEMA_signal_24603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7836 ( .C ( clk ), .D ( new_AGEMA_signal_24610 ), .Q ( new_AGEMA_signal_24611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7844 ( .C ( clk ), .D ( new_AGEMA_signal_24618 ), .Q ( new_AGEMA_signal_24619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7858 ( .C ( clk ), .D ( new_AGEMA_signal_24632 ), .Q ( new_AGEMA_signal_24633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7872 ( .C ( clk ), .D ( new_AGEMA_signal_24646 ), .Q ( new_AGEMA_signal_24647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7886 ( .C ( clk ), .D ( new_AGEMA_signal_24660 ), .Q ( new_AGEMA_signal_24661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7900 ( .C ( clk ), .D ( new_AGEMA_signal_24674 ), .Q ( new_AGEMA_signal_24675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7914 ( .C ( clk ), .D ( new_AGEMA_signal_24688 ), .Q ( new_AGEMA_signal_24689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7922 ( .C ( clk ), .D ( new_AGEMA_signal_24696 ), .Q ( new_AGEMA_signal_24697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7930 ( .C ( clk ), .D ( new_AGEMA_signal_24704 ), .Q ( new_AGEMA_signal_24705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7938 ( .C ( clk ), .D ( new_AGEMA_signal_24712 ), .Q ( new_AGEMA_signal_24713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7946 ( .C ( clk ), .D ( new_AGEMA_signal_24720 ), .Q ( new_AGEMA_signal_24721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7954 ( .C ( clk ), .D ( new_AGEMA_signal_24728 ), .Q ( new_AGEMA_signal_24729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7962 ( .C ( clk ), .D ( new_AGEMA_signal_24736 ), .Q ( new_AGEMA_signal_24737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7970 ( .C ( clk ), .D ( new_AGEMA_signal_24744 ), .Q ( new_AGEMA_signal_24745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7978 ( .C ( clk ), .D ( new_AGEMA_signal_24752 ), .Q ( new_AGEMA_signal_24753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7986 ( .C ( clk ), .D ( new_AGEMA_signal_24760 ), .Q ( new_AGEMA_signal_24761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7994 ( .C ( clk ), .D ( new_AGEMA_signal_24768 ), .Q ( new_AGEMA_signal_24769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8038 ( .C ( clk ), .D ( new_AGEMA_signal_24812 ), .Q ( new_AGEMA_signal_24813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8054 ( .C ( clk ), .D ( new_AGEMA_signal_24828 ), .Q ( new_AGEMA_signal_24829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8070 ( .C ( clk ), .D ( new_AGEMA_signal_24844 ), .Q ( new_AGEMA_signal_24845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8086 ( .C ( clk ), .D ( new_AGEMA_signal_24860 ), .Q ( new_AGEMA_signal_24861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8102 ( .C ( clk ), .D ( new_AGEMA_signal_24876 ), .Q ( new_AGEMA_signal_24877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8148 ( .C ( clk ), .D ( new_AGEMA_signal_24922 ), .Q ( new_AGEMA_signal_24923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8164 ( .C ( clk ), .D ( new_AGEMA_signal_24938 ), .Q ( new_AGEMA_signal_24939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8180 ( .C ( clk ), .D ( new_AGEMA_signal_24954 ), .Q ( new_AGEMA_signal_24955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8196 ( .C ( clk ), .D ( new_AGEMA_signal_24970 ), .Q ( new_AGEMA_signal_24971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8212 ( .C ( clk ), .D ( new_AGEMA_signal_24986 ), .Q ( new_AGEMA_signal_24987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8222 ( .C ( clk ), .D ( new_AGEMA_signal_24996 ), .Q ( new_AGEMA_signal_24997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8232 ( .C ( clk ), .D ( new_AGEMA_signal_25006 ), .Q ( new_AGEMA_signal_25007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8242 ( .C ( clk ), .D ( new_AGEMA_signal_25016 ), .Q ( new_AGEMA_signal_25017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8252 ( .C ( clk ), .D ( new_AGEMA_signal_25026 ), .Q ( new_AGEMA_signal_25027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8262 ( .C ( clk ), .D ( new_AGEMA_signal_25036 ), .Q ( new_AGEMA_signal_25037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8290 ( .C ( clk ), .D ( new_AGEMA_signal_25064 ), .Q ( new_AGEMA_signal_25065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8298 ( .C ( clk ), .D ( new_AGEMA_signal_25072 ), .Q ( new_AGEMA_signal_25073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8306 ( .C ( clk ), .D ( new_AGEMA_signal_25080 ), .Q ( new_AGEMA_signal_25081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8314 ( .C ( clk ), .D ( new_AGEMA_signal_25088 ), .Q ( new_AGEMA_signal_25089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8322 ( .C ( clk ), .D ( new_AGEMA_signal_25096 ), .Q ( new_AGEMA_signal_25097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8396 ( .C ( clk ), .D ( new_AGEMA_signal_25170 ), .Q ( new_AGEMA_signal_25171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8412 ( .C ( clk ), .D ( new_AGEMA_signal_25186 ), .Q ( new_AGEMA_signal_25187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8428 ( .C ( clk ), .D ( new_AGEMA_signal_25202 ), .Q ( new_AGEMA_signal_25203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8444 ( .C ( clk ), .D ( new_AGEMA_signal_25218 ), .Q ( new_AGEMA_signal_25219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8460 ( .C ( clk ), .D ( new_AGEMA_signal_25234 ), .Q ( new_AGEMA_signal_25235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8470 ( .C ( clk ), .D ( new_AGEMA_signal_25244 ), .Q ( new_AGEMA_signal_25245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8480 ( .C ( clk ), .D ( new_AGEMA_signal_25254 ), .Q ( new_AGEMA_signal_25255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8490 ( .C ( clk ), .D ( new_AGEMA_signal_25264 ), .Q ( new_AGEMA_signal_25265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8500 ( .C ( clk ), .D ( new_AGEMA_signal_25274 ), .Q ( new_AGEMA_signal_25275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8510 ( .C ( clk ), .D ( new_AGEMA_signal_25284 ), .Q ( new_AGEMA_signal_25285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8528 ( .C ( clk ), .D ( new_AGEMA_signal_25302 ), .Q ( new_AGEMA_signal_25303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8546 ( .C ( clk ), .D ( new_AGEMA_signal_25320 ), .Q ( new_AGEMA_signal_25321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8564 ( .C ( clk ), .D ( new_AGEMA_signal_25338 ), .Q ( new_AGEMA_signal_25339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8582 ( .C ( clk ), .D ( new_AGEMA_signal_25356 ), .Q ( new_AGEMA_signal_25357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8600 ( .C ( clk ), .D ( new_AGEMA_signal_25374 ), .Q ( new_AGEMA_signal_25375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8628 ( .C ( clk ), .D ( new_AGEMA_signal_25402 ), .Q ( new_AGEMA_signal_25403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8636 ( .C ( clk ), .D ( new_AGEMA_signal_25410 ), .Q ( new_AGEMA_signal_25411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8644 ( .C ( clk ), .D ( new_AGEMA_signal_25418 ), .Q ( new_AGEMA_signal_25419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8652 ( .C ( clk ), .D ( new_AGEMA_signal_25426 ), .Q ( new_AGEMA_signal_25427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8660 ( .C ( clk ), .D ( new_AGEMA_signal_25434 ), .Q ( new_AGEMA_signal_25435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8778 ( .C ( clk ), .D ( new_AGEMA_signal_25552 ), .Q ( new_AGEMA_signal_25553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8798 ( .C ( clk ), .D ( new_AGEMA_signal_25572 ), .Q ( new_AGEMA_signal_25573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8818 ( .C ( clk ), .D ( new_AGEMA_signal_25592 ), .Q ( new_AGEMA_signal_25593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8838 ( .C ( clk ), .D ( new_AGEMA_signal_25612 ), .Q ( new_AGEMA_signal_25613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8858 ( .C ( clk ), .D ( new_AGEMA_signal_25632 ), .Q ( new_AGEMA_signal_25633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8908 ( .C ( clk ), .D ( new_AGEMA_signal_25682 ), .Q ( new_AGEMA_signal_25683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8920 ( .C ( clk ), .D ( new_AGEMA_signal_25694 ), .Q ( new_AGEMA_signal_25695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8932 ( .C ( clk ), .D ( new_AGEMA_signal_25706 ), .Q ( new_AGEMA_signal_25707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8944 ( .C ( clk ), .D ( new_AGEMA_signal_25718 ), .Q ( new_AGEMA_signal_25719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8956 ( .C ( clk ), .D ( new_AGEMA_signal_25730 ), .Q ( new_AGEMA_signal_25731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8968 ( .C ( clk ), .D ( new_AGEMA_signal_25742 ), .Q ( new_AGEMA_signal_25743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8982 ( .C ( clk ), .D ( new_AGEMA_signal_25756 ), .Q ( new_AGEMA_signal_25757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8996 ( .C ( clk ), .D ( new_AGEMA_signal_25770 ), .Q ( new_AGEMA_signal_25771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9010 ( .C ( clk ), .D ( new_AGEMA_signal_25784 ), .Q ( new_AGEMA_signal_25785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9024 ( .C ( clk ), .D ( new_AGEMA_signal_25798 ), .Q ( new_AGEMA_signal_25799 ) ) ;

    /* cells in depth 19 */
    buf_clk new_AGEMA_reg_buffer_7643 ( .C ( clk ), .D ( new_AGEMA_signal_24417 ), .Q ( new_AGEMA_signal_24418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C ( clk ), .D ( new_AGEMA_signal_24425 ), .Q ( new_AGEMA_signal_24426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C ( clk ), .D ( new_AGEMA_signal_24433 ), .Q ( new_AGEMA_signal_24434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7667 ( .C ( clk ), .D ( new_AGEMA_signal_24441 ), .Q ( new_AGEMA_signal_24442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7675 ( .C ( clk ), .D ( new_AGEMA_signal_24449 ), .Q ( new_AGEMA_signal_24450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7687 ( .C ( clk ), .D ( new_AGEMA_signal_24461 ), .Q ( new_AGEMA_signal_24462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7699 ( .C ( clk ), .D ( new_AGEMA_signal_24473 ), .Q ( new_AGEMA_signal_24474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7711 ( .C ( clk ), .D ( new_AGEMA_signal_24485 ), .Q ( new_AGEMA_signal_24486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7723 ( .C ( clk ), .D ( new_AGEMA_signal_24497 ), .Q ( new_AGEMA_signal_24498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7735 ( .C ( clk ), .D ( new_AGEMA_signal_24509 ), .Q ( new_AGEMA_signal_24510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7749 ( .C ( clk ), .D ( new_AGEMA_signal_24523 ), .Q ( new_AGEMA_signal_24524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7763 ( .C ( clk ), .D ( new_AGEMA_signal_24537 ), .Q ( new_AGEMA_signal_24538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7777 ( .C ( clk ), .D ( new_AGEMA_signal_24551 ), .Q ( new_AGEMA_signal_24552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7791 ( .C ( clk ), .D ( new_AGEMA_signal_24565 ), .Q ( new_AGEMA_signal_24566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7805 ( .C ( clk ), .D ( new_AGEMA_signal_24579 ), .Q ( new_AGEMA_signal_24580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7813 ( .C ( clk ), .D ( new_AGEMA_signal_24587 ), .Q ( new_AGEMA_signal_24588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7821 ( .C ( clk ), .D ( new_AGEMA_signal_24595 ), .Q ( new_AGEMA_signal_24596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7829 ( .C ( clk ), .D ( new_AGEMA_signal_24603 ), .Q ( new_AGEMA_signal_24604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7837 ( .C ( clk ), .D ( new_AGEMA_signal_24611 ), .Q ( new_AGEMA_signal_24612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7845 ( .C ( clk ), .D ( new_AGEMA_signal_24619 ), .Q ( new_AGEMA_signal_24620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7859 ( .C ( clk ), .D ( new_AGEMA_signal_24633 ), .Q ( new_AGEMA_signal_24634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7873 ( .C ( clk ), .D ( new_AGEMA_signal_24647 ), .Q ( new_AGEMA_signal_24648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7887 ( .C ( clk ), .D ( new_AGEMA_signal_24661 ), .Q ( new_AGEMA_signal_24662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7901 ( .C ( clk ), .D ( new_AGEMA_signal_24675 ), .Q ( new_AGEMA_signal_24676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7915 ( .C ( clk ), .D ( new_AGEMA_signal_24689 ), .Q ( new_AGEMA_signal_24690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7923 ( .C ( clk ), .D ( new_AGEMA_signal_24697 ), .Q ( new_AGEMA_signal_24698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7931 ( .C ( clk ), .D ( new_AGEMA_signal_24705 ), .Q ( new_AGEMA_signal_24706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7939 ( .C ( clk ), .D ( new_AGEMA_signal_24713 ), .Q ( new_AGEMA_signal_24714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7947 ( .C ( clk ), .D ( new_AGEMA_signal_24721 ), .Q ( new_AGEMA_signal_24722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7955 ( .C ( clk ), .D ( new_AGEMA_signal_24729 ), .Q ( new_AGEMA_signal_24730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7963 ( .C ( clk ), .D ( new_AGEMA_signal_24737 ), .Q ( new_AGEMA_signal_24738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7971 ( .C ( clk ), .D ( new_AGEMA_signal_24745 ), .Q ( new_AGEMA_signal_24746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7979 ( .C ( clk ), .D ( new_AGEMA_signal_24753 ), .Q ( new_AGEMA_signal_24754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7987 ( .C ( clk ), .D ( new_AGEMA_signal_24761 ), .Q ( new_AGEMA_signal_24762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7995 ( .C ( clk ), .D ( new_AGEMA_signal_24769 ), .Q ( new_AGEMA_signal_24770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7997 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_24772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8001 ( .C ( clk ), .D ( new_AGEMA_signal_4366 ), .Q ( new_AGEMA_signal_24776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8005 ( .C ( clk ), .D ( new_AGEMA_signal_4367 ), .Q ( new_AGEMA_signal_24780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8009 ( .C ( clk ), .D ( new_AGEMA_signal_4368 ), .Q ( new_AGEMA_signal_24784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8013 ( .C ( clk ), .D ( new_AGEMA_signal_4369 ), .Q ( new_AGEMA_signal_24788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8039 ( .C ( clk ), .D ( new_AGEMA_signal_24813 ), .Q ( new_AGEMA_signal_24814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8055 ( .C ( clk ), .D ( new_AGEMA_signal_24829 ), .Q ( new_AGEMA_signal_24830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8071 ( .C ( clk ), .D ( new_AGEMA_signal_24845 ), .Q ( new_AGEMA_signal_24846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8087 ( .C ( clk ), .D ( new_AGEMA_signal_24861 ), .Q ( new_AGEMA_signal_24862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8103 ( .C ( clk ), .D ( new_AGEMA_signal_24877 ), .Q ( new_AGEMA_signal_24878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8107 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_24882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8111 ( .C ( clk ), .D ( new_AGEMA_signal_4402 ), .Q ( new_AGEMA_signal_24886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8115 ( .C ( clk ), .D ( new_AGEMA_signal_4403 ), .Q ( new_AGEMA_signal_24890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8119 ( .C ( clk ), .D ( new_AGEMA_signal_4404 ), .Q ( new_AGEMA_signal_24894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8123 ( .C ( clk ), .D ( new_AGEMA_signal_4405 ), .Q ( new_AGEMA_signal_24898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8149 ( .C ( clk ), .D ( new_AGEMA_signal_24923 ), .Q ( new_AGEMA_signal_24924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8165 ( .C ( clk ), .D ( new_AGEMA_signal_24939 ), .Q ( new_AGEMA_signal_24940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8181 ( .C ( clk ), .D ( new_AGEMA_signal_24955 ), .Q ( new_AGEMA_signal_24956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8197 ( .C ( clk ), .D ( new_AGEMA_signal_24971 ), .Q ( new_AGEMA_signal_24972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8213 ( .C ( clk ), .D ( new_AGEMA_signal_24987 ), .Q ( new_AGEMA_signal_24988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8223 ( .C ( clk ), .D ( new_AGEMA_signal_24997 ), .Q ( new_AGEMA_signal_24998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8233 ( .C ( clk ), .D ( new_AGEMA_signal_25007 ), .Q ( new_AGEMA_signal_25008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8243 ( .C ( clk ), .D ( new_AGEMA_signal_25017 ), .Q ( new_AGEMA_signal_25018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8253 ( .C ( clk ), .D ( new_AGEMA_signal_25027 ), .Q ( new_AGEMA_signal_25028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8263 ( .C ( clk ), .D ( new_AGEMA_signal_25037 ), .Q ( new_AGEMA_signal_25038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8267 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_25042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8271 ( .C ( clk ), .D ( new_AGEMA_signal_4446 ), .Q ( new_AGEMA_signal_25046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8275 ( .C ( clk ), .D ( new_AGEMA_signal_4447 ), .Q ( new_AGEMA_signal_25050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8279 ( .C ( clk ), .D ( new_AGEMA_signal_4448 ), .Q ( new_AGEMA_signal_25054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8283 ( .C ( clk ), .D ( new_AGEMA_signal_4449 ), .Q ( new_AGEMA_signal_25058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8291 ( .C ( clk ), .D ( new_AGEMA_signal_25065 ), .Q ( new_AGEMA_signal_25066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8299 ( .C ( clk ), .D ( new_AGEMA_signal_25073 ), .Q ( new_AGEMA_signal_25074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8307 ( .C ( clk ), .D ( new_AGEMA_signal_25081 ), .Q ( new_AGEMA_signal_25082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8315 ( .C ( clk ), .D ( new_AGEMA_signal_25089 ), .Q ( new_AGEMA_signal_25090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8323 ( .C ( clk ), .D ( new_AGEMA_signal_25097 ), .Q ( new_AGEMA_signal_25098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8327 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_25102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8333 ( .C ( clk ), .D ( new_AGEMA_signal_4374 ), .Q ( new_AGEMA_signal_25108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8339 ( .C ( clk ), .D ( new_AGEMA_signal_4375 ), .Q ( new_AGEMA_signal_25114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8345 ( .C ( clk ), .D ( new_AGEMA_signal_4376 ), .Q ( new_AGEMA_signal_25120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8351 ( .C ( clk ), .D ( new_AGEMA_signal_4377 ), .Q ( new_AGEMA_signal_25126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8357 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_25132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8363 ( .C ( clk ), .D ( new_AGEMA_signal_4382 ), .Q ( new_AGEMA_signal_25138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8369 ( .C ( clk ), .D ( new_AGEMA_signal_4383 ), .Q ( new_AGEMA_signal_25144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8375 ( .C ( clk ), .D ( new_AGEMA_signal_4384 ), .Q ( new_AGEMA_signal_25150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8381 ( .C ( clk ), .D ( new_AGEMA_signal_4385 ), .Q ( new_AGEMA_signal_25156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8397 ( .C ( clk ), .D ( new_AGEMA_signal_25171 ), .Q ( new_AGEMA_signal_25172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8413 ( .C ( clk ), .D ( new_AGEMA_signal_25187 ), .Q ( new_AGEMA_signal_25188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8429 ( .C ( clk ), .D ( new_AGEMA_signal_25203 ), .Q ( new_AGEMA_signal_25204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8445 ( .C ( clk ), .D ( new_AGEMA_signal_25219 ), .Q ( new_AGEMA_signal_25220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8461 ( .C ( clk ), .D ( new_AGEMA_signal_25235 ), .Q ( new_AGEMA_signal_25236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8471 ( .C ( clk ), .D ( new_AGEMA_signal_25245 ), .Q ( new_AGEMA_signal_25246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8481 ( .C ( clk ), .D ( new_AGEMA_signal_25255 ), .Q ( new_AGEMA_signal_25256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8491 ( .C ( clk ), .D ( new_AGEMA_signal_25265 ), .Q ( new_AGEMA_signal_25266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8501 ( .C ( clk ), .D ( new_AGEMA_signal_25275 ), .Q ( new_AGEMA_signal_25276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8511 ( .C ( clk ), .D ( new_AGEMA_signal_25285 ), .Q ( new_AGEMA_signal_25286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8529 ( .C ( clk ), .D ( new_AGEMA_signal_25303 ), .Q ( new_AGEMA_signal_25304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8547 ( .C ( clk ), .D ( new_AGEMA_signal_25321 ), .Q ( new_AGEMA_signal_25322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8565 ( .C ( clk ), .D ( new_AGEMA_signal_25339 ), .Q ( new_AGEMA_signal_25340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8583 ( .C ( clk ), .D ( new_AGEMA_signal_25357 ), .Q ( new_AGEMA_signal_25358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8601 ( .C ( clk ), .D ( new_AGEMA_signal_25375 ), .Q ( new_AGEMA_signal_25376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8629 ( .C ( clk ), .D ( new_AGEMA_signal_25403 ), .Q ( new_AGEMA_signal_25404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8637 ( .C ( clk ), .D ( new_AGEMA_signal_25411 ), .Q ( new_AGEMA_signal_25412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8645 ( .C ( clk ), .D ( new_AGEMA_signal_25419 ), .Q ( new_AGEMA_signal_25420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8653 ( .C ( clk ), .D ( new_AGEMA_signal_25427 ), .Q ( new_AGEMA_signal_25428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8661 ( .C ( clk ), .D ( new_AGEMA_signal_25435 ), .Q ( new_AGEMA_signal_25436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8687 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_25462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8695 ( .C ( clk ), .D ( new_AGEMA_signal_4362 ), .Q ( new_AGEMA_signal_25470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8703 ( .C ( clk ), .D ( new_AGEMA_signal_4363 ), .Q ( new_AGEMA_signal_25478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8711 ( .C ( clk ), .D ( new_AGEMA_signal_4364 ), .Q ( new_AGEMA_signal_25486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8719 ( .C ( clk ), .D ( new_AGEMA_signal_4365 ), .Q ( new_AGEMA_signal_25494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8779 ( .C ( clk ), .D ( new_AGEMA_signal_25553 ), .Q ( new_AGEMA_signal_25554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8799 ( .C ( clk ), .D ( new_AGEMA_signal_25573 ), .Q ( new_AGEMA_signal_25574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8819 ( .C ( clk ), .D ( new_AGEMA_signal_25593 ), .Q ( new_AGEMA_signal_25594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8839 ( .C ( clk ), .D ( new_AGEMA_signal_25613 ), .Q ( new_AGEMA_signal_25614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8859 ( .C ( clk ), .D ( new_AGEMA_signal_25633 ), .Q ( new_AGEMA_signal_25634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8909 ( .C ( clk ), .D ( new_AGEMA_signal_25683 ), .Q ( new_AGEMA_signal_25684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8921 ( .C ( clk ), .D ( new_AGEMA_signal_25695 ), .Q ( new_AGEMA_signal_25696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8933 ( .C ( clk ), .D ( new_AGEMA_signal_25707 ), .Q ( new_AGEMA_signal_25708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8945 ( .C ( clk ), .D ( new_AGEMA_signal_25719 ), .Q ( new_AGEMA_signal_25720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8957 ( .C ( clk ), .D ( new_AGEMA_signal_25731 ), .Q ( new_AGEMA_signal_25732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8969 ( .C ( clk ), .D ( new_AGEMA_signal_25743 ), .Q ( new_AGEMA_signal_25744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8983 ( .C ( clk ), .D ( new_AGEMA_signal_25757 ), .Q ( new_AGEMA_signal_25758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8997 ( .C ( clk ), .D ( new_AGEMA_signal_25771 ), .Q ( new_AGEMA_signal_25772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9011 ( .C ( clk ), .D ( new_AGEMA_signal_25785 ), .Q ( new_AGEMA_signal_25786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9025 ( .C ( clk ), .D ( new_AGEMA_signal_25799 ), .Q ( new_AGEMA_signal_25800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9037 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_25812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9051 ( .C ( clk ), .D ( new_AGEMA_signal_4426 ), .Q ( new_AGEMA_signal_25826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9065 ( .C ( clk ), .D ( new_AGEMA_signal_4427 ), .Q ( new_AGEMA_signal_25840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9079 ( .C ( clk ), .D ( new_AGEMA_signal_4428 ), .Q ( new_AGEMA_signal_25854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9093 ( .C ( clk ), .D ( new_AGEMA_signal_4429 ), .Q ( new_AGEMA_signal_25868 ) ) ;

    /* cells in depth 20 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2117 ( .ina ({new_AGEMA_signal_23951, new_AGEMA_signal_23945, new_AGEMA_signal_23939, new_AGEMA_signal_23933, new_AGEMA_signal_23927}), .inb ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, new_AGEMA_signal_4371, new_AGEMA_signal_4370, n1989}), .clk ( clk ), .rnd ({Fresh[12269], Fresh[12268], Fresh[12267], Fresh[12266], Fresh[12265], Fresh[12264], Fresh[12263], Fresh[12262], Fresh[12261], Fresh[12260], Fresh[12259], Fresh[12258], Fresh[12257], Fresh[12256], Fresh[12255]}), .outt ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, new_AGEMA_signal_4458, n2000}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2181 ( .ina ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, new_AGEMA_signal_4266, n2038}), .inb ({new_AGEMA_signal_23971, new_AGEMA_signal_23967, new_AGEMA_signal_23963, new_AGEMA_signal_23959, new_AGEMA_signal_23955}), .clk ( clk ), .rnd ({Fresh[12284], Fresh[12283], Fresh[12282], Fresh[12281], Fresh[12280], Fresh[12279], Fresh[12278], Fresh[12277], Fresh[12276], Fresh[12275], Fresh[12274], Fresh[12273], Fresh[12272], Fresh[12271], Fresh[12270]}), .outt ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, new_AGEMA_signal_4379, new_AGEMA_signal_4378, n2113}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2231 ( .ina ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, new_AGEMA_signal_4386, n2079}), .inb ({new_AGEMA_signal_24001, new_AGEMA_signal_23995, new_AGEMA_signal_23989, new_AGEMA_signal_23983, new_AGEMA_signal_23977}), .clk ( clk ), .rnd ({Fresh[12299], Fresh[12298], Fresh[12297], Fresh[12296], Fresh[12295], Fresh[12294], Fresh[12293], Fresh[12292], Fresh[12291], Fresh[12290], Fresh[12289], Fresh[12288], Fresh[12287], Fresh[12286], Fresh[12285]}), .outt ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, n2109}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2264 ( .ina ({new_AGEMA_signal_24051, new_AGEMA_signal_24041, new_AGEMA_signal_24031, new_AGEMA_signal_24021, new_AGEMA_signal_24011}), .inb ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, new_AGEMA_signal_4391, new_AGEMA_signal_4390, n2104}), .clk ( clk ), .rnd ({Fresh[12314], Fresh[12313], Fresh[12312], Fresh[12311], Fresh[12310], Fresh[12309], Fresh[12308], Fresh[12307], Fresh[12306], Fresh[12305], Fresh[12304], Fresh[12303], Fresh[12302], Fresh[12301], Fresh[12300]}), .outt ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, new_AGEMA_signal_4467, new_AGEMA_signal_4466, n2107}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2290 ( .ina ({new_AGEMA_signal_24081, new_AGEMA_signal_24075, new_AGEMA_signal_24069, new_AGEMA_signal_24063, new_AGEMA_signal_24057}), .inb ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, new_AGEMA_signal_4395, new_AGEMA_signal_4394, n2127}), .clk ( clk ), .rnd ({Fresh[12329], Fresh[12328], Fresh[12327], Fresh[12326], Fresh[12325], Fresh[12324], Fresh[12323], Fresh[12322], Fresh[12321], Fresh[12320], Fresh[12319], Fresh[12318], Fresh[12317], Fresh[12316], Fresh[12315]}), .outt ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, new_AGEMA_signal_4470, n2212}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2316 ( .ina ({new_AGEMA_signal_24111, new_AGEMA_signal_24105, new_AGEMA_signal_24099, new_AGEMA_signal_24093, new_AGEMA_signal_24087}), .inb ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, new_AGEMA_signal_4398, n2147}), .clk ( clk ), .rnd ({Fresh[12344], Fresh[12343], Fresh[12342], Fresh[12341], Fresh[12340], Fresh[12339], Fresh[12338], Fresh[12337], Fresh[12336], Fresh[12335], Fresh[12334], Fresh[12333], Fresh[12332], Fresh[12331], Fresh[12330]}), .outt ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, n2149}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2366 ( .ina ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, new_AGEMA_signal_4407, new_AGEMA_signal_4406, n2199}), .inb ({new_AGEMA_signal_24131, new_AGEMA_signal_24127, new_AGEMA_signal_24123, new_AGEMA_signal_24119, new_AGEMA_signal_24115}), .clk ( clk ), .rnd ({Fresh[12359], Fresh[12358], Fresh[12357], Fresh[12356], Fresh[12355], Fresh[12354], Fresh[12353], Fresh[12352], Fresh[12351], Fresh[12350], Fresh[12349], Fresh[12348], Fresh[12347], Fresh[12346], Fresh[12345]}), .outt ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, new_AGEMA_signal_4479, new_AGEMA_signal_4478, n2206}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2421 ( .ina ({new_AGEMA_signal_24151, new_AGEMA_signal_24147, new_AGEMA_signal_24143, new_AGEMA_signal_24139, new_AGEMA_signal_24135}), .inb ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, new_AGEMA_signal_4410, n2257}), .clk ( clk ), .rnd ({Fresh[12374], Fresh[12373], Fresh[12372], Fresh[12371], Fresh[12370], Fresh[12369], Fresh[12368], Fresh[12367], Fresh[12366], Fresh[12365], Fresh[12364], Fresh[12363], Fresh[12362], Fresh[12361], Fresh[12360]}), .outt ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, new_AGEMA_signal_4482, n2310}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2447 ( .ina ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, new_AGEMA_signal_4415, new_AGEMA_signal_4414, n2281}), .inb ({new_AGEMA_signal_24191, new_AGEMA_signal_24183, new_AGEMA_signal_24175, new_AGEMA_signal_24167, new_AGEMA_signal_24159}), .clk ( clk ), .rnd ({Fresh[12389], Fresh[12388], Fresh[12387], Fresh[12386], Fresh[12385], Fresh[12384], Fresh[12383], Fresh[12382], Fresh[12381], Fresh[12380], Fresh[12379], Fresh[12378], Fresh[12377], Fresh[12376], Fresh[12375]}), .outt ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, n2308}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2476 ( .ina ({new_AGEMA_signal_24221, new_AGEMA_signal_24215, new_AGEMA_signal_24209, new_AGEMA_signal_24203, new_AGEMA_signal_24197}), .inb ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, new_AGEMA_signal_4419, new_AGEMA_signal_4418, n2305}), .clk ( clk ), .rnd ({Fresh[12404], Fresh[12403], Fresh[12402], Fresh[12401], Fresh[12400], Fresh[12399], Fresh[12398], Fresh[12397], Fresh[12396], Fresh[12395], Fresh[12394], Fresh[12393], Fresh[12392], Fresh[12391], Fresh[12390]}), .outt ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, new_AGEMA_signal_4491, new_AGEMA_signal_4490, n2307}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2533 ( .ina ({new_AGEMA_signal_24261, new_AGEMA_signal_24253, new_AGEMA_signal_24245, new_AGEMA_signal_24237, new_AGEMA_signal_24229}), .inb ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, new_AGEMA_signal_4423, new_AGEMA_signal_4422, n2368}), .clk ( clk ), .rnd ({Fresh[12419], Fresh[12418], Fresh[12417], Fresh[12416], Fresh[12415], Fresh[12414], Fresh[12413], Fresh[12412], Fresh[12411], Fresh[12410], Fresh[12409], Fresh[12408], Fresh[12407], Fresh[12406], Fresh[12405]}), .outt ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, new_AGEMA_signal_4494, n2370}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2611 ( .ina ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, new_AGEMA_signal_4431, new_AGEMA_signal_4430, n2457}), .inb ({new_AGEMA_signal_24301, new_AGEMA_signal_24293, new_AGEMA_signal_24285, new_AGEMA_signal_24277, new_AGEMA_signal_24269}), .clk ( clk ), .rnd ({Fresh[12434], Fresh[12433], Fresh[12432], Fresh[12431], Fresh[12430], Fresh[12429], Fresh[12428], Fresh[12427], Fresh[12426], Fresh[12425], Fresh[12424], Fresh[12423], Fresh[12422], Fresh[12421], Fresh[12420]}), .outt ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, n2530}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2660 ( .ina ({new_AGEMA_signal_24311, new_AGEMA_signal_24309, new_AGEMA_signal_24307, new_AGEMA_signal_24305, new_AGEMA_signal_24303}), .inb ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, new_AGEMA_signal_4435, new_AGEMA_signal_4434, n2513}), .clk ( clk ), .rnd ({Fresh[12449], Fresh[12448], Fresh[12447], Fresh[12446], Fresh[12445], Fresh[12444], Fresh[12443], Fresh[12442], Fresh[12441], Fresh[12440], Fresh[12439], Fresh[12438], Fresh[12437], Fresh[12436], Fresh[12435]}), .outt ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, new_AGEMA_signal_4503, new_AGEMA_signal_4502, n2515}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2718 ( .ina ({new_AGEMA_signal_24331, new_AGEMA_signal_24327, new_AGEMA_signal_24323, new_AGEMA_signal_24319, new_AGEMA_signal_24315}), .inb ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, new_AGEMA_signal_4439, new_AGEMA_signal_4438, n2592}), .clk ( clk ), .rnd ({Fresh[12464], Fresh[12463], Fresh[12462], Fresh[12461], Fresh[12460], Fresh[12459], Fresh[12458], Fresh[12457], Fresh[12456], Fresh[12455], Fresh[12454], Fresh[12453], Fresh[12452], Fresh[12451], Fresh[12450]}), .outt ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, new_AGEMA_signal_4506, n2639}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2749 ( .ina ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, new_AGEMA_signal_4347, new_AGEMA_signal_4346, n2637}), .inb ({new_AGEMA_signal_24351, new_AGEMA_signal_24347, new_AGEMA_signal_24343, new_AGEMA_signal_24339, new_AGEMA_signal_24335}), .clk ( clk ), .rnd ({Fresh[12479], Fresh[12478], Fresh[12477], Fresh[12476], Fresh[12475], Fresh[12474], Fresh[12473], Fresh[12472], Fresh[12471], Fresh[12470], Fresh[12469], Fresh[12468], Fresh[12467], Fresh[12466], Fresh[12465]}), .outt ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, new_AGEMA_signal_4443, new_AGEMA_signal_4442, n2638}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2788 ( .ina ({new_AGEMA_signal_24391, new_AGEMA_signal_24383, new_AGEMA_signal_24375, new_AGEMA_signal_24367, new_AGEMA_signal_24359}), .inb ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, n2705}), .clk ( clk ), .rnd ({Fresh[12494], Fresh[12493], Fresh[12492], Fresh[12491], Fresh[12490], Fresh[12489], Fresh[12488], Fresh[12487], Fresh[12486], Fresh[12485], Fresh[12484], Fresh[12483], Fresh[12482], Fresh[12481], Fresh[12480]}), .outt ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, n2832}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2842 ( .ina ({new_AGEMA_signal_24411, new_AGEMA_signal_24407, new_AGEMA_signal_24403, new_AGEMA_signal_24399, new_AGEMA_signal_24395}), .inb ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, new_AGEMA_signal_4359, new_AGEMA_signal_4358, n2805}), .clk ( clk ), .rnd ({Fresh[12509], Fresh[12508], Fresh[12507], Fresh[12506], Fresh[12505], Fresh[12504], Fresh[12503], Fresh[12502], Fresh[12501], Fresh[12500], Fresh[12499], Fresh[12498], Fresh[12497], Fresh[12496], Fresh[12495]}), .outt ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, new_AGEMA_signal_4455, new_AGEMA_signal_4454, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C ( clk ), .D ( new_AGEMA_signal_24418 ), .Q ( new_AGEMA_signal_24419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C ( clk ), .D ( new_AGEMA_signal_24426 ), .Q ( new_AGEMA_signal_24427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C ( clk ), .D ( new_AGEMA_signal_24434 ), .Q ( new_AGEMA_signal_24435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7668 ( .C ( clk ), .D ( new_AGEMA_signal_24442 ), .Q ( new_AGEMA_signal_24443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7676 ( .C ( clk ), .D ( new_AGEMA_signal_24450 ), .Q ( new_AGEMA_signal_24451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7688 ( .C ( clk ), .D ( new_AGEMA_signal_24462 ), .Q ( new_AGEMA_signal_24463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7700 ( .C ( clk ), .D ( new_AGEMA_signal_24474 ), .Q ( new_AGEMA_signal_24475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7712 ( .C ( clk ), .D ( new_AGEMA_signal_24486 ), .Q ( new_AGEMA_signal_24487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7724 ( .C ( clk ), .D ( new_AGEMA_signal_24498 ), .Q ( new_AGEMA_signal_24499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7736 ( .C ( clk ), .D ( new_AGEMA_signal_24510 ), .Q ( new_AGEMA_signal_24511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7750 ( .C ( clk ), .D ( new_AGEMA_signal_24524 ), .Q ( new_AGEMA_signal_24525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7764 ( .C ( clk ), .D ( new_AGEMA_signal_24538 ), .Q ( new_AGEMA_signal_24539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7778 ( .C ( clk ), .D ( new_AGEMA_signal_24552 ), .Q ( new_AGEMA_signal_24553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7792 ( .C ( clk ), .D ( new_AGEMA_signal_24566 ), .Q ( new_AGEMA_signal_24567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7806 ( .C ( clk ), .D ( new_AGEMA_signal_24580 ), .Q ( new_AGEMA_signal_24581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7814 ( .C ( clk ), .D ( new_AGEMA_signal_24588 ), .Q ( new_AGEMA_signal_24589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7822 ( .C ( clk ), .D ( new_AGEMA_signal_24596 ), .Q ( new_AGEMA_signal_24597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7830 ( .C ( clk ), .D ( new_AGEMA_signal_24604 ), .Q ( new_AGEMA_signal_24605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7838 ( .C ( clk ), .D ( new_AGEMA_signal_24612 ), .Q ( new_AGEMA_signal_24613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7846 ( .C ( clk ), .D ( new_AGEMA_signal_24620 ), .Q ( new_AGEMA_signal_24621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7860 ( .C ( clk ), .D ( new_AGEMA_signal_24634 ), .Q ( new_AGEMA_signal_24635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7874 ( .C ( clk ), .D ( new_AGEMA_signal_24648 ), .Q ( new_AGEMA_signal_24649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7888 ( .C ( clk ), .D ( new_AGEMA_signal_24662 ), .Q ( new_AGEMA_signal_24663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7902 ( .C ( clk ), .D ( new_AGEMA_signal_24676 ), .Q ( new_AGEMA_signal_24677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7916 ( .C ( clk ), .D ( new_AGEMA_signal_24690 ), .Q ( new_AGEMA_signal_24691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7924 ( .C ( clk ), .D ( new_AGEMA_signal_24698 ), .Q ( new_AGEMA_signal_24699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7932 ( .C ( clk ), .D ( new_AGEMA_signal_24706 ), .Q ( new_AGEMA_signal_24707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7940 ( .C ( clk ), .D ( new_AGEMA_signal_24714 ), .Q ( new_AGEMA_signal_24715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7948 ( .C ( clk ), .D ( new_AGEMA_signal_24722 ), .Q ( new_AGEMA_signal_24723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7956 ( .C ( clk ), .D ( new_AGEMA_signal_24730 ), .Q ( new_AGEMA_signal_24731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7964 ( .C ( clk ), .D ( new_AGEMA_signal_24738 ), .Q ( new_AGEMA_signal_24739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7972 ( .C ( clk ), .D ( new_AGEMA_signal_24746 ), .Q ( new_AGEMA_signal_24747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7980 ( .C ( clk ), .D ( new_AGEMA_signal_24754 ), .Q ( new_AGEMA_signal_24755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7988 ( .C ( clk ), .D ( new_AGEMA_signal_24762 ), .Q ( new_AGEMA_signal_24763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7996 ( .C ( clk ), .D ( new_AGEMA_signal_24770 ), .Q ( new_AGEMA_signal_24771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7998 ( .C ( clk ), .D ( new_AGEMA_signal_24772 ), .Q ( new_AGEMA_signal_24773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8002 ( .C ( clk ), .D ( new_AGEMA_signal_24776 ), .Q ( new_AGEMA_signal_24777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8006 ( .C ( clk ), .D ( new_AGEMA_signal_24780 ), .Q ( new_AGEMA_signal_24781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8010 ( .C ( clk ), .D ( new_AGEMA_signal_24784 ), .Q ( new_AGEMA_signal_24785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8014 ( .C ( clk ), .D ( new_AGEMA_signal_24788 ), .Q ( new_AGEMA_signal_24789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8040 ( .C ( clk ), .D ( new_AGEMA_signal_24814 ), .Q ( new_AGEMA_signal_24815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8056 ( .C ( clk ), .D ( new_AGEMA_signal_24830 ), .Q ( new_AGEMA_signal_24831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8072 ( .C ( clk ), .D ( new_AGEMA_signal_24846 ), .Q ( new_AGEMA_signal_24847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8088 ( .C ( clk ), .D ( new_AGEMA_signal_24862 ), .Q ( new_AGEMA_signal_24863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8104 ( .C ( clk ), .D ( new_AGEMA_signal_24878 ), .Q ( new_AGEMA_signal_24879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8108 ( .C ( clk ), .D ( new_AGEMA_signal_24882 ), .Q ( new_AGEMA_signal_24883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8112 ( .C ( clk ), .D ( new_AGEMA_signal_24886 ), .Q ( new_AGEMA_signal_24887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8116 ( .C ( clk ), .D ( new_AGEMA_signal_24890 ), .Q ( new_AGEMA_signal_24891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8120 ( .C ( clk ), .D ( new_AGEMA_signal_24894 ), .Q ( new_AGEMA_signal_24895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8124 ( .C ( clk ), .D ( new_AGEMA_signal_24898 ), .Q ( new_AGEMA_signal_24899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8150 ( .C ( clk ), .D ( new_AGEMA_signal_24924 ), .Q ( new_AGEMA_signal_24925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8166 ( .C ( clk ), .D ( new_AGEMA_signal_24940 ), .Q ( new_AGEMA_signal_24941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8182 ( .C ( clk ), .D ( new_AGEMA_signal_24956 ), .Q ( new_AGEMA_signal_24957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8198 ( .C ( clk ), .D ( new_AGEMA_signal_24972 ), .Q ( new_AGEMA_signal_24973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8214 ( .C ( clk ), .D ( new_AGEMA_signal_24988 ), .Q ( new_AGEMA_signal_24989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8224 ( .C ( clk ), .D ( new_AGEMA_signal_24998 ), .Q ( new_AGEMA_signal_24999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8234 ( .C ( clk ), .D ( new_AGEMA_signal_25008 ), .Q ( new_AGEMA_signal_25009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8244 ( .C ( clk ), .D ( new_AGEMA_signal_25018 ), .Q ( new_AGEMA_signal_25019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8254 ( .C ( clk ), .D ( new_AGEMA_signal_25028 ), .Q ( new_AGEMA_signal_25029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8264 ( .C ( clk ), .D ( new_AGEMA_signal_25038 ), .Q ( new_AGEMA_signal_25039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8268 ( .C ( clk ), .D ( new_AGEMA_signal_25042 ), .Q ( new_AGEMA_signal_25043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8272 ( .C ( clk ), .D ( new_AGEMA_signal_25046 ), .Q ( new_AGEMA_signal_25047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8276 ( .C ( clk ), .D ( new_AGEMA_signal_25050 ), .Q ( new_AGEMA_signal_25051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8280 ( .C ( clk ), .D ( new_AGEMA_signal_25054 ), .Q ( new_AGEMA_signal_25055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8284 ( .C ( clk ), .D ( new_AGEMA_signal_25058 ), .Q ( new_AGEMA_signal_25059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8292 ( .C ( clk ), .D ( new_AGEMA_signal_25066 ), .Q ( new_AGEMA_signal_25067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8300 ( .C ( clk ), .D ( new_AGEMA_signal_25074 ), .Q ( new_AGEMA_signal_25075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8308 ( .C ( clk ), .D ( new_AGEMA_signal_25082 ), .Q ( new_AGEMA_signal_25083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8316 ( .C ( clk ), .D ( new_AGEMA_signal_25090 ), .Q ( new_AGEMA_signal_25091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8324 ( .C ( clk ), .D ( new_AGEMA_signal_25098 ), .Q ( new_AGEMA_signal_25099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8328 ( .C ( clk ), .D ( new_AGEMA_signal_25102 ), .Q ( new_AGEMA_signal_25103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8334 ( .C ( clk ), .D ( new_AGEMA_signal_25108 ), .Q ( new_AGEMA_signal_25109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8340 ( .C ( clk ), .D ( new_AGEMA_signal_25114 ), .Q ( new_AGEMA_signal_25115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8346 ( .C ( clk ), .D ( new_AGEMA_signal_25120 ), .Q ( new_AGEMA_signal_25121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8352 ( .C ( clk ), .D ( new_AGEMA_signal_25126 ), .Q ( new_AGEMA_signal_25127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8358 ( .C ( clk ), .D ( new_AGEMA_signal_25132 ), .Q ( new_AGEMA_signal_25133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8364 ( .C ( clk ), .D ( new_AGEMA_signal_25138 ), .Q ( new_AGEMA_signal_25139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8370 ( .C ( clk ), .D ( new_AGEMA_signal_25144 ), .Q ( new_AGEMA_signal_25145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8376 ( .C ( clk ), .D ( new_AGEMA_signal_25150 ), .Q ( new_AGEMA_signal_25151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8382 ( .C ( clk ), .D ( new_AGEMA_signal_25156 ), .Q ( new_AGEMA_signal_25157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8398 ( .C ( clk ), .D ( new_AGEMA_signal_25172 ), .Q ( new_AGEMA_signal_25173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8414 ( .C ( clk ), .D ( new_AGEMA_signal_25188 ), .Q ( new_AGEMA_signal_25189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8430 ( .C ( clk ), .D ( new_AGEMA_signal_25204 ), .Q ( new_AGEMA_signal_25205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8446 ( .C ( clk ), .D ( new_AGEMA_signal_25220 ), .Q ( new_AGEMA_signal_25221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8462 ( .C ( clk ), .D ( new_AGEMA_signal_25236 ), .Q ( new_AGEMA_signal_25237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8472 ( .C ( clk ), .D ( new_AGEMA_signal_25246 ), .Q ( new_AGEMA_signal_25247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8482 ( .C ( clk ), .D ( new_AGEMA_signal_25256 ), .Q ( new_AGEMA_signal_25257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8492 ( .C ( clk ), .D ( new_AGEMA_signal_25266 ), .Q ( new_AGEMA_signal_25267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8502 ( .C ( clk ), .D ( new_AGEMA_signal_25276 ), .Q ( new_AGEMA_signal_25277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8512 ( .C ( clk ), .D ( new_AGEMA_signal_25286 ), .Q ( new_AGEMA_signal_25287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8530 ( .C ( clk ), .D ( new_AGEMA_signal_25304 ), .Q ( new_AGEMA_signal_25305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8548 ( .C ( clk ), .D ( new_AGEMA_signal_25322 ), .Q ( new_AGEMA_signal_25323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8566 ( .C ( clk ), .D ( new_AGEMA_signal_25340 ), .Q ( new_AGEMA_signal_25341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8584 ( .C ( clk ), .D ( new_AGEMA_signal_25358 ), .Q ( new_AGEMA_signal_25359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8602 ( .C ( clk ), .D ( new_AGEMA_signal_25376 ), .Q ( new_AGEMA_signal_25377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8630 ( .C ( clk ), .D ( new_AGEMA_signal_25404 ), .Q ( new_AGEMA_signal_25405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8638 ( .C ( clk ), .D ( new_AGEMA_signal_25412 ), .Q ( new_AGEMA_signal_25413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8646 ( .C ( clk ), .D ( new_AGEMA_signal_25420 ), .Q ( new_AGEMA_signal_25421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8654 ( .C ( clk ), .D ( new_AGEMA_signal_25428 ), .Q ( new_AGEMA_signal_25429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8662 ( .C ( clk ), .D ( new_AGEMA_signal_25436 ), .Q ( new_AGEMA_signal_25437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8688 ( .C ( clk ), .D ( new_AGEMA_signal_25462 ), .Q ( new_AGEMA_signal_25463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8696 ( .C ( clk ), .D ( new_AGEMA_signal_25470 ), .Q ( new_AGEMA_signal_25471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8704 ( .C ( clk ), .D ( new_AGEMA_signal_25478 ), .Q ( new_AGEMA_signal_25479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8712 ( .C ( clk ), .D ( new_AGEMA_signal_25486 ), .Q ( new_AGEMA_signal_25487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8720 ( .C ( clk ), .D ( new_AGEMA_signal_25494 ), .Q ( new_AGEMA_signal_25495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8780 ( .C ( clk ), .D ( new_AGEMA_signal_25554 ), .Q ( new_AGEMA_signal_25555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8800 ( .C ( clk ), .D ( new_AGEMA_signal_25574 ), .Q ( new_AGEMA_signal_25575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8820 ( .C ( clk ), .D ( new_AGEMA_signal_25594 ), .Q ( new_AGEMA_signal_25595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8840 ( .C ( clk ), .D ( new_AGEMA_signal_25614 ), .Q ( new_AGEMA_signal_25615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8860 ( .C ( clk ), .D ( new_AGEMA_signal_25634 ), .Q ( new_AGEMA_signal_25635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8910 ( .C ( clk ), .D ( new_AGEMA_signal_25684 ), .Q ( new_AGEMA_signal_25685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8922 ( .C ( clk ), .D ( new_AGEMA_signal_25696 ), .Q ( new_AGEMA_signal_25697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8934 ( .C ( clk ), .D ( new_AGEMA_signal_25708 ), .Q ( new_AGEMA_signal_25709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8946 ( .C ( clk ), .D ( new_AGEMA_signal_25720 ), .Q ( new_AGEMA_signal_25721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8958 ( .C ( clk ), .D ( new_AGEMA_signal_25732 ), .Q ( new_AGEMA_signal_25733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8970 ( .C ( clk ), .D ( new_AGEMA_signal_25744 ), .Q ( new_AGEMA_signal_25745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8984 ( .C ( clk ), .D ( new_AGEMA_signal_25758 ), .Q ( new_AGEMA_signal_25759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8998 ( .C ( clk ), .D ( new_AGEMA_signal_25772 ), .Q ( new_AGEMA_signal_25773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9012 ( .C ( clk ), .D ( new_AGEMA_signal_25786 ), .Q ( new_AGEMA_signal_25787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9026 ( .C ( clk ), .D ( new_AGEMA_signal_25800 ), .Q ( new_AGEMA_signal_25801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9038 ( .C ( clk ), .D ( new_AGEMA_signal_25812 ), .Q ( new_AGEMA_signal_25813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9052 ( .C ( clk ), .D ( new_AGEMA_signal_25826 ), .Q ( new_AGEMA_signal_25827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9066 ( .C ( clk ), .D ( new_AGEMA_signal_25840 ), .Q ( new_AGEMA_signal_25841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9080 ( .C ( clk ), .D ( new_AGEMA_signal_25854 ), .Q ( new_AGEMA_signal_25855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9094 ( .C ( clk ), .D ( new_AGEMA_signal_25868 ), .Q ( new_AGEMA_signal_25869 ) ) ;

    /* cells in depth 21 */
    buf_clk new_AGEMA_reg_buffer_7999 ( .C ( clk ), .D ( new_AGEMA_signal_24773 ), .Q ( new_AGEMA_signal_24774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8003 ( .C ( clk ), .D ( new_AGEMA_signal_24777 ), .Q ( new_AGEMA_signal_24778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8007 ( .C ( clk ), .D ( new_AGEMA_signal_24781 ), .Q ( new_AGEMA_signal_24782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8011 ( .C ( clk ), .D ( new_AGEMA_signal_24785 ), .Q ( new_AGEMA_signal_24786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8015 ( .C ( clk ), .D ( new_AGEMA_signal_24789 ), .Q ( new_AGEMA_signal_24790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8017 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_24792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8019 ( .C ( clk ), .D ( new_AGEMA_signal_4462 ), .Q ( new_AGEMA_signal_24794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8021 ( .C ( clk ), .D ( new_AGEMA_signal_4463 ), .Q ( new_AGEMA_signal_24796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8023 ( .C ( clk ), .D ( new_AGEMA_signal_4464 ), .Q ( new_AGEMA_signal_24798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8025 ( .C ( clk ), .D ( new_AGEMA_signal_4465 ), .Q ( new_AGEMA_signal_24800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8041 ( .C ( clk ), .D ( new_AGEMA_signal_24815 ), .Q ( new_AGEMA_signal_24816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8057 ( .C ( clk ), .D ( new_AGEMA_signal_24831 ), .Q ( new_AGEMA_signal_24832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8073 ( .C ( clk ), .D ( new_AGEMA_signal_24847 ), .Q ( new_AGEMA_signal_24848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8089 ( .C ( clk ), .D ( new_AGEMA_signal_24863 ), .Q ( new_AGEMA_signal_24864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8105 ( .C ( clk ), .D ( new_AGEMA_signal_24879 ), .Q ( new_AGEMA_signal_24880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8109 ( .C ( clk ), .D ( new_AGEMA_signal_24883 ), .Q ( new_AGEMA_signal_24884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8113 ( .C ( clk ), .D ( new_AGEMA_signal_24887 ), .Q ( new_AGEMA_signal_24888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8117 ( .C ( clk ), .D ( new_AGEMA_signal_24891 ), .Q ( new_AGEMA_signal_24892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8121 ( .C ( clk ), .D ( new_AGEMA_signal_24895 ), .Q ( new_AGEMA_signal_24896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8125 ( .C ( clk ), .D ( new_AGEMA_signal_24899 ), .Q ( new_AGEMA_signal_24900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8127 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_24902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8129 ( .C ( clk ), .D ( new_AGEMA_signal_4482 ), .Q ( new_AGEMA_signal_24904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8131 ( .C ( clk ), .D ( new_AGEMA_signal_4483 ), .Q ( new_AGEMA_signal_24906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8133 ( .C ( clk ), .D ( new_AGEMA_signal_4484 ), .Q ( new_AGEMA_signal_24908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8135 ( .C ( clk ), .D ( new_AGEMA_signal_4485 ), .Q ( new_AGEMA_signal_24910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8151 ( .C ( clk ), .D ( new_AGEMA_signal_24925 ), .Q ( new_AGEMA_signal_24926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8167 ( .C ( clk ), .D ( new_AGEMA_signal_24941 ), .Q ( new_AGEMA_signal_24942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8183 ( .C ( clk ), .D ( new_AGEMA_signal_24957 ), .Q ( new_AGEMA_signal_24958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8199 ( .C ( clk ), .D ( new_AGEMA_signal_24973 ), .Q ( new_AGEMA_signal_24974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8215 ( .C ( clk ), .D ( new_AGEMA_signal_24989 ), .Q ( new_AGEMA_signal_24990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8225 ( .C ( clk ), .D ( new_AGEMA_signal_24999 ), .Q ( new_AGEMA_signal_25000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8235 ( .C ( clk ), .D ( new_AGEMA_signal_25009 ), .Q ( new_AGEMA_signal_25010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8245 ( .C ( clk ), .D ( new_AGEMA_signal_25019 ), .Q ( new_AGEMA_signal_25020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8255 ( .C ( clk ), .D ( new_AGEMA_signal_25029 ), .Q ( new_AGEMA_signal_25030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8265 ( .C ( clk ), .D ( new_AGEMA_signal_25039 ), .Q ( new_AGEMA_signal_25040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8269 ( .C ( clk ), .D ( new_AGEMA_signal_25043 ), .Q ( new_AGEMA_signal_25044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8273 ( .C ( clk ), .D ( new_AGEMA_signal_25047 ), .Q ( new_AGEMA_signal_25048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8277 ( .C ( clk ), .D ( new_AGEMA_signal_25051 ), .Q ( new_AGEMA_signal_25052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8281 ( .C ( clk ), .D ( new_AGEMA_signal_25055 ), .Q ( new_AGEMA_signal_25056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8285 ( .C ( clk ), .D ( new_AGEMA_signal_25059 ), .Q ( new_AGEMA_signal_25060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8293 ( .C ( clk ), .D ( new_AGEMA_signal_25067 ), .Q ( new_AGEMA_signal_25068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8301 ( .C ( clk ), .D ( new_AGEMA_signal_25075 ), .Q ( new_AGEMA_signal_25076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8309 ( .C ( clk ), .D ( new_AGEMA_signal_25083 ), .Q ( new_AGEMA_signal_25084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8317 ( .C ( clk ), .D ( new_AGEMA_signal_25091 ), .Q ( new_AGEMA_signal_25092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8325 ( .C ( clk ), .D ( new_AGEMA_signal_25099 ), .Q ( new_AGEMA_signal_25100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8329 ( .C ( clk ), .D ( new_AGEMA_signal_25103 ), .Q ( new_AGEMA_signal_25104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8335 ( .C ( clk ), .D ( new_AGEMA_signal_25109 ), .Q ( new_AGEMA_signal_25110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8341 ( .C ( clk ), .D ( new_AGEMA_signal_25115 ), .Q ( new_AGEMA_signal_25116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8347 ( .C ( clk ), .D ( new_AGEMA_signal_25121 ), .Q ( new_AGEMA_signal_25122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8353 ( .C ( clk ), .D ( new_AGEMA_signal_25127 ), .Q ( new_AGEMA_signal_25128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8359 ( .C ( clk ), .D ( new_AGEMA_signal_25133 ), .Q ( new_AGEMA_signal_25134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8365 ( .C ( clk ), .D ( new_AGEMA_signal_25139 ), .Q ( new_AGEMA_signal_25140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8371 ( .C ( clk ), .D ( new_AGEMA_signal_25145 ), .Q ( new_AGEMA_signal_25146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8377 ( .C ( clk ), .D ( new_AGEMA_signal_25151 ), .Q ( new_AGEMA_signal_25152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8383 ( .C ( clk ), .D ( new_AGEMA_signal_25157 ), .Q ( new_AGEMA_signal_25158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8399 ( .C ( clk ), .D ( new_AGEMA_signal_25173 ), .Q ( new_AGEMA_signal_25174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8415 ( .C ( clk ), .D ( new_AGEMA_signal_25189 ), .Q ( new_AGEMA_signal_25190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8431 ( .C ( clk ), .D ( new_AGEMA_signal_25205 ), .Q ( new_AGEMA_signal_25206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8447 ( .C ( clk ), .D ( new_AGEMA_signal_25221 ), .Q ( new_AGEMA_signal_25222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8463 ( .C ( clk ), .D ( new_AGEMA_signal_25237 ), .Q ( new_AGEMA_signal_25238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8473 ( .C ( clk ), .D ( new_AGEMA_signal_25247 ), .Q ( new_AGEMA_signal_25248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8483 ( .C ( clk ), .D ( new_AGEMA_signal_25257 ), .Q ( new_AGEMA_signal_25258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8493 ( .C ( clk ), .D ( new_AGEMA_signal_25267 ), .Q ( new_AGEMA_signal_25268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8503 ( .C ( clk ), .D ( new_AGEMA_signal_25277 ), .Q ( new_AGEMA_signal_25278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8513 ( .C ( clk ), .D ( new_AGEMA_signal_25287 ), .Q ( new_AGEMA_signal_25288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8531 ( .C ( clk ), .D ( new_AGEMA_signal_25305 ), .Q ( new_AGEMA_signal_25306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8549 ( .C ( clk ), .D ( new_AGEMA_signal_25323 ), .Q ( new_AGEMA_signal_25324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8567 ( .C ( clk ), .D ( new_AGEMA_signal_25341 ), .Q ( new_AGEMA_signal_25342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8585 ( .C ( clk ), .D ( new_AGEMA_signal_25359 ), .Q ( new_AGEMA_signal_25360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8603 ( .C ( clk ), .D ( new_AGEMA_signal_25377 ), .Q ( new_AGEMA_signal_25378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8607 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_25382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8611 ( .C ( clk ), .D ( new_AGEMA_signal_4498 ), .Q ( new_AGEMA_signal_25386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8615 ( .C ( clk ), .D ( new_AGEMA_signal_4499 ), .Q ( new_AGEMA_signal_25390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8619 ( .C ( clk ), .D ( new_AGEMA_signal_4500 ), .Q ( new_AGEMA_signal_25394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8623 ( .C ( clk ), .D ( new_AGEMA_signal_4501 ), .Q ( new_AGEMA_signal_25398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8631 ( .C ( clk ), .D ( new_AGEMA_signal_25405 ), .Q ( new_AGEMA_signal_25406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8639 ( .C ( clk ), .D ( new_AGEMA_signal_25413 ), .Q ( new_AGEMA_signal_25414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8647 ( .C ( clk ), .D ( new_AGEMA_signal_25421 ), .Q ( new_AGEMA_signal_25422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8655 ( .C ( clk ), .D ( new_AGEMA_signal_25429 ), .Q ( new_AGEMA_signal_25430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8663 ( .C ( clk ), .D ( new_AGEMA_signal_25437 ), .Q ( new_AGEMA_signal_25438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8667 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_25442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8671 ( .C ( clk ), .D ( new_AGEMA_signal_4510 ), .Q ( new_AGEMA_signal_25446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8675 ( .C ( clk ), .D ( new_AGEMA_signal_4511 ), .Q ( new_AGEMA_signal_25450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8679 ( .C ( clk ), .D ( new_AGEMA_signal_4512 ), .Q ( new_AGEMA_signal_25454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8683 ( .C ( clk ), .D ( new_AGEMA_signal_4513 ), .Q ( new_AGEMA_signal_25458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8689 ( .C ( clk ), .D ( new_AGEMA_signal_25463 ), .Q ( new_AGEMA_signal_25464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8697 ( .C ( clk ), .D ( new_AGEMA_signal_25471 ), .Q ( new_AGEMA_signal_25472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8705 ( .C ( clk ), .D ( new_AGEMA_signal_25479 ), .Q ( new_AGEMA_signal_25480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8713 ( .C ( clk ), .D ( new_AGEMA_signal_25487 ), .Q ( new_AGEMA_signal_25488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8721 ( .C ( clk ), .D ( new_AGEMA_signal_25495 ), .Q ( new_AGEMA_signal_25496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8727 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_25502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8733 ( .C ( clk ), .D ( new_AGEMA_signal_4378 ), .Q ( new_AGEMA_signal_25508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8739 ( .C ( clk ), .D ( new_AGEMA_signal_4379 ), .Q ( new_AGEMA_signal_25514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8745 ( .C ( clk ), .D ( new_AGEMA_signal_4380 ), .Q ( new_AGEMA_signal_25520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8751 ( .C ( clk ), .D ( new_AGEMA_signal_4381 ), .Q ( new_AGEMA_signal_25526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8781 ( .C ( clk ), .D ( new_AGEMA_signal_25555 ), .Q ( new_AGEMA_signal_25556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8801 ( .C ( clk ), .D ( new_AGEMA_signal_25575 ), .Q ( new_AGEMA_signal_25576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8821 ( .C ( clk ), .D ( new_AGEMA_signal_25595 ), .Q ( new_AGEMA_signal_25596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8841 ( .C ( clk ), .D ( new_AGEMA_signal_25615 ), .Q ( new_AGEMA_signal_25616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8861 ( .C ( clk ), .D ( new_AGEMA_signal_25635 ), .Q ( new_AGEMA_signal_25636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8867 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_25642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8875 ( .C ( clk ), .D ( new_AGEMA_signal_4470 ), .Q ( new_AGEMA_signal_25650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8883 ( .C ( clk ), .D ( new_AGEMA_signal_4471 ), .Q ( new_AGEMA_signal_25658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8891 ( .C ( clk ), .D ( new_AGEMA_signal_4472 ), .Q ( new_AGEMA_signal_25666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8899 ( .C ( clk ), .D ( new_AGEMA_signal_4473 ), .Q ( new_AGEMA_signal_25674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8911 ( .C ( clk ), .D ( new_AGEMA_signal_25685 ), .Q ( new_AGEMA_signal_25686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8923 ( .C ( clk ), .D ( new_AGEMA_signal_25697 ), .Q ( new_AGEMA_signal_25698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8935 ( .C ( clk ), .D ( new_AGEMA_signal_25709 ), .Q ( new_AGEMA_signal_25710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8947 ( .C ( clk ), .D ( new_AGEMA_signal_25721 ), .Q ( new_AGEMA_signal_25722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8959 ( .C ( clk ), .D ( new_AGEMA_signal_25733 ), .Q ( new_AGEMA_signal_25734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8971 ( .C ( clk ), .D ( new_AGEMA_signal_25745 ), .Q ( new_AGEMA_signal_25746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8985 ( .C ( clk ), .D ( new_AGEMA_signal_25759 ), .Q ( new_AGEMA_signal_25760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8999 ( .C ( clk ), .D ( new_AGEMA_signal_25773 ), .Q ( new_AGEMA_signal_25774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9013 ( .C ( clk ), .D ( new_AGEMA_signal_25787 ), .Q ( new_AGEMA_signal_25788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9027 ( .C ( clk ), .D ( new_AGEMA_signal_25801 ), .Q ( new_AGEMA_signal_25802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9039 ( .C ( clk ), .D ( new_AGEMA_signal_25813 ), .Q ( new_AGEMA_signal_25814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9053 ( .C ( clk ), .D ( new_AGEMA_signal_25827 ), .Q ( new_AGEMA_signal_25828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9067 ( .C ( clk ), .D ( new_AGEMA_signal_25841 ), .Q ( new_AGEMA_signal_25842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9081 ( .C ( clk ), .D ( new_AGEMA_signal_25855 ), .Q ( new_AGEMA_signal_25856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9095 ( .C ( clk ), .D ( new_AGEMA_signal_25869 ), .Q ( new_AGEMA_signal_25870 ) ) ;

    /* cells in depth 22 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2129 ( .ina ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, new_AGEMA_signal_4458, n2000}), .inb ({new_AGEMA_signal_24451, new_AGEMA_signal_24443, new_AGEMA_signal_24435, new_AGEMA_signal_24427, new_AGEMA_signal_24419}), .clk ( clk ), .rnd ({Fresh[12524], Fresh[12523], Fresh[12522], Fresh[12521], Fresh[12520], Fresh[12519], Fresh[12518], Fresh[12517], Fresh[12516], Fresh[12515], Fresh[12514], Fresh[12513], Fresh[12512], Fresh[12511], Fresh[12510]}), .outt ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, new_AGEMA_signal_4518, n2001}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2267 ( .ina ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, new_AGEMA_signal_4467, new_AGEMA_signal_4466, n2107}), .inb ({new_AGEMA_signal_24511, new_AGEMA_signal_24499, new_AGEMA_signal_24487, new_AGEMA_signal_24475, new_AGEMA_signal_24463}), .clk ( clk ), .rnd ({Fresh[12539], Fresh[12538], Fresh[12537], Fresh[12536], Fresh[12535], Fresh[12534], Fresh[12533], Fresh[12532], Fresh[12531], Fresh[12530], Fresh[12529], Fresh[12528], Fresh[12527], Fresh[12526], Fresh[12525]}), .outt ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, n2108}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2317 ( .ina ({new_AGEMA_signal_24581, new_AGEMA_signal_24567, new_AGEMA_signal_24553, new_AGEMA_signal_24539, new_AGEMA_signal_24525}), .inb ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, n2149}), .clk ( clk ), .rnd ({Fresh[12554], Fresh[12553], Fresh[12552], Fresh[12551], Fresh[12550], Fresh[12549], Fresh[12548], Fresh[12547], Fresh[12546], Fresh[12545], Fresh[12544], Fresh[12543], Fresh[12542], Fresh[12541], Fresh[12540]}), .outt ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, n2153}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2374 ( .ina ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, new_AGEMA_signal_4479, new_AGEMA_signal_4478, n2206}), .inb ({new_AGEMA_signal_24621, new_AGEMA_signal_24613, new_AGEMA_signal_24605, new_AGEMA_signal_24597, new_AGEMA_signal_24589}), .clk ( clk ), .rnd ({Fresh[12569], Fresh[12568], Fresh[12567], Fresh[12566], Fresh[12565], Fresh[12564], Fresh[12563], Fresh[12562], Fresh[12561], Fresh[12560], Fresh[12559], Fresh[12558], Fresh[12557], Fresh[12556], Fresh[12555]}), .outt ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, new_AGEMA_signal_4530, n2207}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2477 ( .ina ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, n2308}), .inb ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, new_AGEMA_signal_4491, new_AGEMA_signal_4490, n2307}), .clk ( clk ), .rnd ({Fresh[12584], Fresh[12583], Fresh[12582], Fresh[12581], Fresh[12580], Fresh[12579], Fresh[12578], Fresh[12577], Fresh[12576], Fresh[12575], Fresh[12574], Fresh[12573], Fresh[12572], Fresh[12571], Fresh[12570]}), .outt ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, n2309}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2535 ( .ina ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, new_AGEMA_signal_4494, n2370}), .inb ({new_AGEMA_signal_24691, new_AGEMA_signal_24677, new_AGEMA_signal_24663, new_AGEMA_signal_24649, new_AGEMA_signal_24635}), .clk ( clk ), .rnd ({Fresh[12599], Fresh[12598], Fresh[12597], Fresh[12596], Fresh[12595], Fresh[12594], Fresh[12593], Fresh[12592], Fresh[12591], Fresh[12590], Fresh[12589], Fresh[12588], Fresh[12587], Fresh[12586], Fresh[12585]}), .outt ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, new_AGEMA_signal_4539, new_AGEMA_signal_4538, n2373}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2661 ( .ina ({new_AGEMA_signal_24731, new_AGEMA_signal_24723, new_AGEMA_signal_24715, new_AGEMA_signal_24707, new_AGEMA_signal_24699}), .inb ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, new_AGEMA_signal_4503, new_AGEMA_signal_4502, n2515}), .clk ( clk ), .rnd ({Fresh[12614], Fresh[12613], Fresh[12612], Fresh[12611], Fresh[12610], Fresh[12609], Fresh[12608], Fresh[12607], Fresh[12606], Fresh[12605], Fresh[12604], Fresh[12603], Fresh[12602], Fresh[12601], Fresh[12600]}), .outt ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, new_AGEMA_signal_4542, n2528}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2750 ( .ina ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, new_AGEMA_signal_4506, n2639}), .inb ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, new_AGEMA_signal_4443, new_AGEMA_signal_4442, n2638}), .clk ( clk ), .rnd ({Fresh[12629], Fresh[12628], Fresh[12627], Fresh[12626], Fresh[12625], Fresh[12624], Fresh[12623], Fresh[12622], Fresh[12621], Fresh[12620], Fresh[12619], Fresh[12618], Fresh[12617], Fresh[12616], Fresh[12615]}), .outt ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, n2669}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2843 ( .ina ({new_AGEMA_signal_24771, new_AGEMA_signal_24763, new_AGEMA_signal_24755, new_AGEMA_signal_24747, new_AGEMA_signal_24739}), .inb ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, new_AGEMA_signal_4455, new_AGEMA_signal_4454, n2807}), .clk ( clk ), .rnd ({Fresh[12644], Fresh[12643], Fresh[12642], Fresh[12641], Fresh[12640], Fresh[12639], Fresh[12638], Fresh[12637], Fresh[12636], Fresh[12635], Fresh[12634], Fresh[12633], Fresh[12632], Fresh[12631], Fresh[12630]}), .outt ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_8000 ( .C ( clk ), .D ( new_AGEMA_signal_24774 ), .Q ( new_AGEMA_signal_24775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8004 ( .C ( clk ), .D ( new_AGEMA_signal_24778 ), .Q ( new_AGEMA_signal_24779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8008 ( .C ( clk ), .D ( new_AGEMA_signal_24782 ), .Q ( new_AGEMA_signal_24783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8012 ( .C ( clk ), .D ( new_AGEMA_signal_24786 ), .Q ( new_AGEMA_signal_24787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8016 ( .C ( clk ), .D ( new_AGEMA_signal_24790 ), .Q ( new_AGEMA_signal_24791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8018 ( .C ( clk ), .D ( new_AGEMA_signal_24792 ), .Q ( new_AGEMA_signal_24793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8020 ( .C ( clk ), .D ( new_AGEMA_signal_24794 ), .Q ( new_AGEMA_signal_24795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8022 ( .C ( clk ), .D ( new_AGEMA_signal_24796 ), .Q ( new_AGEMA_signal_24797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8024 ( .C ( clk ), .D ( new_AGEMA_signal_24798 ), .Q ( new_AGEMA_signal_24799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8026 ( .C ( clk ), .D ( new_AGEMA_signal_24800 ), .Q ( new_AGEMA_signal_24801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8042 ( .C ( clk ), .D ( new_AGEMA_signal_24816 ), .Q ( new_AGEMA_signal_24817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8058 ( .C ( clk ), .D ( new_AGEMA_signal_24832 ), .Q ( new_AGEMA_signal_24833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8074 ( .C ( clk ), .D ( new_AGEMA_signal_24848 ), .Q ( new_AGEMA_signal_24849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8090 ( .C ( clk ), .D ( new_AGEMA_signal_24864 ), .Q ( new_AGEMA_signal_24865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8106 ( .C ( clk ), .D ( new_AGEMA_signal_24880 ), .Q ( new_AGEMA_signal_24881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8110 ( .C ( clk ), .D ( new_AGEMA_signal_24884 ), .Q ( new_AGEMA_signal_24885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8114 ( .C ( clk ), .D ( new_AGEMA_signal_24888 ), .Q ( new_AGEMA_signal_24889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8118 ( .C ( clk ), .D ( new_AGEMA_signal_24892 ), .Q ( new_AGEMA_signal_24893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8122 ( .C ( clk ), .D ( new_AGEMA_signal_24896 ), .Q ( new_AGEMA_signal_24897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8126 ( .C ( clk ), .D ( new_AGEMA_signal_24900 ), .Q ( new_AGEMA_signal_24901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8128 ( .C ( clk ), .D ( new_AGEMA_signal_24902 ), .Q ( new_AGEMA_signal_24903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8130 ( .C ( clk ), .D ( new_AGEMA_signal_24904 ), .Q ( new_AGEMA_signal_24905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8132 ( .C ( clk ), .D ( new_AGEMA_signal_24906 ), .Q ( new_AGEMA_signal_24907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8134 ( .C ( clk ), .D ( new_AGEMA_signal_24908 ), .Q ( new_AGEMA_signal_24909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8136 ( .C ( clk ), .D ( new_AGEMA_signal_24910 ), .Q ( new_AGEMA_signal_24911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8152 ( .C ( clk ), .D ( new_AGEMA_signal_24926 ), .Q ( new_AGEMA_signal_24927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8168 ( .C ( clk ), .D ( new_AGEMA_signal_24942 ), .Q ( new_AGEMA_signal_24943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8184 ( .C ( clk ), .D ( new_AGEMA_signal_24958 ), .Q ( new_AGEMA_signal_24959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8200 ( .C ( clk ), .D ( new_AGEMA_signal_24974 ), .Q ( new_AGEMA_signal_24975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8216 ( .C ( clk ), .D ( new_AGEMA_signal_24990 ), .Q ( new_AGEMA_signal_24991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8226 ( .C ( clk ), .D ( new_AGEMA_signal_25000 ), .Q ( new_AGEMA_signal_25001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8236 ( .C ( clk ), .D ( new_AGEMA_signal_25010 ), .Q ( new_AGEMA_signal_25011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8246 ( .C ( clk ), .D ( new_AGEMA_signal_25020 ), .Q ( new_AGEMA_signal_25021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8256 ( .C ( clk ), .D ( new_AGEMA_signal_25030 ), .Q ( new_AGEMA_signal_25031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8266 ( .C ( clk ), .D ( new_AGEMA_signal_25040 ), .Q ( new_AGEMA_signal_25041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8270 ( .C ( clk ), .D ( new_AGEMA_signal_25044 ), .Q ( new_AGEMA_signal_25045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8274 ( .C ( clk ), .D ( new_AGEMA_signal_25048 ), .Q ( new_AGEMA_signal_25049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8278 ( .C ( clk ), .D ( new_AGEMA_signal_25052 ), .Q ( new_AGEMA_signal_25053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8282 ( .C ( clk ), .D ( new_AGEMA_signal_25056 ), .Q ( new_AGEMA_signal_25057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8286 ( .C ( clk ), .D ( new_AGEMA_signal_25060 ), .Q ( new_AGEMA_signal_25061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8294 ( .C ( clk ), .D ( new_AGEMA_signal_25068 ), .Q ( new_AGEMA_signal_25069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8302 ( .C ( clk ), .D ( new_AGEMA_signal_25076 ), .Q ( new_AGEMA_signal_25077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8310 ( .C ( clk ), .D ( new_AGEMA_signal_25084 ), .Q ( new_AGEMA_signal_25085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8318 ( .C ( clk ), .D ( new_AGEMA_signal_25092 ), .Q ( new_AGEMA_signal_25093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8326 ( .C ( clk ), .D ( new_AGEMA_signal_25100 ), .Q ( new_AGEMA_signal_25101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8330 ( .C ( clk ), .D ( new_AGEMA_signal_25104 ), .Q ( new_AGEMA_signal_25105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8336 ( .C ( clk ), .D ( new_AGEMA_signal_25110 ), .Q ( new_AGEMA_signal_25111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8342 ( .C ( clk ), .D ( new_AGEMA_signal_25116 ), .Q ( new_AGEMA_signal_25117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8348 ( .C ( clk ), .D ( new_AGEMA_signal_25122 ), .Q ( new_AGEMA_signal_25123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8354 ( .C ( clk ), .D ( new_AGEMA_signal_25128 ), .Q ( new_AGEMA_signal_25129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8360 ( .C ( clk ), .D ( new_AGEMA_signal_25134 ), .Q ( new_AGEMA_signal_25135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8366 ( .C ( clk ), .D ( new_AGEMA_signal_25140 ), .Q ( new_AGEMA_signal_25141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8372 ( .C ( clk ), .D ( new_AGEMA_signal_25146 ), .Q ( new_AGEMA_signal_25147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8378 ( .C ( clk ), .D ( new_AGEMA_signal_25152 ), .Q ( new_AGEMA_signal_25153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8384 ( .C ( clk ), .D ( new_AGEMA_signal_25158 ), .Q ( new_AGEMA_signal_25159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8400 ( .C ( clk ), .D ( new_AGEMA_signal_25174 ), .Q ( new_AGEMA_signal_25175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8416 ( .C ( clk ), .D ( new_AGEMA_signal_25190 ), .Q ( new_AGEMA_signal_25191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8432 ( .C ( clk ), .D ( new_AGEMA_signal_25206 ), .Q ( new_AGEMA_signal_25207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8448 ( .C ( clk ), .D ( new_AGEMA_signal_25222 ), .Q ( new_AGEMA_signal_25223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8464 ( .C ( clk ), .D ( new_AGEMA_signal_25238 ), .Q ( new_AGEMA_signal_25239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8474 ( .C ( clk ), .D ( new_AGEMA_signal_25248 ), .Q ( new_AGEMA_signal_25249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8484 ( .C ( clk ), .D ( new_AGEMA_signal_25258 ), .Q ( new_AGEMA_signal_25259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8494 ( .C ( clk ), .D ( new_AGEMA_signal_25268 ), .Q ( new_AGEMA_signal_25269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8504 ( .C ( clk ), .D ( new_AGEMA_signal_25278 ), .Q ( new_AGEMA_signal_25279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8514 ( .C ( clk ), .D ( new_AGEMA_signal_25288 ), .Q ( new_AGEMA_signal_25289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8532 ( .C ( clk ), .D ( new_AGEMA_signal_25306 ), .Q ( new_AGEMA_signal_25307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8550 ( .C ( clk ), .D ( new_AGEMA_signal_25324 ), .Q ( new_AGEMA_signal_25325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8568 ( .C ( clk ), .D ( new_AGEMA_signal_25342 ), .Q ( new_AGEMA_signal_25343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8586 ( .C ( clk ), .D ( new_AGEMA_signal_25360 ), .Q ( new_AGEMA_signal_25361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8604 ( .C ( clk ), .D ( new_AGEMA_signal_25378 ), .Q ( new_AGEMA_signal_25379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8608 ( .C ( clk ), .D ( new_AGEMA_signal_25382 ), .Q ( new_AGEMA_signal_25383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8612 ( .C ( clk ), .D ( new_AGEMA_signal_25386 ), .Q ( new_AGEMA_signal_25387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8616 ( .C ( clk ), .D ( new_AGEMA_signal_25390 ), .Q ( new_AGEMA_signal_25391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8620 ( .C ( clk ), .D ( new_AGEMA_signal_25394 ), .Q ( new_AGEMA_signal_25395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8624 ( .C ( clk ), .D ( new_AGEMA_signal_25398 ), .Q ( new_AGEMA_signal_25399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8632 ( .C ( clk ), .D ( new_AGEMA_signal_25406 ), .Q ( new_AGEMA_signal_25407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8640 ( .C ( clk ), .D ( new_AGEMA_signal_25414 ), .Q ( new_AGEMA_signal_25415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8648 ( .C ( clk ), .D ( new_AGEMA_signal_25422 ), .Q ( new_AGEMA_signal_25423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8656 ( .C ( clk ), .D ( new_AGEMA_signal_25430 ), .Q ( new_AGEMA_signal_25431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8664 ( .C ( clk ), .D ( new_AGEMA_signal_25438 ), .Q ( new_AGEMA_signal_25439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8668 ( .C ( clk ), .D ( new_AGEMA_signal_25442 ), .Q ( new_AGEMA_signal_25443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8672 ( .C ( clk ), .D ( new_AGEMA_signal_25446 ), .Q ( new_AGEMA_signal_25447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8676 ( .C ( clk ), .D ( new_AGEMA_signal_25450 ), .Q ( new_AGEMA_signal_25451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8680 ( .C ( clk ), .D ( new_AGEMA_signal_25454 ), .Q ( new_AGEMA_signal_25455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8684 ( .C ( clk ), .D ( new_AGEMA_signal_25458 ), .Q ( new_AGEMA_signal_25459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8690 ( .C ( clk ), .D ( new_AGEMA_signal_25464 ), .Q ( new_AGEMA_signal_25465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8698 ( .C ( clk ), .D ( new_AGEMA_signal_25472 ), .Q ( new_AGEMA_signal_25473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8706 ( .C ( clk ), .D ( new_AGEMA_signal_25480 ), .Q ( new_AGEMA_signal_25481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8714 ( .C ( clk ), .D ( new_AGEMA_signal_25488 ), .Q ( new_AGEMA_signal_25489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8722 ( .C ( clk ), .D ( new_AGEMA_signal_25496 ), .Q ( new_AGEMA_signal_25497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8728 ( .C ( clk ), .D ( new_AGEMA_signal_25502 ), .Q ( new_AGEMA_signal_25503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8734 ( .C ( clk ), .D ( new_AGEMA_signal_25508 ), .Q ( new_AGEMA_signal_25509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8740 ( .C ( clk ), .D ( new_AGEMA_signal_25514 ), .Q ( new_AGEMA_signal_25515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8746 ( .C ( clk ), .D ( new_AGEMA_signal_25520 ), .Q ( new_AGEMA_signal_25521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8752 ( .C ( clk ), .D ( new_AGEMA_signal_25526 ), .Q ( new_AGEMA_signal_25527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8782 ( .C ( clk ), .D ( new_AGEMA_signal_25556 ), .Q ( new_AGEMA_signal_25557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8802 ( .C ( clk ), .D ( new_AGEMA_signal_25576 ), .Q ( new_AGEMA_signal_25577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8822 ( .C ( clk ), .D ( new_AGEMA_signal_25596 ), .Q ( new_AGEMA_signal_25597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8842 ( .C ( clk ), .D ( new_AGEMA_signal_25616 ), .Q ( new_AGEMA_signal_25617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8862 ( .C ( clk ), .D ( new_AGEMA_signal_25636 ), .Q ( new_AGEMA_signal_25637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8868 ( .C ( clk ), .D ( new_AGEMA_signal_25642 ), .Q ( new_AGEMA_signal_25643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8876 ( .C ( clk ), .D ( new_AGEMA_signal_25650 ), .Q ( new_AGEMA_signal_25651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8884 ( .C ( clk ), .D ( new_AGEMA_signal_25658 ), .Q ( new_AGEMA_signal_25659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8892 ( .C ( clk ), .D ( new_AGEMA_signal_25666 ), .Q ( new_AGEMA_signal_25667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8900 ( .C ( clk ), .D ( new_AGEMA_signal_25674 ), .Q ( new_AGEMA_signal_25675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8912 ( .C ( clk ), .D ( new_AGEMA_signal_25686 ), .Q ( new_AGEMA_signal_25687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8924 ( .C ( clk ), .D ( new_AGEMA_signal_25698 ), .Q ( new_AGEMA_signal_25699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8936 ( .C ( clk ), .D ( new_AGEMA_signal_25710 ), .Q ( new_AGEMA_signal_25711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8948 ( .C ( clk ), .D ( new_AGEMA_signal_25722 ), .Q ( new_AGEMA_signal_25723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8960 ( .C ( clk ), .D ( new_AGEMA_signal_25734 ), .Q ( new_AGEMA_signal_25735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8972 ( .C ( clk ), .D ( new_AGEMA_signal_25746 ), .Q ( new_AGEMA_signal_25747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8986 ( .C ( clk ), .D ( new_AGEMA_signal_25760 ), .Q ( new_AGEMA_signal_25761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9000 ( .C ( clk ), .D ( new_AGEMA_signal_25774 ), .Q ( new_AGEMA_signal_25775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9014 ( .C ( clk ), .D ( new_AGEMA_signal_25788 ), .Q ( new_AGEMA_signal_25789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9028 ( .C ( clk ), .D ( new_AGEMA_signal_25802 ), .Q ( new_AGEMA_signal_25803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9040 ( .C ( clk ), .D ( new_AGEMA_signal_25814 ), .Q ( new_AGEMA_signal_25815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9054 ( .C ( clk ), .D ( new_AGEMA_signal_25828 ), .Q ( new_AGEMA_signal_25829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9068 ( .C ( clk ), .D ( new_AGEMA_signal_25842 ), .Q ( new_AGEMA_signal_25843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9082 ( .C ( clk ), .D ( new_AGEMA_signal_25856 ), .Q ( new_AGEMA_signal_25857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9096 ( .C ( clk ), .D ( new_AGEMA_signal_25870 ), .Q ( new_AGEMA_signal_25871 ) ) ;

    /* cells in depth 23 */
    buf_clk new_AGEMA_reg_buffer_8331 ( .C ( clk ), .D ( new_AGEMA_signal_25105 ), .Q ( new_AGEMA_signal_25106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8337 ( .C ( clk ), .D ( new_AGEMA_signal_25111 ), .Q ( new_AGEMA_signal_25112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8343 ( .C ( clk ), .D ( new_AGEMA_signal_25117 ), .Q ( new_AGEMA_signal_25118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8349 ( .C ( clk ), .D ( new_AGEMA_signal_25123 ), .Q ( new_AGEMA_signal_25124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8355 ( .C ( clk ), .D ( new_AGEMA_signal_25129 ), .Q ( new_AGEMA_signal_25130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8361 ( .C ( clk ), .D ( new_AGEMA_signal_25135 ), .Q ( new_AGEMA_signal_25136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8367 ( .C ( clk ), .D ( new_AGEMA_signal_25141 ), .Q ( new_AGEMA_signal_25142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8373 ( .C ( clk ), .D ( new_AGEMA_signal_25147 ), .Q ( new_AGEMA_signal_25148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8379 ( .C ( clk ), .D ( new_AGEMA_signal_25153 ), .Q ( new_AGEMA_signal_25154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8385 ( .C ( clk ), .D ( new_AGEMA_signal_25159 ), .Q ( new_AGEMA_signal_25160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8401 ( .C ( clk ), .D ( new_AGEMA_signal_25175 ), .Q ( new_AGEMA_signal_25176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8417 ( .C ( clk ), .D ( new_AGEMA_signal_25191 ), .Q ( new_AGEMA_signal_25192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8433 ( .C ( clk ), .D ( new_AGEMA_signal_25207 ), .Q ( new_AGEMA_signal_25208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8449 ( .C ( clk ), .D ( new_AGEMA_signal_25223 ), .Q ( new_AGEMA_signal_25224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8465 ( .C ( clk ), .D ( new_AGEMA_signal_25239 ), .Q ( new_AGEMA_signal_25240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8475 ( .C ( clk ), .D ( new_AGEMA_signal_25249 ), .Q ( new_AGEMA_signal_25250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8485 ( .C ( clk ), .D ( new_AGEMA_signal_25259 ), .Q ( new_AGEMA_signal_25260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8495 ( .C ( clk ), .D ( new_AGEMA_signal_25269 ), .Q ( new_AGEMA_signal_25270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8505 ( .C ( clk ), .D ( new_AGEMA_signal_25279 ), .Q ( new_AGEMA_signal_25280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8515 ( .C ( clk ), .D ( new_AGEMA_signal_25289 ), .Q ( new_AGEMA_signal_25290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8533 ( .C ( clk ), .D ( new_AGEMA_signal_25307 ), .Q ( new_AGEMA_signal_25308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8551 ( .C ( clk ), .D ( new_AGEMA_signal_25325 ), .Q ( new_AGEMA_signal_25326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8569 ( .C ( clk ), .D ( new_AGEMA_signal_25343 ), .Q ( new_AGEMA_signal_25344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8587 ( .C ( clk ), .D ( new_AGEMA_signal_25361 ), .Q ( new_AGEMA_signal_25362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8605 ( .C ( clk ), .D ( new_AGEMA_signal_25379 ), .Q ( new_AGEMA_signal_25380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8609 ( .C ( clk ), .D ( new_AGEMA_signal_25383 ), .Q ( new_AGEMA_signal_25384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8613 ( .C ( clk ), .D ( new_AGEMA_signal_25387 ), .Q ( new_AGEMA_signal_25388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8617 ( .C ( clk ), .D ( new_AGEMA_signal_25391 ), .Q ( new_AGEMA_signal_25392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8621 ( .C ( clk ), .D ( new_AGEMA_signal_25395 ), .Q ( new_AGEMA_signal_25396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8625 ( .C ( clk ), .D ( new_AGEMA_signal_25399 ), .Q ( new_AGEMA_signal_25400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8633 ( .C ( clk ), .D ( new_AGEMA_signal_25407 ), .Q ( new_AGEMA_signal_25408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8641 ( .C ( clk ), .D ( new_AGEMA_signal_25415 ), .Q ( new_AGEMA_signal_25416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8649 ( .C ( clk ), .D ( new_AGEMA_signal_25423 ), .Q ( new_AGEMA_signal_25424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8657 ( .C ( clk ), .D ( new_AGEMA_signal_25431 ), .Q ( new_AGEMA_signal_25432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8665 ( .C ( clk ), .D ( new_AGEMA_signal_25439 ), .Q ( new_AGEMA_signal_25440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8669 ( .C ( clk ), .D ( new_AGEMA_signal_25443 ), .Q ( new_AGEMA_signal_25444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8673 ( .C ( clk ), .D ( new_AGEMA_signal_25447 ), .Q ( new_AGEMA_signal_25448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8677 ( .C ( clk ), .D ( new_AGEMA_signal_25451 ), .Q ( new_AGEMA_signal_25452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8681 ( .C ( clk ), .D ( new_AGEMA_signal_25455 ), .Q ( new_AGEMA_signal_25456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8685 ( .C ( clk ), .D ( new_AGEMA_signal_25459 ), .Q ( new_AGEMA_signal_25460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8691 ( .C ( clk ), .D ( new_AGEMA_signal_25465 ), .Q ( new_AGEMA_signal_25466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8699 ( .C ( clk ), .D ( new_AGEMA_signal_25473 ), .Q ( new_AGEMA_signal_25474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8707 ( .C ( clk ), .D ( new_AGEMA_signal_25481 ), .Q ( new_AGEMA_signal_25482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8715 ( .C ( clk ), .D ( new_AGEMA_signal_25489 ), .Q ( new_AGEMA_signal_25490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8723 ( .C ( clk ), .D ( new_AGEMA_signal_25497 ), .Q ( new_AGEMA_signal_25498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8729 ( .C ( clk ), .D ( new_AGEMA_signal_25503 ), .Q ( new_AGEMA_signal_25504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8735 ( .C ( clk ), .D ( new_AGEMA_signal_25509 ), .Q ( new_AGEMA_signal_25510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8741 ( .C ( clk ), .D ( new_AGEMA_signal_25515 ), .Q ( new_AGEMA_signal_25516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8747 ( .C ( clk ), .D ( new_AGEMA_signal_25521 ), .Q ( new_AGEMA_signal_25522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8753 ( .C ( clk ), .D ( new_AGEMA_signal_25527 ), .Q ( new_AGEMA_signal_25528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8783 ( .C ( clk ), .D ( new_AGEMA_signal_25557 ), .Q ( new_AGEMA_signal_25558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8803 ( .C ( clk ), .D ( new_AGEMA_signal_25577 ), .Q ( new_AGEMA_signal_25578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8823 ( .C ( clk ), .D ( new_AGEMA_signal_25597 ), .Q ( new_AGEMA_signal_25598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8843 ( .C ( clk ), .D ( new_AGEMA_signal_25617 ), .Q ( new_AGEMA_signal_25618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8863 ( .C ( clk ), .D ( new_AGEMA_signal_25637 ), .Q ( new_AGEMA_signal_25638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8869 ( .C ( clk ), .D ( new_AGEMA_signal_25643 ), .Q ( new_AGEMA_signal_25644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8877 ( .C ( clk ), .D ( new_AGEMA_signal_25651 ), .Q ( new_AGEMA_signal_25652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8885 ( .C ( clk ), .D ( new_AGEMA_signal_25659 ), .Q ( new_AGEMA_signal_25660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8893 ( .C ( clk ), .D ( new_AGEMA_signal_25667 ), .Q ( new_AGEMA_signal_25668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8901 ( .C ( clk ), .D ( new_AGEMA_signal_25675 ), .Q ( new_AGEMA_signal_25676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8913 ( .C ( clk ), .D ( new_AGEMA_signal_25687 ), .Q ( new_AGEMA_signal_25688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8925 ( .C ( clk ), .D ( new_AGEMA_signal_25699 ), .Q ( new_AGEMA_signal_25700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8937 ( .C ( clk ), .D ( new_AGEMA_signal_25711 ), .Q ( new_AGEMA_signal_25712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8949 ( .C ( clk ), .D ( new_AGEMA_signal_25723 ), .Q ( new_AGEMA_signal_25724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8961 ( .C ( clk ), .D ( new_AGEMA_signal_25735 ), .Q ( new_AGEMA_signal_25736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8973 ( .C ( clk ), .D ( new_AGEMA_signal_25747 ), .Q ( new_AGEMA_signal_25748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8987 ( .C ( clk ), .D ( new_AGEMA_signal_25761 ), .Q ( new_AGEMA_signal_25762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9001 ( .C ( clk ), .D ( new_AGEMA_signal_25775 ), .Q ( new_AGEMA_signal_25776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9015 ( .C ( clk ), .D ( new_AGEMA_signal_25789 ), .Q ( new_AGEMA_signal_25790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9029 ( .C ( clk ), .D ( new_AGEMA_signal_25803 ), .Q ( new_AGEMA_signal_25804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9041 ( .C ( clk ), .D ( new_AGEMA_signal_25815 ), .Q ( new_AGEMA_signal_25816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9055 ( .C ( clk ), .D ( new_AGEMA_signal_25829 ), .Q ( new_AGEMA_signal_25830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9069 ( .C ( clk ), .D ( new_AGEMA_signal_25843 ), .Q ( new_AGEMA_signal_25844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9083 ( .C ( clk ), .D ( new_AGEMA_signal_25857 ), .Q ( new_AGEMA_signal_25858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9097 ( .C ( clk ), .D ( new_AGEMA_signal_25871 ), .Q ( new_AGEMA_signal_25872 ) ) ;

    /* cells in depth 24 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2130 ( .ina ({new_AGEMA_signal_24791, new_AGEMA_signal_24787, new_AGEMA_signal_24783, new_AGEMA_signal_24779, new_AGEMA_signal_24775}), .inb ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, new_AGEMA_signal_4518, n2001}), .clk ( clk ), .rnd ({Fresh[12659], Fresh[12658], Fresh[12657], Fresh[12656], Fresh[12655], Fresh[12654], Fresh[12653], Fresh[12652], Fresh[12651], Fresh[12650], Fresh[12649], Fresh[12648], Fresh[12647], Fresh[12646], Fresh[12645]}), .outt ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, new_AGEMA_signal_4554, n2017}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2268 ( .ina ({new_AGEMA_signal_24801, new_AGEMA_signal_24799, new_AGEMA_signal_24797, new_AGEMA_signal_24795, new_AGEMA_signal_24793}), .inb ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, n2108}), .clk ( clk ), .rnd ({Fresh[12674], Fresh[12673], Fresh[12672], Fresh[12671], Fresh[12670], Fresh[12669], Fresh[12668], Fresh[12667], Fresh[12666], Fresh[12665], Fresh[12664], Fresh[12663], Fresh[12662], Fresh[12661], Fresh[12660]}), .outt ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, n2110}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2319 ( .ina ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, new_AGEMA_signal_4527, new_AGEMA_signal_4526, n2153}), .inb ({new_AGEMA_signal_24881, new_AGEMA_signal_24865, new_AGEMA_signal_24849, new_AGEMA_signal_24833, new_AGEMA_signal_24817}), .clk ( clk ), .rnd ({Fresh[12689], Fresh[12688], Fresh[12687], Fresh[12686], Fresh[12685], Fresh[12684], Fresh[12683], Fresh[12682], Fresh[12681], Fresh[12680], Fresh[12679], Fresh[12678], Fresh[12677], Fresh[12676], Fresh[12675]}), .outt ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, new_AGEMA_signal_4563, new_AGEMA_signal_4562, n2154}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2375 ( .ina ({new_AGEMA_signal_24901, new_AGEMA_signal_24897, new_AGEMA_signal_24893, new_AGEMA_signal_24889, new_AGEMA_signal_24885}), .inb ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, new_AGEMA_signal_4530, n2207}), .clk ( clk ), .rnd ({Fresh[12704], Fresh[12703], Fresh[12702], Fresh[12701], Fresh[12700], Fresh[12699], Fresh[12698], Fresh[12697], Fresh[12696], Fresh[12695], Fresh[12694], Fresh[12693], Fresh[12692], Fresh[12691], Fresh[12690]}), .outt ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, new_AGEMA_signal_4566, n2209}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2478 ( .ina ({new_AGEMA_signal_24911, new_AGEMA_signal_24909, new_AGEMA_signal_24907, new_AGEMA_signal_24905, new_AGEMA_signal_24903}), .inb ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, n2309}), .clk ( clk ), .rnd ({Fresh[12719], Fresh[12718], Fresh[12717], Fresh[12716], Fresh[12715], Fresh[12714], Fresh[12713], Fresh[12712], Fresh[12711], Fresh[12710], Fresh[12709], Fresh[12708], Fresh[12707], Fresh[12706], Fresh[12705]}), .outt ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, n2311}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2537 ( .ina ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, new_AGEMA_signal_4539, new_AGEMA_signal_4538, n2373}), .inb ({new_AGEMA_signal_24991, new_AGEMA_signal_24975, new_AGEMA_signal_24959, new_AGEMA_signal_24943, new_AGEMA_signal_24927}), .clk ( clk ), .rnd ({Fresh[12734], Fresh[12733], Fresh[12732], Fresh[12731], Fresh[12730], Fresh[12729], Fresh[12728], Fresh[12727], Fresh[12726], Fresh[12725], Fresh[12724], Fresh[12723], Fresh[12722], Fresh[12721], Fresh[12720]}), .outt ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, new_AGEMA_signal_4575, new_AGEMA_signal_4574, n2374}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2672 ( .ina ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, new_AGEMA_signal_4542, n2528}), .inb ({new_AGEMA_signal_25041, new_AGEMA_signal_25031, new_AGEMA_signal_25021, new_AGEMA_signal_25011, new_AGEMA_signal_25001}), .clk ( clk ), .rnd ({Fresh[12749], Fresh[12748], Fresh[12747], Fresh[12746], Fresh[12745], Fresh[12744], Fresh[12743], Fresh[12742], Fresh[12741], Fresh[12740], Fresh[12739], Fresh[12738], Fresh[12737], Fresh[12736], Fresh[12735]}), .outt ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, new_AGEMA_signal_4578, n2529}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2768 ( .ina ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, n2669}), .inb ({new_AGEMA_signal_25061, new_AGEMA_signal_25057, new_AGEMA_signal_25053, new_AGEMA_signal_25049, new_AGEMA_signal_25045}), .clk ( clk ), .rnd ({Fresh[12764], Fresh[12763], Fresh[12762], Fresh[12761], Fresh[12760], Fresh[12759], Fresh[12758], Fresh[12757], Fresh[12756], Fresh[12755], Fresh[12754], Fresh[12753], Fresh[12752], Fresh[12751], Fresh[12750]}), .outt ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, n2670}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2854 ( .ina ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, new_AGEMA_signal_4515, new_AGEMA_signal_4514, n2830}), .inb ({new_AGEMA_signal_25101, new_AGEMA_signal_25093, new_AGEMA_signal_25085, new_AGEMA_signal_25077, new_AGEMA_signal_25069}), .clk ( clk ), .rnd ({Fresh[12779], Fresh[12778], Fresh[12777], Fresh[12776], Fresh[12775], Fresh[12774], Fresh[12773], Fresh[12772], Fresh[12771], Fresh[12770], Fresh[12769], Fresh[12768], Fresh[12767], Fresh[12766], Fresh[12765]}), .outt ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, new_AGEMA_signal_4551, new_AGEMA_signal_4550, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_8332 ( .C ( clk ), .D ( new_AGEMA_signal_25106 ), .Q ( new_AGEMA_signal_25107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8338 ( .C ( clk ), .D ( new_AGEMA_signal_25112 ), .Q ( new_AGEMA_signal_25113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8344 ( .C ( clk ), .D ( new_AGEMA_signal_25118 ), .Q ( new_AGEMA_signal_25119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8350 ( .C ( clk ), .D ( new_AGEMA_signal_25124 ), .Q ( new_AGEMA_signal_25125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8356 ( .C ( clk ), .D ( new_AGEMA_signal_25130 ), .Q ( new_AGEMA_signal_25131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8362 ( .C ( clk ), .D ( new_AGEMA_signal_25136 ), .Q ( new_AGEMA_signal_25137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8368 ( .C ( clk ), .D ( new_AGEMA_signal_25142 ), .Q ( new_AGEMA_signal_25143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8374 ( .C ( clk ), .D ( new_AGEMA_signal_25148 ), .Q ( new_AGEMA_signal_25149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8380 ( .C ( clk ), .D ( new_AGEMA_signal_25154 ), .Q ( new_AGEMA_signal_25155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8386 ( .C ( clk ), .D ( new_AGEMA_signal_25160 ), .Q ( new_AGEMA_signal_25161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8402 ( .C ( clk ), .D ( new_AGEMA_signal_25176 ), .Q ( new_AGEMA_signal_25177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8418 ( .C ( clk ), .D ( new_AGEMA_signal_25192 ), .Q ( new_AGEMA_signal_25193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8434 ( .C ( clk ), .D ( new_AGEMA_signal_25208 ), .Q ( new_AGEMA_signal_25209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8450 ( .C ( clk ), .D ( new_AGEMA_signal_25224 ), .Q ( new_AGEMA_signal_25225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8466 ( .C ( clk ), .D ( new_AGEMA_signal_25240 ), .Q ( new_AGEMA_signal_25241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8476 ( .C ( clk ), .D ( new_AGEMA_signal_25250 ), .Q ( new_AGEMA_signal_25251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8486 ( .C ( clk ), .D ( new_AGEMA_signal_25260 ), .Q ( new_AGEMA_signal_25261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8496 ( .C ( clk ), .D ( new_AGEMA_signal_25270 ), .Q ( new_AGEMA_signal_25271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8506 ( .C ( clk ), .D ( new_AGEMA_signal_25280 ), .Q ( new_AGEMA_signal_25281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8516 ( .C ( clk ), .D ( new_AGEMA_signal_25290 ), .Q ( new_AGEMA_signal_25291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8534 ( .C ( clk ), .D ( new_AGEMA_signal_25308 ), .Q ( new_AGEMA_signal_25309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8552 ( .C ( clk ), .D ( new_AGEMA_signal_25326 ), .Q ( new_AGEMA_signal_25327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8570 ( .C ( clk ), .D ( new_AGEMA_signal_25344 ), .Q ( new_AGEMA_signal_25345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8588 ( .C ( clk ), .D ( new_AGEMA_signal_25362 ), .Q ( new_AGEMA_signal_25363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8606 ( .C ( clk ), .D ( new_AGEMA_signal_25380 ), .Q ( new_AGEMA_signal_25381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8610 ( .C ( clk ), .D ( new_AGEMA_signal_25384 ), .Q ( new_AGEMA_signal_25385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8614 ( .C ( clk ), .D ( new_AGEMA_signal_25388 ), .Q ( new_AGEMA_signal_25389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8618 ( .C ( clk ), .D ( new_AGEMA_signal_25392 ), .Q ( new_AGEMA_signal_25393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8622 ( .C ( clk ), .D ( new_AGEMA_signal_25396 ), .Q ( new_AGEMA_signal_25397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8626 ( .C ( clk ), .D ( new_AGEMA_signal_25400 ), .Q ( new_AGEMA_signal_25401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8634 ( .C ( clk ), .D ( new_AGEMA_signal_25408 ), .Q ( new_AGEMA_signal_25409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8642 ( .C ( clk ), .D ( new_AGEMA_signal_25416 ), .Q ( new_AGEMA_signal_25417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8650 ( .C ( clk ), .D ( new_AGEMA_signal_25424 ), .Q ( new_AGEMA_signal_25425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8658 ( .C ( clk ), .D ( new_AGEMA_signal_25432 ), .Q ( new_AGEMA_signal_25433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8666 ( .C ( clk ), .D ( new_AGEMA_signal_25440 ), .Q ( new_AGEMA_signal_25441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8670 ( .C ( clk ), .D ( new_AGEMA_signal_25444 ), .Q ( new_AGEMA_signal_25445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8674 ( .C ( clk ), .D ( new_AGEMA_signal_25448 ), .Q ( new_AGEMA_signal_25449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8678 ( .C ( clk ), .D ( new_AGEMA_signal_25452 ), .Q ( new_AGEMA_signal_25453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8682 ( .C ( clk ), .D ( new_AGEMA_signal_25456 ), .Q ( new_AGEMA_signal_25457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8686 ( .C ( clk ), .D ( new_AGEMA_signal_25460 ), .Q ( new_AGEMA_signal_25461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8692 ( .C ( clk ), .D ( new_AGEMA_signal_25466 ), .Q ( new_AGEMA_signal_25467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8700 ( .C ( clk ), .D ( new_AGEMA_signal_25474 ), .Q ( new_AGEMA_signal_25475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8708 ( .C ( clk ), .D ( new_AGEMA_signal_25482 ), .Q ( new_AGEMA_signal_25483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8716 ( .C ( clk ), .D ( new_AGEMA_signal_25490 ), .Q ( new_AGEMA_signal_25491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8724 ( .C ( clk ), .D ( new_AGEMA_signal_25498 ), .Q ( new_AGEMA_signal_25499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8730 ( .C ( clk ), .D ( new_AGEMA_signal_25504 ), .Q ( new_AGEMA_signal_25505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8736 ( .C ( clk ), .D ( new_AGEMA_signal_25510 ), .Q ( new_AGEMA_signal_25511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8742 ( .C ( clk ), .D ( new_AGEMA_signal_25516 ), .Q ( new_AGEMA_signal_25517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8748 ( .C ( clk ), .D ( new_AGEMA_signal_25522 ), .Q ( new_AGEMA_signal_25523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8754 ( .C ( clk ), .D ( new_AGEMA_signal_25528 ), .Q ( new_AGEMA_signal_25529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8784 ( .C ( clk ), .D ( new_AGEMA_signal_25558 ), .Q ( new_AGEMA_signal_25559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8804 ( .C ( clk ), .D ( new_AGEMA_signal_25578 ), .Q ( new_AGEMA_signal_25579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8824 ( .C ( clk ), .D ( new_AGEMA_signal_25598 ), .Q ( new_AGEMA_signal_25599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8844 ( .C ( clk ), .D ( new_AGEMA_signal_25618 ), .Q ( new_AGEMA_signal_25619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8864 ( .C ( clk ), .D ( new_AGEMA_signal_25638 ), .Q ( new_AGEMA_signal_25639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8870 ( .C ( clk ), .D ( new_AGEMA_signal_25644 ), .Q ( new_AGEMA_signal_25645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8878 ( .C ( clk ), .D ( new_AGEMA_signal_25652 ), .Q ( new_AGEMA_signal_25653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8886 ( .C ( clk ), .D ( new_AGEMA_signal_25660 ), .Q ( new_AGEMA_signal_25661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8894 ( .C ( clk ), .D ( new_AGEMA_signal_25668 ), .Q ( new_AGEMA_signal_25669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8902 ( .C ( clk ), .D ( new_AGEMA_signal_25676 ), .Q ( new_AGEMA_signal_25677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8914 ( .C ( clk ), .D ( new_AGEMA_signal_25688 ), .Q ( new_AGEMA_signal_25689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8926 ( .C ( clk ), .D ( new_AGEMA_signal_25700 ), .Q ( new_AGEMA_signal_25701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8938 ( .C ( clk ), .D ( new_AGEMA_signal_25712 ), .Q ( new_AGEMA_signal_25713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8950 ( .C ( clk ), .D ( new_AGEMA_signal_25724 ), .Q ( new_AGEMA_signal_25725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8962 ( .C ( clk ), .D ( new_AGEMA_signal_25736 ), .Q ( new_AGEMA_signal_25737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8974 ( .C ( clk ), .D ( new_AGEMA_signal_25748 ), .Q ( new_AGEMA_signal_25749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8988 ( .C ( clk ), .D ( new_AGEMA_signal_25762 ), .Q ( new_AGEMA_signal_25763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9002 ( .C ( clk ), .D ( new_AGEMA_signal_25776 ), .Q ( new_AGEMA_signal_25777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9016 ( .C ( clk ), .D ( new_AGEMA_signal_25790 ), .Q ( new_AGEMA_signal_25791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9030 ( .C ( clk ), .D ( new_AGEMA_signal_25804 ), .Q ( new_AGEMA_signal_25805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9042 ( .C ( clk ), .D ( new_AGEMA_signal_25816 ), .Q ( new_AGEMA_signal_25817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9056 ( .C ( clk ), .D ( new_AGEMA_signal_25830 ), .Q ( new_AGEMA_signal_25831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9070 ( .C ( clk ), .D ( new_AGEMA_signal_25844 ), .Q ( new_AGEMA_signal_25845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9084 ( .C ( clk ), .D ( new_AGEMA_signal_25858 ), .Q ( new_AGEMA_signal_25859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9098 ( .C ( clk ), .D ( new_AGEMA_signal_25872 ), .Q ( new_AGEMA_signal_25873 ) ) ;

    /* cells in depth 25 */
    buf_clk new_AGEMA_reg_buffer_8693 ( .C ( clk ), .D ( new_AGEMA_signal_25467 ), .Q ( new_AGEMA_signal_25468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8701 ( .C ( clk ), .D ( new_AGEMA_signal_25475 ), .Q ( new_AGEMA_signal_25476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8709 ( .C ( clk ), .D ( new_AGEMA_signal_25483 ), .Q ( new_AGEMA_signal_25484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8717 ( .C ( clk ), .D ( new_AGEMA_signal_25491 ), .Q ( new_AGEMA_signal_25492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8725 ( .C ( clk ), .D ( new_AGEMA_signal_25499 ), .Q ( new_AGEMA_signal_25500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8731 ( .C ( clk ), .D ( new_AGEMA_signal_25505 ), .Q ( new_AGEMA_signal_25506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8737 ( .C ( clk ), .D ( new_AGEMA_signal_25511 ), .Q ( new_AGEMA_signal_25512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8743 ( .C ( clk ), .D ( new_AGEMA_signal_25517 ), .Q ( new_AGEMA_signal_25518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8749 ( .C ( clk ), .D ( new_AGEMA_signal_25523 ), .Q ( new_AGEMA_signal_25524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8755 ( .C ( clk ), .D ( new_AGEMA_signal_25529 ), .Q ( new_AGEMA_signal_25530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8757 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_25532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8759 ( .C ( clk ), .D ( new_AGEMA_signal_4566 ), .Q ( new_AGEMA_signal_25534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8761 ( .C ( clk ), .D ( new_AGEMA_signal_4567 ), .Q ( new_AGEMA_signal_25536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8763 ( .C ( clk ), .D ( new_AGEMA_signal_4568 ), .Q ( new_AGEMA_signal_25538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8765 ( .C ( clk ), .D ( new_AGEMA_signal_4569 ), .Q ( new_AGEMA_signal_25540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8785 ( .C ( clk ), .D ( new_AGEMA_signal_25559 ), .Q ( new_AGEMA_signal_25560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8805 ( .C ( clk ), .D ( new_AGEMA_signal_25579 ), .Q ( new_AGEMA_signal_25580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8825 ( .C ( clk ), .D ( new_AGEMA_signal_25599 ), .Q ( new_AGEMA_signal_25600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8845 ( .C ( clk ), .D ( new_AGEMA_signal_25619 ), .Q ( new_AGEMA_signal_25620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8865 ( .C ( clk ), .D ( new_AGEMA_signal_25639 ), .Q ( new_AGEMA_signal_25640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8871 ( .C ( clk ), .D ( new_AGEMA_signal_25645 ), .Q ( new_AGEMA_signal_25646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8879 ( .C ( clk ), .D ( new_AGEMA_signal_25653 ), .Q ( new_AGEMA_signal_25654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8887 ( .C ( clk ), .D ( new_AGEMA_signal_25661 ), .Q ( new_AGEMA_signal_25662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8895 ( .C ( clk ), .D ( new_AGEMA_signal_25669 ), .Q ( new_AGEMA_signal_25670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8903 ( .C ( clk ), .D ( new_AGEMA_signal_25677 ), .Q ( new_AGEMA_signal_25678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8915 ( .C ( clk ), .D ( new_AGEMA_signal_25689 ), .Q ( new_AGEMA_signal_25690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8927 ( .C ( clk ), .D ( new_AGEMA_signal_25701 ), .Q ( new_AGEMA_signal_25702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8939 ( .C ( clk ), .D ( new_AGEMA_signal_25713 ), .Q ( new_AGEMA_signal_25714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8951 ( .C ( clk ), .D ( new_AGEMA_signal_25725 ), .Q ( new_AGEMA_signal_25726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8963 ( .C ( clk ), .D ( new_AGEMA_signal_25737 ), .Q ( new_AGEMA_signal_25738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8975 ( .C ( clk ), .D ( new_AGEMA_signal_25749 ), .Q ( new_AGEMA_signal_25750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8989 ( .C ( clk ), .D ( new_AGEMA_signal_25763 ), .Q ( new_AGEMA_signal_25764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9003 ( .C ( clk ), .D ( new_AGEMA_signal_25777 ), .Q ( new_AGEMA_signal_25778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9017 ( .C ( clk ), .D ( new_AGEMA_signal_25791 ), .Q ( new_AGEMA_signal_25792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9031 ( .C ( clk ), .D ( new_AGEMA_signal_25805 ), .Q ( new_AGEMA_signal_25806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9043 ( .C ( clk ), .D ( new_AGEMA_signal_25817 ), .Q ( new_AGEMA_signal_25818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9057 ( .C ( clk ), .D ( new_AGEMA_signal_25831 ), .Q ( new_AGEMA_signal_25832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9071 ( .C ( clk ), .D ( new_AGEMA_signal_25845 ), .Q ( new_AGEMA_signal_25846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9085 ( .C ( clk ), .D ( new_AGEMA_signal_25859 ), .Q ( new_AGEMA_signal_25860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9099 ( .C ( clk ), .D ( new_AGEMA_signal_25873 ), .Q ( new_AGEMA_signal_25874 ) ) ;

    /* cells in depth 26 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2155 ( .ina ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, new_AGEMA_signal_4554, n2017}), .inb ({new_AGEMA_signal_25131, new_AGEMA_signal_25125, new_AGEMA_signal_25119, new_AGEMA_signal_25113, new_AGEMA_signal_25107}), .clk ( clk ), .rnd ({Fresh[12794], Fresh[12793], Fresh[12792], Fresh[12791], Fresh[12790], Fresh[12789], Fresh[12788], Fresh[12787], Fresh[12786], Fresh[12785], Fresh[12784], Fresh[12783], Fresh[12782], Fresh[12781], Fresh[12780]}), .outt ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, new_AGEMA_signal_4590, n2018}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2269 ( .ina ({new_AGEMA_signal_25161, new_AGEMA_signal_25155, new_AGEMA_signal_25149, new_AGEMA_signal_25143, new_AGEMA_signal_25137}), .inb ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, n2110}), .clk ( clk ), .rnd ({Fresh[12809], Fresh[12808], Fresh[12807], Fresh[12806], Fresh[12805], Fresh[12804], Fresh[12803], Fresh[12802], Fresh[12801], Fresh[12800], Fresh[12799], Fresh[12798], Fresh[12797], Fresh[12796], Fresh[12795]}), .outt ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, n2112}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2320 ( .ina ({new_AGEMA_signal_25241, new_AGEMA_signal_25225, new_AGEMA_signal_25209, new_AGEMA_signal_25193, new_AGEMA_signal_25177}), .inb ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, new_AGEMA_signal_4563, new_AGEMA_signal_4562, n2154}), .clk ( clk ), .rnd ({Fresh[12824], Fresh[12823], Fresh[12822], Fresh[12821], Fresh[12820], Fresh[12819], Fresh[12818], Fresh[12817], Fresh[12816], Fresh[12815], Fresh[12814], Fresh[12813], Fresh[12812], Fresh[12811], Fresh[12810]}), .outt ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, n2210}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2479 ( .ina ({new_AGEMA_signal_25291, new_AGEMA_signal_25281, new_AGEMA_signal_25271, new_AGEMA_signal_25261, new_AGEMA_signal_25251}), .inb ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, n2311}), .clk ( clk ), .rnd ({Fresh[12839], Fresh[12838], Fresh[12837], Fresh[12836], Fresh[12835], Fresh[12834], Fresh[12833], Fresh[12832], Fresh[12831], Fresh[12830], Fresh[12829], Fresh[12828], Fresh[12827], Fresh[12826], Fresh[12825]}), .outt ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, new_AGEMA_signal_4602, N470}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2538 ( .ina ({new_AGEMA_signal_25381, new_AGEMA_signal_25363, new_AGEMA_signal_25345, new_AGEMA_signal_25327, new_AGEMA_signal_25309}), .inb ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, new_AGEMA_signal_4575, new_AGEMA_signal_4574, n2374}), .clk ( clk ), .rnd ({Fresh[12854], Fresh[12853], Fresh[12852], Fresh[12851], Fresh[12850], Fresh[12849], Fresh[12848], Fresh[12847], Fresh[12846], Fresh[12845], Fresh[12844], Fresh[12843], Fresh[12842], Fresh[12841], Fresh[12840]}), .outt ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, n2378}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2673 ( .ina ({new_AGEMA_signal_25401, new_AGEMA_signal_25397, new_AGEMA_signal_25393, new_AGEMA_signal_25389, new_AGEMA_signal_25385}), .inb ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, new_AGEMA_signal_4578, n2529}), .clk ( clk ), .rnd ({Fresh[12869], Fresh[12868], Fresh[12867], Fresh[12866], Fresh[12865], Fresh[12864], Fresh[12863], Fresh[12862], Fresh[12861], Fresh[12860], Fresh[12859], Fresh[12858], Fresh[12857], Fresh[12856], Fresh[12855]}), .outt ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, new_AGEMA_signal_4611, new_AGEMA_signal_4610, N639}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2769 ( .ina ({new_AGEMA_signal_25441, new_AGEMA_signal_25433, new_AGEMA_signal_25425, new_AGEMA_signal_25417, new_AGEMA_signal_25409}), .inb ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, n2670}), .clk ( clk ), .rnd ({Fresh[12884], Fresh[12883], Fresh[12882], Fresh[12881], Fresh[12880], Fresh[12879], Fresh[12878], Fresh[12877], Fresh[12876], Fresh[12875], Fresh[12874], Fresh[12873], Fresh[12872], Fresh[12871], Fresh[12870]}), .outt ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, new_AGEMA_signal_4614, N723}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2855 ( .ina ({new_AGEMA_signal_25461, new_AGEMA_signal_25457, new_AGEMA_signal_25453, new_AGEMA_signal_25449, new_AGEMA_signal_25445}), .inb ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, new_AGEMA_signal_4551, new_AGEMA_signal_4550, n2831}), .clk ( clk ), .rnd ({Fresh[12899], Fresh[12898], Fresh[12897], Fresh[12896], Fresh[12895], Fresh[12894], Fresh[12893], Fresh[12892], Fresh[12891], Fresh[12890], Fresh[12889], Fresh[12888], Fresh[12887], Fresh[12886], Fresh[12885]}), .outt ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, new_AGEMA_signal_4587, new_AGEMA_signal_4586, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_8694 ( .C ( clk ), .D ( new_AGEMA_signal_25468 ), .Q ( new_AGEMA_signal_25469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8702 ( .C ( clk ), .D ( new_AGEMA_signal_25476 ), .Q ( new_AGEMA_signal_25477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8710 ( .C ( clk ), .D ( new_AGEMA_signal_25484 ), .Q ( new_AGEMA_signal_25485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8718 ( .C ( clk ), .D ( new_AGEMA_signal_25492 ), .Q ( new_AGEMA_signal_25493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8726 ( .C ( clk ), .D ( new_AGEMA_signal_25500 ), .Q ( new_AGEMA_signal_25501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8732 ( .C ( clk ), .D ( new_AGEMA_signal_25506 ), .Q ( new_AGEMA_signal_25507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8738 ( .C ( clk ), .D ( new_AGEMA_signal_25512 ), .Q ( new_AGEMA_signal_25513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8744 ( .C ( clk ), .D ( new_AGEMA_signal_25518 ), .Q ( new_AGEMA_signal_25519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8750 ( .C ( clk ), .D ( new_AGEMA_signal_25524 ), .Q ( new_AGEMA_signal_25525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8756 ( .C ( clk ), .D ( new_AGEMA_signal_25530 ), .Q ( new_AGEMA_signal_25531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8758 ( .C ( clk ), .D ( new_AGEMA_signal_25532 ), .Q ( new_AGEMA_signal_25533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8760 ( .C ( clk ), .D ( new_AGEMA_signal_25534 ), .Q ( new_AGEMA_signal_25535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8762 ( .C ( clk ), .D ( new_AGEMA_signal_25536 ), .Q ( new_AGEMA_signal_25537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8764 ( .C ( clk ), .D ( new_AGEMA_signal_25538 ), .Q ( new_AGEMA_signal_25539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8766 ( .C ( clk ), .D ( new_AGEMA_signal_25540 ), .Q ( new_AGEMA_signal_25541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8786 ( .C ( clk ), .D ( new_AGEMA_signal_25560 ), .Q ( new_AGEMA_signal_25561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8806 ( .C ( clk ), .D ( new_AGEMA_signal_25580 ), .Q ( new_AGEMA_signal_25581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8826 ( .C ( clk ), .D ( new_AGEMA_signal_25600 ), .Q ( new_AGEMA_signal_25601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8846 ( .C ( clk ), .D ( new_AGEMA_signal_25620 ), .Q ( new_AGEMA_signal_25621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8866 ( .C ( clk ), .D ( new_AGEMA_signal_25640 ), .Q ( new_AGEMA_signal_25641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8872 ( .C ( clk ), .D ( new_AGEMA_signal_25646 ), .Q ( new_AGEMA_signal_25647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8880 ( .C ( clk ), .D ( new_AGEMA_signal_25654 ), .Q ( new_AGEMA_signal_25655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8888 ( .C ( clk ), .D ( new_AGEMA_signal_25662 ), .Q ( new_AGEMA_signal_25663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8896 ( .C ( clk ), .D ( new_AGEMA_signal_25670 ), .Q ( new_AGEMA_signal_25671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8904 ( .C ( clk ), .D ( new_AGEMA_signal_25678 ), .Q ( new_AGEMA_signal_25679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8916 ( .C ( clk ), .D ( new_AGEMA_signal_25690 ), .Q ( new_AGEMA_signal_25691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8928 ( .C ( clk ), .D ( new_AGEMA_signal_25702 ), .Q ( new_AGEMA_signal_25703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8940 ( .C ( clk ), .D ( new_AGEMA_signal_25714 ), .Q ( new_AGEMA_signal_25715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8952 ( .C ( clk ), .D ( new_AGEMA_signal_25726 ), .Q ( new_AGEMA_signal_25727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8964 ( .C ( clk ), .D ( new_AGEMA_signal_25738 ), .Q ( new_AGEMA_signal_25739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8976 ( .C ( clk ), .D ( new_AGEMA_signal_25750 ), .Q ( new_AGEMA_signal_25751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8990 ( .C ( clk ), .D ( new_AGEMA_signal_25764 ), .Q ( new_AGEMA_signal_25765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9004 ( .C ( clk ), .D ( new_AGEMA_signal_25778 ), .Q ( new_AGEMA_signal_25779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9018 ( .C ( clk ), .D ( new_AGEMA_signal_25792 ), .Q ( new_AGEMA_signal_25793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9032 ( .C ( clk ), .D ( new_AGEMA_signal_25806 ), .Q ( new_AGEMA_signal_25807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9044 ( .C ( clk ), .D ( new_AGEMA_signal_25818 ), .Q ( new_AGEMA_signal_25819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9058 ( .C ( clk ), .D ( new_AGEMA_signal_25832 ), .Q ( new_AGEMA_signal_25833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9072 ( .C ( clk ), .D ( new_AGEMA_signal_25846 ), .Q ( new_AGEMA_signal_25847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9086 ( .C ( clk ), .D ( new_AGEMA_signal_25860 ), .Q ( new_AGEMA_signal_25861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9100 ( .C ( clk ), .D ( new_AGEMA_signal_25874 ), .Q ( new_AGEMA_signal_25875 ) ) ;

    /* cells in depth 27 */
    buf_clk new_AGEMA_reg_buffer_8873 ( .C ( clk ), .D ( new_AGEMA_signal_25647 ), .Q ( new_AGEMA_signal_25648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8881 ( .C ( clk ), .D ( new_AGEMA_signal_25655 ), .Q ( new_AGEMA_signal_25656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8889 ( .C ( clk ), .D ( new_AGEMA_signal_25663 ), .Q ( new_AGEMA_signal_25664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8897 ( .C ( clk ), .D ( new_AGEMA_signal_25671 ), .Q ( new_AGEMA_signal_25672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8905 ( .C ( clk ), .D ( new_AGEMA_signal_25679 ), .Q ( new_AGEMA_signal_25680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8917 ( .C ( clk ), .D ( new_AGEMA_signal_25691 ), .Q ( new_AGEMA_signal_25692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8929 ( .C ( clk ), .D ( new_AGEMA_signal_25703 ), .Q ( new_AGEMA_signal_25704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8941 ( .C ( clk ), .D ( new_AGEMA_signal_25715 ), .Q ( new_AGEMA_signal_25716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8953 ( .C ( clk ), .D ( new_AGEMA_signal_25727 ), .Q ( new_AGEMA_signal_25728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8965 ( .C ( clk ), .D ( new_AGEMA_signal_25739 ), .Q ( new_AGEMA_signal_25740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8977 ( .C ( clk ), .D ( new_AGEMA_signal_25751 ), .Q ( new_AGEMA_signal_25752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8991 ( .C ( clk ), .D ( new_AGEMA_signal_25765 ), .Q ( new_AGEMA_signal_25766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9005 ( .C ( clk ), .D ( new_AGEMA_signal_25779 ), .Q ( new_AGEMA_signal_25780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9019 ( .C ( clk ), .D ( new_AGEMA_signal_25793 ), .Q ( new_AGEMA_signal_25794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9033 ( .C ( clk ), .D ( new_AGEMA_signal_25807 ), .Q ( new_AGEMA_signal_25808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9045 ( .C ( clk ), .D ( new_AGEMA_signal_25819 ), .Q ( new_AGEMA_signal_25820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9059 ( .C ( clk ), .D ( new_AGEMA_signal_25833 ), .Q ( new_AGEMA_signal_25834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9073 ( .C ( clk ), .D ( new_AGEMA_signal_25847 ), .Q ( new_AGEMA_signal_25848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9087 ( .C ( clk ), .D ( new_AGEMA_signal_25861 ), .Q ( new_AGEMA_signal_25862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9101 ( .C ( clk ), .D ( new_AGEMA_signal_25875 ), .Q ( new_AGEMA_signal_25876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9187 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_25962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9195 ( .C ( clk ), .D ( new_AGEMA_signal_4602 ), .Q ( new_AGEMA_signal_25970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9203 ( .C ( clk ), .D ( new_AGEMA_signal_4603 ), .Q ( new_AGEMA_signal_25978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9211 ( .C ( clk ), .D ( new_AGEMA_signal_4604 ), .Q ( new_AGEMA_signal_25986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9219 ( .C ( clk ), .D ( new_AGEMA_signal_4605 ), .Q ( new_AGEMA_signal_25994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9227 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_26002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9235 ( .C ( clk ), .D ( new_AGEMA_signal_4610 ), .Q ( new_AGEMA_signal_26010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9243 ( .C ( clk ), .D ( new_AGEMA_signal_4611 ), .Q ( new_AGEMA_signal_26018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9251 ( .C ( clk ), .D ( new_AGEMA_signal_4612 ), .Q ( new_AGEMA_signal_26026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9259 ( .C ( clk ), .D ( new_AGEMA_signal_4613 ), .Q ( new_AGEMA_signal_26034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9267 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_26042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9275 ( .C ( clk ), .D ( new_AGEMA_signal_4614 ), .Q ( new_AGEMA_signal_26050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9283 ( .C ( clk ), .D ( new_AGEMA_signal_4615 ), .Q ( new_AGEMA_signal_26058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9291 ( .C ( clk ), .D ( new_AGEMA_signal_4616 ), .Q ( new_AGEMA_signal_26066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9299 ( .C ( clk ), .D ( new_AGEMA_signal_4617 ), .Q ( new_AGEMA_signal_26074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9307 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_26082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9315 ( .C ( clk ), .D ( new_AGEMA_signal_4586 ), .Q ( new_AGEMA_signal_26090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9323 ( .C ( clk ), .D ( new_AGEMA_signal_4587 ), .Q ( new_AGEMA_signal_26098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9331 ( .C ( clk ), .D ( new_AGEMA_signal_4588 ), .Q ( new_AGEMA_signal_26106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9339 ( .C ( clk ), .D ( new_AGEMA_signal_4589 ), .Q ( new_AGEMA_signal_26114 ) ) ;

    /* cells in depth 28 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2156 ( .ina ({new_AGEMA_signal_25501, new_AGEMA_signal_25493, new_AGEMA_signal_25485, new_AGEMA_signal_25477, new_AGEMA_signal_25469}), .inb ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, new_AGEMA_signal_4590, n2018}), .clk ( clk ), .rnd ({Fresh[12914], Fresh[12913], Fresh[12912], Fresh[12911], Fresh[12910], Fresh[12909], Fresh[12908], Fresh[12907], Fresh[12906], Fresh[12905], Fresh[12904], Fresh[12903], Fresh[12902], Fresh[12901], Fresh[12900]}), .outt ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, N169}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2270 ( .ina ({new_AGEMA_signal_25531, new_AGEMA_signal_25525, new_AGEMA_signal_25519, new_AGEMA_signal_25513, new_AGEMA_signal_25507}), .inb ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, n2112}), .clk ( clk ), .rnd ({Fresh[12929], Fresh[12928], Fresh[12927], Fresh[12926], Fresh[12925], Fresh[12924], Fresh[12923], Fresh[12922], Fresh[12921], Fresh[12920], Fresh[12919], Fresh[12918], Fresh[12917], Fresh[12916], Fresh[12915]}), .outt ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, new_AGEMA_signal_4623, new_AGEMA_signal_4622, N277}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2376 ( .ina ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, new_AGEMA_signal_4599, new_AGEMA_signal_4598, n2210}), .inb ({new_AGEMA_signal_25541, new_AGEMA_signal_25539, new_AGEMA_signal_25537, new_AGEMA_signal_25535, new_AGEMA_signal_25533}), .clk ( clk ), .rnd ({Fresh[12944], Fresh[12943], Fresh[12942], Fresh[12941], Fresh[12940], Fresh[12939], Fresh[12938], Fresh[12937], Fresh[12936], Fresh[12935], Fresh[12934], Fresh[12933], Fresh[12932], Fresh[12931], Fresh[12930]}), .outt ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, new_AGEMA_signal_4626, n2211}) ) ;
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2540 ( .ina ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, n2378}), .inb ({new_AGEMA_signal_25641, new_AGEMA_signal_25621, new_AGEMA_signal_25601, new_AGEMA_signal_25581, new_AGEMA_signal_25561}), .clk ( clk ), .rnd ({Fresh[12959], Fresh[12958], Fresh[12957], Fresh[12956], Fresh[12955], Fresh[12954], Fresh[12953], Fresh[12952], Fresh[12951], Fresh[12950], Fresh[12949], Fresh[12948], Fresh[12947], Fresh[12946], Fresh[12945]}), .outt ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_8874 ( .C ( clk ), .D ( new_AGEMA_signal_25648 ), .Q ( new_AGEMA_signal_25649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8882 ( .C ( clk ), .D ( new_AGEMA_signal_25656 ), .Q ( new_AGEMA_signal_25657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8890 ( .C ( clk ), .D ( new_AGEMA_signal_25664 ), .Q ( new_AGEMA_signal_25665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8898 ( .C ( clk ), .D ( new_AGEMA_signal_25672 ), .Q ( new_AGEMA_signal_25673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8906 ( .C ( clk ), .D ( new_AGEMA_signal_25680 ), .Q ( new_AGEMA_signal_25681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8918 ( .C ( clk ), .D ( new_AGEMA_signal_25692 ), .Q ( new_AGEMA_signal_25693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8930 ( .C ( clk ), .D ( new_AGEMA_signal_25704 ), .Q ( new_AGEMA_signal_25705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8942 ( .C ( clk ), .D ( new_AGEMA_signal_25716 ), .Q ( new_AGEMA_signal_25717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8954 ( .C ( clk ), .D ( new_AGEMA_signal_25728 ), .Q ( new_AGEMA_signal_25729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8966 ( .C ( clk ), .D ( new_AGEMA_signal_25740 ), .Q ( new_AGEMA_signal_25741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8978 ( .C ( clk ), .D ( new_AGEMA_signal_25752 ), .Q ( new_AGEMA_signal_25753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8992 ( .C ( clk ), .D ( new_AGEMA_signal_25766 ), .Q ( new_AGEMA_signal_25767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9006 ( .C ( clk ), .D ( new_AGEMA_signal_25780 ), .Q ( new_AGEMA_signal_25781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9020 ( .C ( clk ), .D ( new_AGEMA_signal_25794 ), .Q ( new_AGEMA_signal_25795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9034 ( .C ( clk ), .D ( new_AGEMA_signal_25808 ), .Q ( new_AGEMA_signal_25809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9046 ( .C ( clk ), .D ( new_AGEMA_signal_25820 ), .Q ( new_AGEMA_signal_25821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9060 ( .C ( clk ), .D ( new_AGEMA_signal_25834 ), .Q ( new_AGEMA_signal_25835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9074 ( .C ( clk ), .D ( new_AGEMA_signal_25848 ), .Q ( new_AGEMA_signal_25849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9088 ( .C ( clk ), .D ( new_AGEMA_signal_25862 ), .Q ( new_AGEMA_signal_25863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9102 ( .C ( clk ), .D ( new_AGEMA_signal_25876 ), .Q ( new_AGEMA_signal_25877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9188 ( .C ( clk ), .D ( new_AGEMA_signal_25962 ), .Q ( new_AGEMA_signal_25963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9196 ( .C ( clk ), .D ( new_AGEMA_signal_25970 ), .Q ( new_AGEMA_signal_25971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9204 ( .C ( clk ), .D ( new_AGEMA_signal_25978 ), .Q ( new_AGEMA_signal_25979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9212 ( .C ( clk ), .D ( new_AGEMA_signal_25986 ), .Q ( new_AGEMA_signal_25987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9220 ( .C ( clk ), .D ( new_AGEMA_signal_25994 ), .Q ( new_AGEMA_signal_25995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9228 ( .C ( clk ), .D ( new_AGEMA_signal_26002 ), .Q ( new_AGEMA_signal_26003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9236 ( .C ( clk ), .D ( new_AGEMA_signal_26010 ), .Q ( new_AGEMA_signal_26011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9244 ( .C ( clk ), .D ( new_AGEMA_signal_26018 ), .Q ( new_AGEMA_signal_26019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9252 ( .C ( clk ), .D ( new_AGEMA_signal_26026 ), .Q ( new_AGEMA_signal_26027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9260 ( .C ( clk ), .D ( new_AGEMA_signal_26034 ), .Q ( new_AGEMA_signal_26035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9268 ( .C ( clk ), .D ( new_AGEMA_signal_26042 ), .Q ( new_AGEMA_signal_26043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9276 ( .C ( clk ), .D ( new_AGEMA_signal_26050 ), .Q ( new_AGEMA_signal_26051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9284 ( .C ( clk ), .D ( new_AGEMA_signal_26058 ), .Q ( new_AGEMA_signal_26059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9292 ( .C ( clk ), .D ( new_AGEMA_signal_26066 ), .Q ( new_AGEMA_signal_26067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9300 ( .C ( clk ), .D ( new_AGEMA_signal_26074 ), .Q ( new_AGEMA_signal_26075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9308 ( .C ( clk ), .D ( new_AGEMA_signal_26082 ), .Q ( new_AGEMA_signal_26083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9316 ( .C ( clk ), .D ( new_AGEMA_signal_26090 ), .Q ( new_AGEMA_signal_26091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9324 ( .C ( clk ), .D ( new_AGEMA_signal_26098 ), .Q ( new_AGEMA_signal_26099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9332 ( .C ( clk ), .D ( new_AGEMA_signal_26106 ), .Q ( new_AGEMA_signal_26107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9340 ( .C ( clk ), .D ( new_AGEMA_signal_26114 ), .Q ( new_AGEMA_signal_26115 ) ) ;

    /* cells in depth 29 */
    buf_clk new_AGEMA_reg_buffer_8979 ( .C ( clk ), .D ( new_AGEMA_signal_25753 ), .Q ( new_AGEMA_signal_25754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8993 ( .C ( clk ), .D ( new_AGEMA_signal_25767 ), .Q ( new_AGEMA_signal_25768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9007 ( .C ( clk ), .D ( new_AGEMA_signal_25781 ), .Q ( new_AGEMA_signal_25782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9021 ( .C ( clk ), .D ( new_AGEMA_signal_25795 ), .Q ( new_AGEMA_signal_25796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9035 ( .C ( clk ), .D ( new_AGEMA_signal_25809 ), .Q ( new_AGEMA_signal_25810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9047 ( .C ( clk ), .D ( new_AGEMA_signal_25821 ), .Q ( new_AGEMA_signal_25822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9061 ( .C ( clk ), .D ( new_AGEMA_signal_25835 ), .Q ( new_AGEMA_signal_25836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9075 ( .C ( clk ), .D ( new_AGEMA_signal_25849 ), .Q ( new_AGEMA_signal_25850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9089 ( .C ( clk ), .D ( new_AGEMA_signal_25863 ), .Q ( new_AGEMA_signal_25864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9103 ( .C ( clk ), .D ( new_AGEMA_signal_25877 ), .Q ( new_AGEMA_signal_25878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9107 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_25882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9113 ( .C ( clk ), .D ( new_AGEMA_signal_4618 ), .Q ( new_AGEMA_signal_25888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9119 ( .C ( clk ), .D ( new_AGEMA_signal_4619 ), .Q ( new_AGEMA_signal_25894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9125 ( .C ( clk ), .D ( new_AGEMA_signal_4620 ), .Q ( new_AGEMA_signal_25900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9131 ( .C ( clk ), .D ( new_AGEMA_signal_4621 ), .Q ( new_AGEMA_signal_25906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9137 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_25912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9143 ( .C ( clk ), .D ( new_AGEMA_signal_4622 ), .Q ( new_AGEMA_signal_25918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9149 ( .C ( clk ), .D ( new_AGEMA_signal_4623 ), .Q ( new_AGEMA_signal_25924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9155 ( .C ( clk ), .D ( new_AGEMA_signal_4624 ), .Q ( new_AGEMA_signal_25930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9161 ( .C ( clk ), .D ( new_AGEMA_signal_4625 ), .Q ( new_AGEMA_signal_25936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9189 ( .C ( clk ), .D ( new_AGEMA_signal_25963 ), .Q ( new_AGEMA_signal_25964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9197 ( .C ( clk ), .D ( new_AGEMA_signal_25971 ), .Q ( new_AGEMA_signal_25972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9205 ( .C ( clk ), .D ( new_AGEMA_signal_25979 ), .Q ( new_AGEMA_signal_25980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9213 ( .C ( clk ), .D ( new_AGEMA_signal_25987 ), .Q ( new_AGEMA_signal_25988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9221 ( .C ( clk ), .D ( new_AGEMA_signal_25995 ), .Q ( new_AGEMA_signal_25996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9229 ( .C ( clk ), .D ( new_AGEMA_signal_26003 ), .Q ( new_AGEMA_signal_26004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9237 ( .C ( clk ), .D ( new_AGEMA_signal_26011 ), .Q ( new_AGEMA_signal_26012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9245 ( .C ( clk ), .D ( new_AGEMA_signal_26019 ), .Q ( new_AGEMA_signal_26020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9253 ( .C ( clk ), .D ( new_AGEMA_signal_26027 ), .Q ( new_AGEMA_signal_26028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9261 ( .C ( clk ), .D ( new_AGEMA_signal_26035 ), .Q ( new_AGEMA_signal_26036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9269 ( .C ( clk ), .D ( new_AGEMA_signal_26043 ), .Q ( new_AGEMA_signal_26044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9277 ( .C ( clk ), .D ( new_AGEMA_signal_26051 ), .Q ( new_AGEMA_signal_26052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9285 ( .C ( clk ), .D ( new_AGEMA_signal_26059 ), .Q ( new_AGEMA_signal_26060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9293 ( .C ( clk ), .D ( new_AGEMA_signal_26067 ), .Q ( new_AGEMA_signal_26068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9301 ( .C ( clk ), .D ( new_AGEMA_signal_26075 ), .Q ( new_AGEMA_signal_26076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9309 ( .C ( clk ), .D ( new_AGEMA_signal_26083 ), .Q ( new_AGEMA_signal_26084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9317 ( .C ( clk ), .D ( new_AGEMA_signal_26091 ), .Q ( new_AGEMA_signal_26092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9325 ( .C ( clk ), .D ( new_AGEMA_signal_26099 ), .Q ( new_AGEMA_signal_26100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9333 ( .C ( clk ), .D ( new_AGEMA_signal_26107 ), .Q ( new_AGEMA_signal_26108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9341 ( .C ( clk ), .D ( new_AGEMA_signal_26115 ), .Q ( new_AGEMA_signal_26116 ) ) ;

    /* cells in depth 30 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2377 ( .ina ({new_AGEMA_signal_25681, new_AGEMA_signal_25673, new_AGEMA_signal_25665, new_AGEMA_signal_25657, new_AGEMA_signal_25649}), .inb ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, new_AGEMA_signal_4626, n2211}), .clk ( clk ), .rnd ({Fresh[12974], Fresh[12973], Fresh[12972], Fresh[12971], Fresh[12970], Fresh[12969], Fresh[12968], Fresh[12967], Fresh[12966], Fresh[12965], Fresh[12964], Fresh[12963], Fresh[12962], Fresh[12961], Fresh[12960]}), .outt ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, new_AGEMA_signal_4635, new_AGEMA_signal_4634, N379}) ) ;
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2541 ( .ina ({new_AGEMA_signal_25741, new_AGEMA_signal_25729, new_AGEMA_signal_25717, new_AGEMA_signal_25705, new_AGEMA_signal_25693}), .inb ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, n2379}), .clk ( clk ), .rnd ({Fresh[12989], Fresh[12988], Fresh[12987], Fresh[12986], Fresh[12985], Fresh[12984], Fresh[12983], Fresh[12982], Fresh[12981], Fresh[12980], Fresh[12979], Fresh[12978], Fresh[12977], Fresh[12976], Fresh[12975]}), .outt ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, new_AGEMA_signal_4638, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_8980 ( .C ( clk ), .D ( new_AGEMA_signal_25754 ), .Q ( new_AGEMA_signal_25755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_8994 ( .C ( clk ), .D ( new_AGEMA_signal_25768 ), .Q ( new_AGEMA_signal_25769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9008 ( .C ( clk ), .D ( new_AGEMA_signal_25782 ), .Q ( new_AGEMA_signal_25783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9022 ( .C ( clk ), .D ( new_AGEMA_signal_25796 ), .Q ( new_AGEMA_signal_25797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9036 ( .C ( clk ), .D ( new_AGEMA_signal_25810 ), .Q ( new_AGEMA_signal_25811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9048 ( .C ( clk ), .D ( new_AGEMA_signal_25822 ), .Q ( new_AGEMA_signal_25823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9062 ( .C ( clk ), .D ( new_AGEMA_signal_25836 ), .Q ( new_AGEMA_signal_25837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9076 ( .C ( clk ), .D ( new_AGEMA_signal_25850 ), .Q ( new_AGEMA_signal_25851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9090 ( .C ( clk ), .D ( new_AGEMA_signal_25864 ), .Q ( new_AGEMA_signal_25865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9104 ( .C ( clk ), .D ( new_AGEMA_signal_25878 ), .Q ( new_AGEMA_signal_25879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9108 ( .C ( clk ), .D ( new_AGEMA_signal_25882 ), .Q ( new_AGEMA_signal_25883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9114 ( .C ( clk ), .D ( new_AGEMA_signal_25888 ), .Q ( new_AGEMA_signal_25889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9120 ( .C ( clk ), .D ( new_AGEMA_signal_25894 ), .Q ( new_AGEMA_signal_25895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9126 ( .C ( clk ), .D ( new_AGEMA_signal_25900 ), .Q ( new_AGEMA_signal_25901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9132 ( .C ( clk ), .D ( new_AGEMA_signal_25906 ), .Q ( new_AGEMA_signal_25907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9138 ( .C ( clk ), .D ( new_AGEMA_signal_25912 ), .Q ( new_AGEMA_signal_25913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9144 ( .C ( clk ), .D ( new_AGEMA_signal_25918 ), .Q ( new_AGEMA_signal_25919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9150 ( .C ( clk ), .D ( new_AGEMA_signal_25924 ), .Q ( new_AGEMA_signal_25925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9156 ( .C ( clk ), .D ( new_AGEMA_signal_25930 ), .Q ( new_AGEMA_signal_25931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9162 ( .C ( clk ), .D ( new_AGEMA_signal_25936 ), .Q ( new_AGEMA_signal_25937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9190 ( .C ( clk ), .D ( new_AGEMA_signal_25964 ), .Q ( new_AGEMA_signal_25965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9198 ( .C ( clk ), .D ( new_AGEMA_signal_25972 ), .Q ( new_AGEMA_signal_25973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9206 ( .C ( clk ), .D ( new_AGEMA_signal_25980 ), .Q ( new_AGEMA_signal_25981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9214 ( .C ( clk ), .D ( new_AGEMA_signal_25988 ), .Q ( new_AGEMA_signal_25989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9222 ( .C ( clk ), .D ( new_AGEMA_signal_25996 ), .Q ( new_AGEMA_signal_25997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9230 ( .C ( clk ), .D ( new_AGEMA_signal_26004 ), .Q ( new_AGEMA_signal_26005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9238 ( .C ( clk ), .D ( new_AGEMA_signal_26012 ), .Q ( new_AGEMA_signal_26013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9246 ( .C ( clk ), .D ( new_AGEMA_signal_26020 ), .Q ( new_AGEMA_signal_26021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9254 ( .C ( clk ), .D ( new_AGEMA_signal_26028 ), .Q ( new_AGEMA_signal_26029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9262 ( .C ( clk ), .D ( new_AGEMA_signal_26036 ), .Q ( new_AGEMA_signal_26037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9270 ( .C ( clk ), .D ( new_AGEMA_signal_26044 ), .Q ( new_AGEMA_signal_26045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9278 ( .C ( clk ), .D ( new_AGEMA_signal_26052 ), .Q ( new_AGEMA_signal_26053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9286 ( .C ( clk ), .D ( new_AGEMA_signal_26060 ), .Q ( new_AGEMA_signal_26061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9294 ( .C ( clk ), .D ( new_AGEMA_signal_26068 ), .Q ( new_AGEMA_signal_26069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9302 ( .C ( clk ), .D ( new_AGEMA_signal_26076 ), .Q ( new_AGEMA_signal_26077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9310 ( .C ( clk ), .D ( new_AGEMA_signal_26084 ), .Q ( new_AGEMA_signal_26085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9318 ( .C ( clk ), .D ( new_AGEMA_signal_26092 ), .Q ( new_AGEMA_signal_26093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9326 ( .C ( clk ), .D ( new_AGEMA_signal_26100 ), .Q ( new_AGEMA_signal_26101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9334 ( .C ( clk ), .D ( new_AGEMA_signal_26108 ), .Q ( new_AGEMA_signal_26109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9342 ( .C ( clk ), .D ( new_AGEMA_signal_26116 ), .Q ( new_AGEMA_signal_26117 ) ) ;

    /* cells in depth 31 */
    buf_clk new_AGEMA_reg_buffer_9049 ( .C ( clk ), .D ( new_AGEMA_signal_25823 ), .Q ( new_AGEMA_signal_25824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9063 ( .C ( clk ), .D ( new_AGEMA_signal_25837 ), .Q ( new_AGEMA_signal_25838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9077 ( .C ( clk ), .D ( new_AGEMA_signal_25851 ), .Q ( new_AGEMA_signal_25852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9091 ( .C ( clk ), .D ( new_AGEMA_signal_25865 ), .Q ( new_AGEMA_signal_25866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9105 ( .C ( clk ), .D ( new_AGEMA_signal_25879 ), .Q ( new_AGEMA_signal_25880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9109 ( .C ( clk ), .D ( new_AGEMA_signal_25883 ), .Q ( new_AGEMA_signal_25884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9115 ( .C ( clk ), .D ( new_AGEMA_signal_25889 ), .Q ( new_AGEMA_signal_25890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9121 ( .C ( clk ), .D ( new_AGEMA_signal_25895 ), .Q ( new_AGEMA_signal_25896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9127 ( .C ( clk ), .D ( new_AGEMA_signal_25901 ), .Q ( new_AGEMA_signal_25902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9133 ( .C ( clk ), .D ( new_AGEMA_signal_25907 ), .Q ( new_AGEMA_signal_25908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9139 ( .C ( clk ), .D ( new_AGEMA_signal_25913 ), .Q ( new_AGEMA_signal_25914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9145 ( .C ( clk ), .D ( new_AGEMA_signal_25919 ), .Q ( new_AGEMA_signal_25920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9151 ( .C ( clk ), .D ( new_AGEMA_signal_25925 ), .Q ( new_AGEMA_signal_25926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9157 ( .C ( clk ), .D ( new_AGEMA_signal_25931 ), .Q ( new_AGEMA_signal_25932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9163 ( .C ( clk ), .D ( new_AGEMA_signal_25937 ), .Q ( new_AGEMA_signal_25938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9167 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_25942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9171 ( .C ( clk ), .D ( new_AGEMA_signal_4634 ), .Q ( new_AGEMA_signal_25946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9175 ( .C ( clk ), .D ( new_AGEMA_signal_4635 ), .Q ( new_AGEMA_signal_25950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9179 ( .C ( clk ), .D ( new_AGEMA_signal_4636 ), .Q ( new_AGEMA_signal_25954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9183 ( .C ( clk ), .D ( new_AGEMA_signal_4637 ), .Q ( new_AGEMA_signal_25958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9191 ( .C ( clk ), .D ( new_AGEMA_signal_25965 ), .Q ( new_AGEMA_signal_25966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9199 ( .C ( clk ), .D ( new_AGEMA_signal_25973 ), .Q ( new_AGEMA_signal_25974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9207 ( .C ( clk ), .D ( new_AGEMA_signal_25981 ), .Q ( new_AGEMA_signal_25982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9215 ( .C ( clk ), .D ( new_AGEMA_signal_25989 ), .Q ( new_AGEMA_signal_25990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9223 ( .C ( clk ), .D ( new_AGEMA_signal_25997 ), .Q ( new_AGEMA_signal_25998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9231 ( .C ( clk ), .D ( new_AGEMA_signal_26005 ), .Q ( new_AGEMA_signal_26006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9239 ( .C ( clk ), .D ( new_AGEMA_signal_26013 ), .Q ( new_AGEMA_signal_26014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9247 ( .C ( clk ), .D ( new_AGEMA_signal_26021 ), .Q ( new_AGEMA_signal_26022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9255 ( .C ( clk ), .D ( new_AGEMA_signal_26029 ), .Q ( new_AGEMA_signal_26030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9263 ( .C ( clk ), .D ( new_AGEMA_signal_26037 ), .Q ( new_AGEMA_signal_26038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9271 ( .C ( clk ), .D ( new_AGEMA_signal_26045 ), .Q ( new_AGEMA_signal_26046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9279 ( .C ( clk ), .D ( new_AGEMA_signal_26053 ), .Q ( new_AGEMA_signal_26054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9287 ( .C ( clk ), .D ( new_AGEMA_signal_26061 ), .Q ( new_AGEMA_signal_26062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9295 ( .C ( clk ), .D ( new_AGEMA_signal_26069 ), .Q ( new_AGEMA_signal_26070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9303 ( .C ( clk ), .D ( new_AGEMA_signal_26077 ), .Q ( new_AGEMA_signal_26078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9311 ( .C ( clk ), .D ( new_AGEMA_signal_26085 ), .Q ( new_AGEMA_signal_26086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9319 ( .C ( clk ), .D ( new_AGEMA_signal_26093 ), .Q ( new_AGEMA_signal_26094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9327 ( .C ( clk ), .D ( new_AGEMA_signal_26101 ), .Q ( new_AGEMA_signal_26102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9335 ( .C ( clk ), .D ( new_AGEMA_signal_26109 ), .Q ( new_AGEMA_signal_26110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9343 ( .C ( clk ), .D ( new_AGEMA_signal_26117 ), .Q ( new_AGEMA_signal_26118 ) ) ;

    /* cells in depth 32 */
    nor_HPC1 #(.security_order(4), .pipeline(1)) U2542 ( .ina ({new_AGEMA_signal_25811, new_AGEMA_signal_25797, new_AGEMA_signal_25783, new_AGEMA_signal_25769, new_AGEMA_signal_25755}), .inb ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, new_AGEMA_signal_4638, n2381}), .clk ( clk ), .rnd ({Fresh[13004], Fresh[13003], Fresh[13002], Fresh[13001], Fresh[13000], Fresh[12999], Fresh[12998], Fresh[12997], Fresh[12996], Fresh[12995], Fresh[12994], Fresh[12993], Fresh[12992], Fresh[12991], Fresh[12990]}), .outt ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_9050 ( .C ( clk ), .D ( new_AGEMA_signal_25824 ), .Q ( new_AGEMA_signal_25825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9064 ( .C ( clk ), .D ( new_AGEMA_signal_25838 ), .Q ( new_AGEMA_signal_25839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9078 ( .C ( clk ), .D ( new_AGEMA_signal_25852 ), .Q ( new_AGEMA_signal_25853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9092 ( .C ( clk ), .D ( new_AGEMA_signal_25866 ), .Q ( new_AGEMA_signal_25867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9106 ( .C ( clk ), .D ( new_AGEMA_signal_25880 ), .Q ( new_AGEMA_signal_25881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9110 ( .C ( clk ), .D ( new_AGEMA_signal_25884 ), .Q ( new_AGEMA_signal_25885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9116 ( .C ( clk ), .D ( new_AGEMA_signal_25890 ), .Q ( new_AGEMA_signal_25891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9122 ( .C ( clk ), .D ( new_AGEMA_signal_25896 ), .Q ( new_AGEMA_signal_25897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9128 ( .C ( clk ), .D ( new_AGEMA_signal_25902 ), .Q ( new_AGEMA_signal_25903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9134 ( .C ( clk ), .D ( new_AGEMA_signal_25908 ), .Q ( new_AGEMA_signal_25909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9140 ( .C ( clk ), .D ( new_AGEMA_signal_25914 ), .Q ( new_AGEMA_signal_25915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9146 ( .C ( clk ), .D ( new_AGEMA_signal_25920 ), .Q ( new_AGEMA_signal_25921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9152 ( .C ( clk ), .D ( new_AGEMA_signal_25926 ), .Q ( new_AGEMA_signal_25927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9158 ( .C ( clk ), .D ( new_AGEMA_signal_25932 ), .Q ( new_AGEMA_signal_25933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9164 ( .C ( clk ), .D ( new_AGEMA_signal_25938 ), .Q ( new_AGEMA_signal_25939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9168 ( .C ( clk ), .D ( new_AGEMA_signal_25942 ), .Q ( new_AGEMA_signal_25943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9172 ( .C ( clk ), .D ( new_AGEMA_signal_25946 ), .Q ( new_AGEMA_signal_25947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9176 ( .C ( clk ), .D ( new_AGEMA_signal_25950 ), .Q ( new_AGEMA_signal_25951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9180 ( .C ( clk ), .D ( new_AGEMA_signal_25954 ), .Q ( new_AGEMA_signal_25955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9184 ( .C ( clk ), .D ( new_AGEMA_signal_25958 ), .Q ( new_AGEMA_signal_25959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9192 ( .C ( clk ), .D ( new_AGEMA_signal_25966 ), .Q ( new_AGEMA_signal_25967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9200 ( .C ( clk ), .D ( new_AGEMA_signal_25974 ), .Q ( new_AGEMA_signal_25975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9208 ( .C ( clk ), .D ( new_AGEMA_signal_25982 ), .Q ( new_AGEMA_signal_25983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9216 ( .C ( clk ), .D ( new_AGEMA_signal_25990 ), .Q ( new_AGEMA_signal_25991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9224 ( .C ( clk ), .D ( new_AGEMA_signal_25998 ), .Q ( new_AGEMA_signal_25999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9232 ( .C ( clk ), .D ( new_AGEMA_signal_26006 ), .Q ( new_AGEMA_signal_26007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9240 ( .C ( clk ), .D ( new_AGEMA_signal_26014 ), .Q ( new_AGEMA_signal_26015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9248 ( .C ( clk ), .D ( new_AGEMA_signal_26022 ), .Q ( new_AGEMA_signal_26023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9256 ( .C ( clk ), .D ( new_AGEMA_signal_26030 ), .Q ( new_AGEMA_signal_26031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9264 ( .C ( clk ), .D ( new_AGEMA_signal_26038 ), .Q ( new_AGEMA_signal_26039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9272 ( .C ( clk ), .D ( new_AGEMA_signal_26046 ), .Q ( new_AGEMA_signal_26047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9280 ( .C ( clk ), .D ( new_AGEMA_signal_26054 ), .Q ( new_AGEMA_signal_26055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9288 ( .C ( clk ), .D ( new_AGEMA_signal_26062 ), .Q ( new_AGEMA_signal_26063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9296 ( .C ( clk ), .D ( new_AGEMA_signal_26070 ), .Q ( new_AGEMA_signal_26071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9304 ( .C ( clk ), .D ( new_AGEMA_signal_26078 ), .Q ( new_AGEMA_signal_26079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9312 ( .C ( clk ), .D ( new_AGEMA_signal_26086 ), .Q ( new_AGEMA_signal_26087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9320 ( .C ( clk ), .D ( new_AGEMA_signal_26094 ), .Q ( new_AGEMA_signal_26095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9328 ( .C ( clk ), .D ( new_AGEMA_signal_26102 ), .Q ( new_AGEMA_signal_26103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9336 ( .C ( clk ), .D ( new_AGEMA_signal_26110 ), .Q ( new_AGEMA_signal_26111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9344 ( .C ( clk ), .D ( new_AGEMA_signal_26118 ), .Q ( new_AGEMA_signal_26119 ) ) ;

    /* cells in depth 33 */
    buf_clk new_AGEMA_reg_buffer_9111 ( .C ( clk ), .D ( new_AGEMA_signal_25885 ), .Q ( new_AGEMA_signal_25886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9117 ( .C ( clk ), .D ( new_AGEMA_signal_25891 ), .Q ( new_AGEMA_signal_25892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9123 ( .C ( clk ), .D ( new_AGEMA_signal_25897 ), .Q ( new_AGEMA_signal_25898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9129 ( .C ( clk ), .D ( new_AGEMA_signal_25903 ), .Q ( new_AGEMA_signal_25904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9135 ( .C ( clk ), .D ( new_AGEMA_signal_25909 ), .Q ( new_AGEMA_signal_25910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9141 ( .C ( clk ), .D ( new_AGEMA_signal_25915 ), .Q ( new_AGEMA_signal_25916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9147 ( .C ( clk ), .D ( new_AGEMA_signal_25921 ), .Q ( new_AGEMA_signal_25922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9153 ( .C ( clk ), .D ( new_AGEMA_signal_25927 ), .Q ( new_AGEMA_signal_25928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9159 ( .C ( clk ), .D ( new_AGEMA_signal_25933 ), .Q ( new_AGEMA_signal_25934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9165 ( .C ( clk ), .D ( new_AGEMA_signal_25939 ), .Q ( new_AGEMA_signal_25940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9169 ( .C ( clk ), .D ( new_AGEMA_signal_25943 ), .Q ( new_AGEMA_signal_25944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9173 ( .C ( clk ), .D ( new_AGEMA_signal_25947 ), .Q ( new_AGEMA_signal_25948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9177 ( .C ( clk ), .D ( new_AGEMA_signal_25951 ), .Q ( new_AGEMA_signal_25952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9181 ( .C ( clk ), .D ( new_AGEMA_signal_25955 ), .Q ( new_AGEMA_signal_25956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9185 ( .C ( clk ), .D ( new_AGEMA_signal_25959 ), .Q ( new_AGEMA_signal_25960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9193 ( .C ( clk ), .D ( new_AGEMA_signal_25967 ), .Q ( new_AGEMA_signal_25968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9201 ( .C ( clk ), .D ( new_AGEMA_signal_25975 ), .Q ( new_AGEMA_signal_25976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9209 ( .C ( clk ), .D ( new_AGEMA_signal_25983 ), .Q ( new_AGEMA_signal_25984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9217 ( .C ( clk ), .D ( new_AGEMA_signal_25991 ), .Q ( new_AGEMA_signal_25992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9225 ( .C ( clk ), .D ( new_AGEMA_signal_25999 ), .Q ( new_AGEMA_signal_26000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9233 ( .C ( clk ), .D ( new_AGEMA_signal_26007 ), .Q ( new_AGEMA_signal_26008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9241 ( .C ( clk ), .D ( new_AGEMA_signal_26015 ), .Q ( new_AGEMA_signal_26016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9249 ( .C ( clk ), .D ( new_AGEMA_signal_26023 ), .Q ( new_AGEMA_signal_26024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9257 ( .C ( clk ), .D ( new_AGEMA_signal_26031 ), .Q ( new_AGEMA_signal_26032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9265 ( .C ( clk ), .D ( new_AGEMA_signal_26039 ), .Q ( new_AGEMA_signal_26040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9273 ( .C ( clk ), .D ( new_AGEMA_signal_26047 ), .Q ( new_AGEMA_signal_26048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9281 ( .C ( clk ), .D ( new_AGEMA_signal_26055 ), .Q ( new_AGEMA_signal_26056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9289 ( .C ( clk ), .D ( new_AGEMA_signal_26063 ), .Q ( new_AGEMA_signal_26064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9297 ( .C ( clk ), .D ( new_AGEMA_signal_26071 ), .Q ( new_AGEMA_signal_26072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9305 ( .C ( clk ), .D ( new_AGEMA_signal_26079 ), .Q ( new_AGEMA_signal_26080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9313 ( .C ( clk ), .D ( new_AGEMA_signal_26087 ), .Q ( new_AGEMA_signal_26088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9321 ( .C ( clk ), .D ( new_AGEMA_signal_26095 ), .Q ( new_AGEMA_signal_26096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9329 ( .C ( clk ), .D ( new_AGEMA_signal_26103 ), .Q ( new_AGEMA_signal_26104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9337 ( .C ( clk ), .D ( new_AGEMA_signal_26111 ), .Q ( new_AGEMA_signal_26112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9345 ( .C ( clk ), .D ( new_AGEMA_signal_26119 ), .Q ( new_AGEMA_signal_26120 ) ) ;

    /* cells in depth 34 */
    nand_HPC1 #(.security_order(4), .pipeline(1)) U2584 ( .ina ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, n2427}), .inb ({new_AGEMA_signal_25881, new_AGEMA_signal_25867, new_AGEMA_signal_25853, new_AGEMA_signal_25839, new_AGEMA_signal_25825}), .clk ( clk ), .rnd ({Fresh[13019], Fresh[13018], Fresh[13017], Fresh[13016], Fresh[13015], Fresh[13014], Fresh[13013], Fresh[13012], Fresh[13011], Fresh[13010], Fresh[13009], Fresh[13008], Fresh[13007], Fresh[13006], Fresh[13005]}), .outt ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, new_AGEMA_signal_4647, new_AGEMA_signal_4646, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_9112 ( .C ( clk ), .D ( new_AGEMA_signal_25886 ), .Q ( new_AGEMA_signal_25887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9118 ( .C ( clk ), .D ( new_AGEMA_signal_25892 ), .Q ( new_AGEMA_signal_25893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9124 ( .C ( clk ), .D ( new_AGEMA_signal_25898 ), .Q ( new_AGEMA_signal_25899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9130 ( .C ( clk ), .D ( new_AGEMA_signal_25904 ), .Q ( new_AGEMA_signal_25905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9136 ( .C ( clk ), .D ( new_AGEMA_signal_25910 ), .Q ( new_AGEMA_signal_25911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9142 ( .C ( clk ), .D ( new_AGEMA_signal_25916 ), .Q ( new_AGEMA_signal_25917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9148 ( .C ( clk ), .D ( new_AGEMA_signal_25922 ), .Q ( new_AGEMA_signal_25923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9154 ( .C ( clk ), .D ( new_AGEMA_signal_25928 ), .Q ( new_AGEMA_signal_25929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9160 ( .C ( clk ), .D ( new_AGEMA_signal_25934 ), .Q ( new_AGEMA_signal_25935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9166 ( .C ( clk ), .D ( new_AGEMA_signal_25940 ), .Q ( new_AGEMA_signal_25941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9170 ( .C ( clk ), .D ( new_AGEMA_signal_25944 ), .Q ( new_AGEMA_signal_25945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9174 ( .C ( clk ), .D ( new_AGEMA_signal_25948 ), .Q ( new_AGEMA_signal_25949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9178 ( .C ( clk ), .D ( new_AGEMA_signal_25952 ), .Q ( new_AGEMA_signal_25953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9182 ( .C ( clk ), .D ( new_AGEMA_signal_25956 ), .Q ( new_AGEMA_signal_25957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9186 ( .C ( clk ), .D ( new_AGEMA_signal_25960 ), .Q ( new_AGEMA_signal_25961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9194 ( .C ( clk ), .D ( new_AGEMA_signal_25968 ), .Q ( new_AGEMA_signal_25969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9202 ( .C ( clk ), .D ( new_AGEMA_signal_25976 ), .Q ( new_AGEMA_signal_25977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9210 ( .C ( clk ), .D ( new_AGEMA_signal_25984 ), .Q ( new_AGEMA_signal_25985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9218 ( .C ( clk ), .D ( new_AGEMA_signal_25992 ), .Q ( new_AGEMA_signal_25993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9226 ( .C ( clk ), .D ( new_AGEMA_signal_26000 ), .Q ( new_AGEMA_signal_26001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9234 ( .C ( clk ), .D ( new_AGEMA_signal_26008 ), .Q ( new_AGEMA_signal_26009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9242 ( .C ( clk ), .D ( new_AGEMA_signal_26016 ), .Q ( new_AGEMA_signal_26017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9250 ( .C ( clk ), .D ( new_AGEMA_signal_26024 ), .Q ( new_AGEMA_signal_26025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9258 ( .C ( clk ), .D ( new_AGEMA_signal_26032 ), .Q ( new_AGEMA_signal_26033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9266 ( .C ( clk ), .D ( new_AGEMA_signal_26040 ), .Q ( new_AGEMA_signal_26041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9274 ( .C ( clk ), .D ( new_AGEMA_signal_26048 ), .Q ( new_AGEMA_signal_26049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9282 ( .C ( clk ), .D ( new_AGEMA_signal_26056 ), .Q ( new_AGEMA_signal_26057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9290 ( .C ( clk ), .D ( new_AGEMA_signal_26064 ), .Q ( new_AGEMA_signal_26065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9298 ( .C ( clk ), .D ( new_AGEMA_signal_26072 ), .Q ( new_AGEMA_signal_26073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9306 ( .C ( clk ), .D ( new_AGEMA_signal_26080 ), .Q ( new_AGEMA_signal_26081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9314 ( .C ( clk ), .D ( new_AGEMA_signal_26088 ), .Q ( new_AGEMA_signal_26089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9322 ( .C ( clk ), .D ( new_AGEMA_signal_26096 ), .Q ( new_AGEMA_signal_26097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9330 ( .C ( clk ), .D ( new_AGEMA_signal_26104 ), .Q ( new_AGEMA_signal_26105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9338 ( .C ( clk ), .D ( new_AGEMA_signal_26112 ), .Q ( new_AGEMA_signal_26113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_9346 ( .C ( clk ), .D ( new_AGEMA_signal_26120 ), .Q ( new_AGEMA_signal_26121 ) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_25911, new_AGEMA_signal_25905, new_AGEMA_signal_25899, new_AGEMA_signal_25893, new_AGEMA_signal_25887}), .Q ({SO_s4[7], SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_25941, new_AGEMA_signal_25935, new_AGEMA_signal_25929, new_AGEMA_signal_25923, new_AGEMA_signal_25917}), .Q ({SO_s4[6], SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_25961, new_AGEMA_signal_25957, new_AGEMA_signal_25953, new_AGEMA_signal_25949, new_AGEMA_signal_25945}), .Q ({SO_s4[5], SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_26001, new_AGEMA_signal_25993, new_AGEMA_signal_25985, new_AGEMA_signal_25977, new_AGEMA_signal_25969}), .Q ({SO_s4[4], SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, new_AGEMA_signal_4647, new_AGEMA_signal_4646, N563}), .Q ({SO_s4[3], SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_26041, new_AGEMA_signal_26033, new_AGEMA_signal_26025, new_AGEMA_signal_26017, new_AGEMA_signal_26009}), .Q ({SO_s4[2], SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_26081, new_AGEMA_signal_26073, new_AGEMA_signal_26065, new_AGEMA_signal_26057, new_AGEMA_signal_26049}), .Q ({SO_s4[1], SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_26121, new_AGEMA_signal_26113, new_AGEMA_signal_26105, new_AGEMA_signal_26097, new_AGEMA_signal_26089}), .Q ({SO_s4[0], SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
