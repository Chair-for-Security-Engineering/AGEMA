/* modified netlist. Source: module AES in file ../CaseStudies/08_AES128_round_based_encryption/FPGA_based/AES_synthesis.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module AES_GHPC_ClockGating_d1 (clk, reset, plaintext_s0, key_s0, key_s1, plaintext_s1, Fresh, done, ciphertext_s0, ciphertext_s1, Synch);
    input clk ;
    input reset ;
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [799:0] Fresh ;
    output done ;
    output [127:0] ciphertext_s0 ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_258 ;
    wire \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_259 ;
    wire \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_260 ;
    wire \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_261 ;
    wire \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_262 ;
    wire \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_263 ;
    wire \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_264 ;
    wire \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_265 ;
    wire \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_266 ;
    wire \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_267 ;
    wire \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_268 ;
    wire \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_269 ;
    wire \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_270 ;
    wire \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_271 ;
    wire \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_272 ;
    wire \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_273 ;
    wire \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_274 ;
    wire \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_275 ;
    wire \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_276 ;
    wire \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_277 ;
    wire \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_278 ;
    wire \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_279 ;
    wire \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_280 ;
    wire \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_281 ;
    wire \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_282 ;
    wire \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_283 ;
    wire \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_284 ;
    wire \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_285 ;
    wire \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_286 ;
    wire \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_287 ;
    wire \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_288 ;
    wire \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_289 ;
    wire \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_290 ;
    wire \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_291 ;
    wire \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_292 ;
    wire \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_293 ;
    wire \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_294 ;
    wire \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_295 ;
    wire \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_296 ;
    wire \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_297 ;
    wire \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_298 ;
    wire \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_299 ;
    wire \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_300 ;
    wire \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_301 ;
    wire \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_302 ;
    wire \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_303 ;
    wire \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_304 ;
    wire \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_305 ;
    wire \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_306 ;
    wire \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_307 ;
    wire \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_308 ;
    wire \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_309 ;
    wire \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_310 ;
    wire \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_311 ;
    wire \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_312 ;
    wire \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_313 ;
    wire \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_314 ;
    wire \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_315 ;
    wire \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_316 ;
    wire \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_317 ;
    wire \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_318 ;
    wire \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_319 ;
    wire \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_320 ;
    wire \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_321 ;
    wire \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_322 ;
    wire \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_323 ;
    wire \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_324 ;
    wire \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_325 ;
    wire \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_326 ;
    wire \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_327 ;
    wire \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_328 ;
    wire \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_329 ;
    wire \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_330 ;
    wire \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_331 ;
    wire \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_332 ;
    wire \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_333 ;
    wire \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_334 ;
    wire \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_335 ;
    wire \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_336 ;
    wire \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_337 ;
    wire \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_338 ;
    wire \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_339 ;
    wire \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_340 ;
    wire \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_341 ;
    wire \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_342 ;
    wire \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_343 ;
    wire \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_344 ;
    wire \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_345 ;
    wire \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_346 ;
    wire \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_347 ;
    wire \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_348 ;
    wire \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_349 ;
    wire \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_350 ;
    wire \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_351 ;
    wire \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_352 ;
    wire \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_353 ;
    wire \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_354 ;
    wire \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_355 ;
    wire \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_356 ;
    wire \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_357 ;
    wire \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_358 ;
    wire \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_359 ;
    wire \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_360 ;
    wire \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_361 ;
    wire \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_362 ;
    wire \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_363 ;
    wire \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_364 ;
    wire \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_365 ;
    wire \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_366 ;
    wire \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_367 ;
    wire \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_368 ;
    wire \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_369 ;
    wire \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_370 ;
    wire \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_371 ;
    wire \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_372 ;
    wire \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_373 ;
    wire \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_374 ;
    wire \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_375 ;
    wire \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_376 ;
    wire \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_377 ;
    wire \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_378 ;
    wire \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_379 ;
    wire \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_380 ;
    wire \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_381 ;
    wire \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_382 ;
    wire \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_383 ;
    wire \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_384 ;
    wire \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_385 ;
    wire \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_386 ;
    wire \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_387 ;
    wire \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_388 ;
    wire \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_389 ;
    wire \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_390 ;
    wire \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_391 ;
    wire \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_392 ;
    wire \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_393 ;
    wire \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 ;
    wire \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 ;
    wire \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 ;
    wire \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 ;
    wire \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 ;
    wire \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 ;
    wire \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 ;
    wire \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 ;
    wire \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 ;
    wire \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 ;
    wire \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 ;
    wire \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 ;
    wire \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 ;
    wire \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 ;
    wire \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 ;
    wire \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 ;
    wire \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 ;
    wire \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 ;
    wire \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 ;
    wire \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 ;
    wire \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 ;
    wire \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 ;
    wire \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 ;
    wire \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 ;
    wire \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 ;
    wire \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 ;
    wire \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 ;
    wire \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 ;
    wire \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 ;
    wire \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_423 ;
    wire \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 ;
    wire \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 ;
    wire \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 ;
    wire \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 ;
    wire \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 ;
    wire \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 ;
    wire \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 ;
    wire \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 ;
    wire \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 ;
    wire \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 ;
    wire \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 ;
    wire \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 ;
    wire \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 ;
    wire \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 ;
    wire \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 ;
    wire \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 ;
    wire \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 ;
    wire \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 ;
    wire \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 ;
    wire \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 ;
    wire \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 ;
    wire \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 ;
    wire \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 ;
    wire \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 ;
    wire \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 ;
    wire \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 ;
    wire \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_450 ;
    wire \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_451 ;
    wire \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_452 ;
    wire \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_453 ;
    wire \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_454 ;
    wire \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_455 ;
    wire \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_456 ;
    wire \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_457 ;
    wire \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_458 ;
    wire \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_459 ;
    wire \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_460 ;
    wire \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_461 ;
    wire \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_462 ;
    wire \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_463 ;
    wire \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_464 ;
    wire \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_465 ;
    wire \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_466 ;
    wire \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_467 ;
    wire \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_468 ;
    wire \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_469 ;
    wire \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_470 ;
    wire \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_471 ;
    wire \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_472 ;
    wire \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_473 ;
    wire \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_474 ;
    wire \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_475 ;
    wire \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_476 ;
    wire \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_477 ;
    wire \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_478 ;
    wire \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_479 ;
    wire \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_480 ;
    wire \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_481 ;
    wire \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 ;
    wire \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 ;
    wire \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 ;
    wire \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 ;
    wire \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 ;
    wire \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 ;
    wire \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 ;
    wire \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 ;
    wire \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 ;
    wire \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 ;
    wire \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 ;
    wire \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 ;
    wire \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 ;
    wire \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 ;
    wire \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 ;
    wire \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 ;
    wire \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 ;
    wire \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 ;
    wire \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 ;
    wire \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 ;
    wire \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 ;
    wire \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 ;
    wire \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 ;
    wire \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 ;
    wire \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 ;
    wire \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 ;
    wire \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 ;
    wire \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 ;
    wire \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 ;
    wire \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 ;
    wire \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 ;
    wire \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 ;
    wire \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><4> ;
    wire \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><3> ;
    wire \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><1> ;
    wire \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><3> ;
    wire \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><4> ;
    wire \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><4> ;
    wire \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><1> ;
    wire \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><3> ;
    wire \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><4> ;
    wire \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><1> ;
    wire \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><3> ;
    wire \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><1> ;
    wire LastRound ;
    wire \KeyExpansionOutput<24>_bdd4 ;
    wire \KeyExpansionOutput<31>_bdd4 ;
    wire \KeyExpansionOutput<27>_bdd4 ;
    wire \KeyExpansionOutput<30>_bdd4 ;
    wire \KeyExpansionOutput<28>_bdd4 ;
    wire \KeyExpansionOutput<29>_bdd4 ;
    wire \KeyExpansionOutput<25>_bdd4 ;
    wire \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state ;
    wire \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state ;
    wire \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<0> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<3> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<2> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<1> ;
    wire \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<3> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<0> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<1> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<2> ;
    wire \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<3> ;
    wire N01 ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N10 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N30 ;
    wire N32 ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N50 ;
    wire N52 ;
    wire N54 ;
    wire N56 ;
    wire N58 ;
    wire N60 ;
    wire N62 ;
    wire N64 ;
    wire N66 ;
    wire N68 ;
    wire N70 ;
    wire N72 ;
    wire N74 ;
    wire N76 ;
    wire N78 ;
    wire N80 ;
    wire N82 ;
    wire N84 ;
    wire N86 ;
    wire N88 ;
    wire N90 ;
    wire N92 ;
    wire N94 ;
    wire N96 ;
    wire N98 ;
    wire N100 ;
    wire N102 ;
    wire N104 ;
    wire N106 ;
    wire N108 ;
    wire N110 ;
    wire N112 ;
    wire N114 ;
    wire N116 ;
    wire N118 ;
    wire N120 ;
    wire N122 ;
    wire N124 ;
    wire N126 ;
    wire N128 ;
    wire N130 ;
    wire N132 ;
    wire N134 ;
    wire N136 ;
    wire N138 ;
    wire N140 ;
    wire N142 ;
    wire N144 ;
    wire N146 ;
    wire N148 ;
    wire N150 ;
    wire N152 ;
    wire N154 ;
    wire N156 ;
    wire N158 ;
    wire N160 ;
    wire N162 ;
    wire N164 ;
    wire N166 ;
    wire N168 ;
    wire N170 ;
    wire N172 ;
    wire N174 ;
    wire N176 ;
    wire N178 ;
    wire N180 ;
    wire N182 ;
    wire N184 ;
    wire N186 ;
    wire N188 ;
    wire N190 ;
    wire N192 ;
    wire N194 ;
    wire N196 ;
    wire N198 ;
    wire N200 ;
    wire N202 ;
    wire N204 ;
    wire N206 ;
    wire N208 ;
    wire N210 ;
    wire N212 ;
    wire N214 ;
    wire N216 ;
    wire N218 ;
    wire N220 ;
    wire N222 ;
    wire N224 ;
    wire N226 ;
    wire N228 ;
    wire N230 ;
    wire N232 ;
    wire N234 ;
    wire N236 ;
    wire N238 ;
    wire N240 ;
    wire N242 ;
    wire N244 ;
    wire N246 ;
    wire N248 ;
    wire N250 ;
    wire N252 ;
    wire N254 ;
    wire N256 ;
    wire N258 ;
    wire N260 ;
    wire N262 ;
    wire N264 ;
    wire N266 ;
    wire N268 ;
    wire N270 ;
    wire N272 ;
    wire N274 ;
    wire N276 ;
    wire N278 ;
    wire N280 ;
    wire N282 ;
    wire N284 ;
    wire N286 ;
    wire N288 ;
    wire N290 ;
    wire N292 ;
    wire N294 ;
    wire N296 ;
    wire N298 ;
    wire N300 ;
    wire N302 ;
    wire N304 ;
    wire N306 ;
    wire N308 ;
    wire N310 ;
    wire N312 ;
    wire N314 ;
    wire N316 ;
    wire N318 ;
    wire N320 ;
    wire \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_1_2276 ;
    wire \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_1_2277 ;
    wire \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_1_2278 ;
    wire \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_1_2279 ;
    wire \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_1_2280 ;
    wire \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_1_2281 ;
    wire \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_1_2282 ;
    wire \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_1_2283 ;
    wire \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_1_2284 ;
    wire \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_1_2285 ;
    wire \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_1_2286 ;
    wire \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_1_2287 ;
    wire \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_1_2288 ;
    wire \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_1_2289 ;
    wire \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_1_2290 ;
    wire \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_1_2291 ;
    wire \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_1_2292 ;
    wire \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_1_2293 ;
    wire \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_1_2294 ;
    wire \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_1_2295 ;
    wire \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_1_2296 ;
    wire \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_1_2297 ;
    wire \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_1_2298 ;
    wire \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_1_2299 ;
    wire [3:0] \RoundCounterIns/count ;
    wire [90:90] KeyExpansionOutput ;
    wire [127:0] ShiftRowsInput ;
    wire [23:0] \KeyExpansionIns/tmp ;
    wire [7:0] \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> ;
    wire [3:0] Result ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4197 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT2 #( .INIT ( 4'h6 ) ) \RoundCounterIns/Mcount_count_xor<1>11 ( .I0 (\RoundCounterIns/count [1]), .I1 (\RoundCounterIns/count [0]), .O (Result[1]) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_127_xo<0>1 ( .I0 ({new_AGEMA_signal_2458, \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_258 }), .I1 ({new_AGEMA_signal_2459, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_386 }), .O ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_126_xo<0>1 ( .I0 ({new_AGEMA_signal_2461, \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_259 }), .I1 ({new_AGEMA_signal_2462, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_387 }), .O ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_125_xo<0>1 ( .I0 ({new_AGEMA_signal_2464, \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_260 }), .I1 ({new_AGEMA_signal_2465, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_388 }), .O ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_124_xo<0>1 ( .I0 ({new_AGEMA_signal_2467, \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_261 }), .I1 ({new_AGEMA_signal_2468, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_389 }), .O ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_123_xo<0>1 ( .I0 ({new_AGEMA_signal_2470, \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_262 }), .I1 ({new_AGEMA_signal_2471, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_390 }), .O ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_122_xo<0>1 ( .I0 ({new_AGEMA_signal_2473, \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_263 }), .I1 ({new_AGEMA_signal_2474, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_391 }), .O ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_121_xo<0>1 ( .I0 ({new_AGEMA_signal_2476, \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_264 }), .I1 ({new_AGEMA_signal_2477, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_392 }), .O ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_120_xo<0>1 ( .I0 ({new_AGEMA_signal_2479, \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_265 }), .I1 ({new_AGEMA_signal_2480, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_393 }), .O ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_119_xo<0>1 ( .I0 ({new_AGEMA_signal_2482, \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_266 }), .I1 ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }), .O ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_118_xo<0>1 ( .I0 ({new_AGEMA_signal_2485, \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_267 }), .I1 ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }), .O ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_117_xo<0>1 ( .I0 ({new_AGEMA_signal_2488, \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_268 }), .I1 ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }), .O ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_116_xo<0>1 ( .I0 ({new_AGEMA_signal_2491, \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_269 }), .I1 ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }), .O ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_115_xo<0>1 ( .I0 ({new_AGEMA_signal_2494, \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_270 }), .I1 ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }), .O ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_114_xo<0>1 ( .I0 ({new_AGEMA_signal_2497, \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_271 }), .I1 ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }), .O ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_113_xo<0>1 ( .I0 ({new_AGEMA_signal_2500, \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_272 }), .I1 ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }), .O ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_112_xo<0>1 ( .I0 ({new_AGEMA_signal_2503, \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_273 }), .I1 ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }), .O ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_111_xo<0>1 ( .I0 ({new_AGEMA_signal_2506, \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_274 }), .I1 ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }), .O ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_110_xo<0>1 ( .I0 ({new_AGEMA_signal_2509, \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_275 }), .I1 ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }), .O ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_109_xo<0>1 ( .I0 ({new_AGEMA_signal_2512, \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_276 }), .I1 ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }), .O ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_108_xo<0>1 ( .I0 ({new_AGEMA_signal_2515, \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_277 }), .I1 ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }), .O ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_107_xo<0>1 ( .I0 ({new_AGEMA_signal_2518, \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_278 }), .I1 ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }), .O ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_106_xo<0>1 ( .I0 ({new_AGEMA_signal_2521, \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_279 }), .I1 ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }), .O ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_105_xo<0>1 ( .I0 ({new_AGEMA_signal_2524, \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_280 }), .I1 ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }), .O ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_104_xo<0>1 ( .I0 ({new_AGEMA_signal_2527, \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_281 }), .I1 ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }), .O ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_103_xo<0>1 ( .I0 ({new_AGEMA_signal_2530, \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_282 }), .I1 ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }), .O ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_102_xo<0>1 ( .I0 ({new_AGEMA_signal_2533, \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_283 }), .I1 ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }), .O ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_101_xo<0>1 ( .I0 ({new_AGEMA_signal_2536, \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_284 }), .I1 ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }), .O ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_100_xo<0>1 ( .I0 ({new_AGEMA_signal_2539, \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_285 }), .I1 ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }), .O ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_99_xo<0>1 ( .I0 ({new_AGEMA_signal_2542, \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_286 }), .I1 ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }), .O ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_98_xo<0>1 ( .I0 ({new_AGEMA_signal_2545, \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_287 }), .I1 ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }), .O ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_97_xo<0>1 ( .I0 ({new_AGEMA_signal_2548, \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_288 }), .I1 ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }), .O ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_96_xo<0>1 ( .I0 ({new_AGEMA_signal_2551, \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_289 }), .I1 ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }), .O ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_95_xo<0>1 ( .I0 ({new_AGEMA_signal_2554, \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_290 }), .I1 ({new_AGEMA_signal_2555, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 }), .O ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_94_xo<0>1 ( .I0 ({new_AGEMA_signal_2557, \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_291 }), .I1 ({new_AGEMA_signal_2558, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 }), .O ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_93_xo<0>1 ( .I0 ({new_AGEMA_signal_2560, \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_292 }), .I1 ({new_AGEMA_signal_2561, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 }), .O ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_92_xo<0>1 ( .I0 ({new_AGEMA_signal_2563, \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_293 }), .I1 ({new_AGEMA_signal_2564, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 }), .O ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_91_xo<0>1 ( .I0 ({new_AGEMA_signal_2566, \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_294 }), .I1 ({new_AGEMA_signal_2567, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 }), .O ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_90_xo<0>1 ( .I0 ({new_AGEMA_signal_2569, \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_295 }), .I1 ({new_AGEMA_signal_2570, \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_423 }), .O ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_89_xo<0>1 ( .I0 ({new_AGEMA_signal_2572, \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_296 }), .I1 ({new_AGEMA_signal_2573, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 }), .O ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_88_xo<0>1 ( .I0 ({new_AGEMA_signal_2575, \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_297 }), .I1 ({new_AGEMA_signal_2576, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 }), .O ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_87_xo<0>1 ( .I0 ({new_AGEMA_signal_2578, \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_298 }), .I1 ({new_AGEMA_signal_2579, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 }), .O ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_86_xo<0>1 ( .I0 ({new_AGEMA_signal_2581, \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_299 }), .I1 ({new_AGEMA_signal_2582, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 }), .O ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_85_xo<0>1 ( .I0 ({new_AGEMA_signal_2584, \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_300 }), .I1 ({new_AGEMA_signal_2585, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 }), .O ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_84_xo<0>1 ( .I0 ({new_AGEMA_signal_2587, \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_301 }), .I1 ({new_AGEMA_signal_2588, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 }), .O ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_83_xo<0>1 ( .I0 ({new_AGEMA_signal_2590, \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_302 }), .I1 ({new_AGEMA_signal_2591, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 }), .O ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_82_xo<0>1 ( .I0 ({new_AGEMA_signal_2593, \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_303 }), .I1 ({new_AGEMA_signal_2594, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 }), .O ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_81_xo<0>1 ( .I0 ({new_AGEMA_signal_2596, \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_304 }), .I1 ({new_AGEMA_signal_2597, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 }), .O ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_80_xo<0>1 ( .I0 ({new_AGEMA_signal_2599, \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_305 }), .I1 ({new_AGEMA_signal_2600, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 }), .O ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_79_xo<0>1 ( .I0 ({new_AGEMA_signal_2602, \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_306 }), .I1 ({new_AGEMA_signal_2603, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 }), .O ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_78_xo<0>1 ( .I0 ({new_AGEMA_signal_2605, \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_307 }), .I1 ({new_AGEMA_signal_2606, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 }), .O ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_77_xo<0>1 ( .I0 ({new_AGEMA_signal_2608, \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_308 }), .I1 ({new_AGEMA_signal_2609, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 }), .O ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_76_xo<0>1 ( .I0 ({new_AGEMA_signal_2611, \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_309 }), .I1 ({new_AGEMA_signal_2612, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 }), .O ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_75_xo<0>1 ( .I0 ({new_AGEMA_signal_2614, \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_310 }), .I1 ({new_AGEMA_signal_2615, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 }), .O ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_74_xo<0>1 ( .I0 ({new_AGEMA_signal_2617, \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_311 }), .I1 ({new_AGEMA_signal_2618, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 }), .O ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_73_xo<0>1 ( .I0 ({new_AGEMA_signal_2620, \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_312 }), .I1 ({new_AGEMA_signal_2621, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 }), .O ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_72_xo<0>1 ( .I0 ({new_AGEMA_signal_2623, \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_313 }), .I1 ({new_AGEMA_signal_2624, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 }), .O ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_71_xo<0>1 ( .I0 ({new_AGEMA_signal_2626, \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_314 }), .I1 ({new_AGEMA_signal_2627, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 }), .O ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_70_xo<0>1 ( .I0 ({new_AGEMA_signal_2629, \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_315 }), .I1 ({new_AGEMA_signal_2630, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 }), .O ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_69_xo<0>1 ( .I0 ({new_AGEMA_signal_2632, \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_316 }), .I1 ({new_AGEMA_signal_2633, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 }), .O ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_68_xo<0>1 ( .I0 ({new_AGEMA_signal_2635, \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_317 }), .I1 ({new_AGEMA_signal_2636, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 }), .O ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_67_xo<0>1 ( .I0 ({new_AGEMA_signal_2638, \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_318 }), .I1 ({new_AGEMA_signal_2639, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 }), .O ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_66_xo<0>1 ( .I0 ({new_AGEMA_signal_2641, \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_319 }), .I1 ({new_AGEMA_signal_2642, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 }), .O ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_65_xo<0>1 ( .I0 ({new_AGEMA_signal_2644, \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_320 }), .I1 ({new_AGEMA_signal_2645, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 }), .O ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_64_xo<0>1 ( .I0 ({new_AGEMA_signal_2647, \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_321 }), .I1 ({new_AGEMA_signal_2648, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 }), .O ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_63_xo<0>1 ( .I0 ({new_AGEMA_signal_2650, \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_322 }), .I1 ({new_AGEMA_signal_2651, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_450 }), .O ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_62_xo<0>1 ( .I0 ({new_AGEMA_signal_2653, \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_323 }), .I1 ({new_AGEMA_signal_2654, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_451 }), .O ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_61_xo<0>1 ( .I0 ({new_AGEMA_signal_2656, \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_324 }), .I1 ({new_AGEMA_signal_2657, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_452 }), .O ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_60_xo<0>1 ( .I0 ({new_AGEMA_signal_2659, \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_325 }), .I1 ({new_AGEMA_signal_2660, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_453 }), .O ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_59_xo<0>1 ( .I0 ({new_AGEMA_signal_2662, \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_326 }), .I1 ({new_AGEMA_signal_2663, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_454 }), .O ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_58_xo<0>1 ( .I0 ({new_AGEMA_signal_2665, \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_327 }), .I1 ({new_AGEMA_signal_2666, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_455 }), .O ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_57_xo<0>1 ( .I0 ({new_AGEMA_signal_2668, \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_328 }), .I1 ({new_AGEMA_signal_2669, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_456 }), .O ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_56_xo<0>1 ( .I0 ({new_AGEMA_signal_2671, \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_329 }), .I1 ({new_AGEMA_signal_2672, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_457 }), .O ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_55_xo<0>1 ( .I0 ({new_AGEMA_signal_2674, \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_330 }), .I1 ({new_AGEMA_signal_2675, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_458 }), .O ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_54_xo<0>1 ( .I0 ({new_AGEMA_signal_2677, \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_331 }), .I1 ({new_AGEMA_signal_2678, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_459 }), .O ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_53_xo<0>1 ( .I0 ({new_AGEMA_signal_2680, \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_332 }), .I1 ({new_AGEMA_signal_2681, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_460 }), .O ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_52_xo<0>1 ( .I0 ({new_AGEMA_signal_2683, \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_333 }), .I1 ({new_AGEMA_signal_2684, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_461 }), .O ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_51_xo<0>1 ( .I0 ({new_AGEMA_signal_2686, \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_334 }), .I1 ({new_AGEMA_signal_2687, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_462 }), .O ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_50_xo<0>1 ( .I0 ({new_AGEMA_signal_2689, \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_335 }), .I1 ({new_AGEMA_signal_2690, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_463 }), .O ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_49_xo<0>1 ( .I0 ({new_AGEMA_signal_2692, \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_336 }), .I1 ({new_AGEMA_signal_2693, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_464 }), .O ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_48_xo<0>1 ( .I0 ({new_AGEMA_signal_2695, \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_337 }), .I1 ({new_AGEMA_signal_2696, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_465 }), .O ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_47_xo<0>1 ( .I0 ({new_AGEMA_signal_2698, \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_338 }), .I1 ({new_AGEMA_signal_2699, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_466 }), .O ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_46_xo<0>1 ( .I0 ({new_AGEMA_signal_2701, \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_339 }), .I1 ({new_AGEMA_signal_2702, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_467 }), .O ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_45_xo<0>1 ( .I0 ({new_AGEMA_signal_2704, \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_340 }), .I1 ({new_AGEMA_signal_2705, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_468 }), .O ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_44_xo<0>1 ( .I0 ({new_AGEMA_signal_2707, \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_341 }), .I1 ({new_AGEMA_signal_2708, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_469 }), .O ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_43_xo<0>1 ( .I0 ({new_AGEMA_signal_2710, \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_342 }), .I1 ({new_AGEMA_signal_2711, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_470 }), .O ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_42_xo<0>1 ( .I0 ({new_AGEMA_signal_2713, \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_343 }), .I1 ({new_AGEMA_signal_2714, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_471 }), .O ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_41_xo<0>1 ( .I0 ({new_AGEMA_signal_2716, \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_344 }), .I1 ({new_AGEMA_signal_2717, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_472 }), .O ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_40_xo<0>1 ( .I0 ({new_AGEMA_signal_2719, \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_345 }), .I1 ({new_AGEMA_signal_2720, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_473 }), .O ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_39_xo<0>1 ( .I0 ({new_AGEMA_signal_2722, \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_346 }), .I1 ({new_AGEMA_signal_2723, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_474 }), .O ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_38_xo<0>1 ( .I0 ({new_AGEMA_signal_2725, \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_347 }), .I1 ({new_AGEMA_signal_2726, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_475 }), .O ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_37_xo<0>1 ( .I0 ({new_AGEMA_signal_2728, \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_348 }), .I1 ({new_AGEMA_signal_2729, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_476 }), .O ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_36_xo<0>1 ( .I0 ({new_AGEMA_signal_2731, \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_349 }), .I1 ({new_AGEMA_signal_2732, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_477 }), .O ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_35_xo<0>1 ( .I0 ({new_AGEMA_signal_2734, \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_350 }), .I1 ({new_AGEMA_signal_2735, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_478 }), .O ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_34_xo<0>1 ( .I0 ({new_AGEMA_signal_2737, \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_351 }), .I1 ({new_AGEMA_signal_2738, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_479 }), .O ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_33_xo<0>1 ( .I0 ({new_AGEMA_signal_2740, \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_352 }), .I1 ({new_AGEMA_signal_2741, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_480 }), .O ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_32_xo<0>1 ( .I0 ({new_AGEMA_signal_2743, \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_353 }), .I1 ({new_AGEMA_signal_2744, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_481 }), .O ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_31_xo<0>1 ( .I0 ({new_AGEMA_signal_2746, \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_354 }), .I1 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .O ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_30_xo<0>1 ( .I0 ({new_AGEMA_signal_2749, \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_355 }), .I1 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .O ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_29_xo<0>1 ( .I0 ({new_AGEMA_signal_2752, \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_356 }), .I1 ({new_AGEMA_signal_2753, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_1_2286 }), .O ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_28_xo<0>1 ( .I0 ({new_AGEMA_signal_2755, \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_357 }), .I1 ({new_AGEMA_signal_2756, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_1_2285 }), .O ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_27_xo<0>1 ( .I0 ({new_AGEMA_signal_2758, \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_358 }), .I1 ({new_AGEMA_signal_2759, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_1_2284 }), .O ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_26_xo<0>1 ( .I0 ({new_AGEMA_signal_2761, \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_359 }), .I1 ({new_AGEMA_signal_2762, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_1_2299 }), .O ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_25_xo<0>1 ( .I0 ({new_AGEMA_signal_2764, \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_360 }), .I1 ({new_AGEMA_signal_2765, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_1_2283 }), .O ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_24_xo<0>1 ( .I0 ({new_AGEMA_signal_2767, \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_361 }), .I1 ({new_AGEMA_signal_2768, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_1_2282 }), .O ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_23_xo<0>1 ( .I0 ({new_AGEMA_signal_2770, \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_362 }), .I1 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .O ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_22_xo<0>1 ( .I0 ({new_AGEMA_signal_2773, \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_363 }), .I1 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .O ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_21_xo<0>1 ( .I0 ({new_AGEMA_signal_2776, \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_364 }), .I1 ({new_AGEMA_signal_2777, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_1_2281 }), .O ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_20_xo<0>1 ( .I0 ({new_AGEMA_signal_2779, \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_365 }), .I1 ({new_AGEMA_signal_2780, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_1_2280 }), .O ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_19_xo<0>1 ( .I0 ({new_AGEMA_signal_2782, \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_366 }), .I1 ({new_AGEMA_signal_2783, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_1_2279 }), .O ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_18_xo<0>1 ( .I0 ({new_AGEMA_signal_2785, \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_367 }), .I1 ({new_AGEMA_signal_2786, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_1_2278 }), .O ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_17_xo<0>1 ( .I0 ({new_AGEMA_signal_2788, \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_368 }), .I1 ({new_AGEMA_signal_2789, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_1_2277 }), .O ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_16_xo<0>1 ( .I0 ({new_AGEMA_signal_2791, \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_369 }), .I1 ({new_AGEMA_signal_2792, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_1_2276 }), .O ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_15_xo<0>1 ( .I0 ({new_AGEMA_signal_2794, \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_370 }), .I1 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .O ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_14_xo<0>1 ( .I0 ({new_AGEMA_signal_2797, \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_371 }), .I1 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .O ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_13_xo<0>1 ( .I0 ({new_AGEMA_signal_2800, \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_372 }), .I1 ({new_AGEMA_signal_2801, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_1_2298 }), .O ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_12_xo<0>1 ( .I0 ({new_AGEMA_signal_2803, \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_373 }), .I1 ({new_AGEMA_signal_2804, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_1_2297 }), .O ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_11_xo<0>1 ( .I0 ({new_AGEMA_signal_2806, \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_374 }), .I1 ({new_AGEMA_signal_2807, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_1_2296 }), .O ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_10_xo<0>1 ( .I0 ({new_AGEMA_signal_2809, \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_375 }), .I1 ({new_AGEMA_signal_2810, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_1_2295 }), .O ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_9_xo<0>1 ( .I0 ({new_AGEMA_signal_2812, \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_376 }), .I1 ({new_AGEMA_signal_2813, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_1_2294 }), .O ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_8_xo<0>1 ( .I0 ({new_AGEMA_signal_2815, \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_377 }), .I1 ({new_AGEMA_signal_2816, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_1_2293 }), .O ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_7_xo<0>1 ( .I0 ({new_AGEMA_signal_2818, \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_378 }), .I1 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .O ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_6_xo<0>1 ( .I0 ({new_AGEMA_signal_2821, \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_379 }), .I1 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .O ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_5_xo<0>1 ( .I0 ({new_AGEMA_signal_2824, \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_380 }), .I1 ({new_AGEMA_signal_2825, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_1_2292 }), .O ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_4_xo<0>1 ( .I0 ({new_AGEMA_signal_2827, \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_381 }), .I1 ({new_AGEMA_signal_2828, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_1_2291 }), .O ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_3_xo<0>1 ( .I0 ({new_AGEMA_signal_2830, \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_382 }), .I1 ({new_AGEMA_signal_2831, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_1_2290 }), .O ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_2_xo<0>1 ( .I0 ({new_AGEMA_signal_2833, \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_383 }), .I1 ({new_AGEMA_signal_2834, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_1_2289 }), .O ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_1_xo<0>1 ( .I0 ({new_AGEMA_signal_2836, \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_384 }), .I1 ({new_AGEMA_signal_2837, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_1_2288 }), .O ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \Mxor_ciphertext_0_xo<0>1 ( .I0 ({new_AGEMA_signal_2839, \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_385 }), .I1 ({new_AGEMA_signal_2840, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_1_2287 }), .O ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    LUT4 #( .INIT ( 16'h0200 ) ) \done<3>1 ( .I0 (\RoundCounterIns/count [3]), .I1 (\RoundCounterIns/count [0]), .I2 (\RoundCounterIns/count [2]), .I3 (\RoundCounterIns/count [1]), .O (done) ) ;
    LUT4 #( .INIT ( 16'h6CCC ) ) \Result<3>1 ( .I0 (\RoundCounterIns/count [2]), .I1 (\RoundCounterIns/count [3]), .I2 (\RoundCounterIns/count [0]), .I3 (\RoundCounterIns/count [1]), .O (Result[3]) ) ;
    LUT3 #( .INIT ( 8'h6A ) ) \Result<2>1 ( .I0 (\RoundCounterIns/count [2]), .I1 (\RoundCounterIns/count [0]), .I2 (\RoundCounterIns/count [1]), .O (Result[2]) ) ;
    LUT4 #( .INIT ( 16'h0200 ) ) \LastRound<3>1 ( .I0 (\RoundCounterIns/count [0]), .I1 (\RoundCounterIns/count [2]), .I2 (\RoundCounterIns/count [1]), .I3 (\RoundCounterIns/count [3]), .O (LastRound) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2744, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_481 }), .I1 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .O ({new_AGEMA_signal_2842, N01}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2741, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_480 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .O ({new_AGEMA_signal_2843, N2}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2738, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_479 }), .I1 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .O ({new_AGEMA_signal_2844, N4}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I1 ({new_AGEMA_signal_2735, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_478 }), .O ({new_AGEMA_signal_2845, N6}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2732, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_477 }), .I1 ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }), .O ({new_AGEMA_signal_2846, N8}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2729, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_476 }), .I1 ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }), .O ({new_AGEMA_signal_2847, N10}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2726, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_475 }), .I1 ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }), .O ({new_AGEMA_signal_2848, N12}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2723, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_474 }), .I1 ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }), .O ({new_AGEMA_signal_2849, N14}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2720, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_473 }), .I1 ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }), .O ({new_AGEMA_signal_2850, N16}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2717, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_472 }), .I1 ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }), .O ({new_AGEMA_signal_2851, N18}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I1 ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }), .O ({new_AGEMA_signal_2852, N20}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I1 ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }), .O ({new_AGEMA_signal_2853, N22}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I1 ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }), .O ({new_AGEMA_signal_2854, N24}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .I1 ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }), .O ({new_AGEMA_signal_2855, N26}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I1 ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }), .O ({new_AGEMA_signal_2856, N28}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .I1 ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }), .O ({new_AGEMA_signal_2857, N30}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }), .O ({new_AGEMA_signal_2858, N32}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I1 ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }), .O ({new_AGEMA_signal_2859, N34}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I1 ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }), .O ({new_AGEMA_signal_2860, N36}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I1 ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }), .O ({new_AGEMA_signal_2861, N38}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I1 ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }), .O ({new_AGEMA_signal_2862, N40}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .I1 ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }), .O ({new_AGEMA_signal_2863, N42}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I1 ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }), .O ({new_AGEMA_signal_2864, N44}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .I1 ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }), .O ({new_AGEMA_signal_2865, N46}) ) ;
    LUT2 #( .INIT ( 4'h1 ) ) \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [0]), .I1 (\RoundCounterIns/count [2]), .O (N48) ) ;
    LUT3 #( .INIT ( 8'h54 ) ) \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [2]), .I1 (\RoundCounterIns/count [3]), .I2 (\RoundCounterIns/count [0]), .O (N50) ) ;
    LUT3 #( .INIT ( 8'h42 ) ) \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [3]), .I1 (\RoundCounterIns/count [1]), .I2 (\RoundCounterIns/count [0]), .O (N52) ) ;
    LUT3 #( .INIT ( 8'h26 ) ) \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [3]), .I1 (\RoundCounterIns/count [2]), .I2 (\RoundCounterIns/count [0]), .O (N54) ) ;
    LUT3 #( .INIT ( 8'h28 ) ) \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [0]), .I1 (\RoundCounterIns/count [3]), .I2 (\RoundCounterIns/count [2]), .O (N56) ) ;
    LUT3 #( .INIT ( 8'h20 ) ) \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [1]), .I1 (\RoundCounterIns/count [0]), .I2 (\RoundCounterIns/count [2]), .O (N58) ) ;
    LUT3 #( .INIT ( 8'h80 ) ) \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 (\RoundCounterIns/count [1]), .I1 (\RoundCounterIns/count [0]), .I2 (\RoundCounterIns/count [2]), .O (N60) ) ;
    LUT3 #( .INIT ( 8'hE7 ) ) \KeyExpansionIns/Mxor_OutWords<0>_26_xo<0>1_SW0 ( .I0 (\RoundCounterIns/count [0]), .I1 (\RoundCounterIns/count [3]), .I2 (\RoundCounterIns/count [1]), .O (N318) ) ;
    LUT3 #( .INIT ( 8'h42 ) ) \KeyExpansionIns/Mxor_OutWords<0>_26_xo<0>1_SW1 ( .I0 (\RoundCounterIns/count [1]), .I1 (\RoundCounterIns/count [3]), .I2 (\RoundCounterIns/count [0]), .O (N320) ) ;
    INV \RoundCounterIns/Mcount_count_xor<0>11_INV_0 ( .I (\RoundCounterIns/count [0]), .O (Result[0]) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[0]), .O ({new_AGEMA_signal_2312, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[1]), .O ({new_AGEMA_signal_2313, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[2]), .O ({new_AGEMA_signal_2314, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[3]), .O ({new_AGEMA_signal_2315, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[4]), .O ({new_AGEMA_signal_2316, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[5]), .O ({new_AGEMA_signal_2317, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[6]), .O ({new_AGEMA_signal_2318, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[7]), .O ({new_AGEMA_signal_2319, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[8]), .O ({new_AGEMA_signal_2320, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[9]), .O ({new_AGEMA_signal_2321, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[10]), .O ({new_AGEMA_signal_2322, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[11]), .O ({new_AGEMA_signal_2323, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[12]), .O ({new_AGEMA_signal_2324, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[13]), .O ({new_AGEMA_signal_2325, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[14]), .O ({new_AGEMA_signal_2326, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[15]), .O ({new_AGEMA_signal_2327, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[16]), .O ({new_AGEMA_signal_2328, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[17]), .O ({new_AGEMA_signal_2329, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[18]), .O ({new_AGEMA_signal_2330, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[19]), .O ({new_AGEMA_signal_2331, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[20]), .O ({new_AGEMA_signal_2332, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[21]), .O ({new_AGEMA_signal_2333, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[22]), .O ({new_AGEMA_signal_2334, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[23]), .O ({new_AGEMA_signal_2335, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[24]), .O ({new_AGEMA_signal_2336, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[25]), .O ({new_AGEMA_signal_2337, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[26]), .O ({new_AGEMA_signal_2338, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[27]), .O ({new_AGEMA_signal_2339, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0_3 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[28]), .O ({new_AGEMA_signal_2340, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0_2 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[29]), .O ({new_AGEMA_signal_2341, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0_1 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[30]), .O ({new_AGEMA_signal_2342, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0_0 ( .I0 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I1 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I2 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I3 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I4 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I5 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .clk (clk), .r (Fresh[31]), .O ({new_AGEMA_signal_2343, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[32]), .O ({new_AGEMA_signal_2350, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[33]), .O ({new_AGEMA_signal_2351, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[34]), .O ({new_AGEMA_signal_2352, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[35]), .O ({new_AGEMA_signal_2353, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[36]), .O ({new_AGEMA_signal_2354, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[37]), .O ({new_AGEMA_signal_2355, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[38]), .O ({new_AGEMA_signal_2356, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[39]), .O ({new_AGEMA_signal_2357, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[40]), .O ({new_AGEMA_signal_2358, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[41]), .O ({new_AGEMA_signal_2359, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[42]), .O ({new_AGEMA_signal_2360, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[43]), .O ({new_AGEMA_signal_2361, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[44]), .O ({new_AGEMA_signal_2362, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[45]), .O ({new_AGEMA_signal_2363, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[46]), .O ({new_AGEMA_signal_2364, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[47]), .O ({new_AGEMA_signal_2365, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[48]), .O ({new_AGEMA_signal_2366, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[49]), .O ({new_AGEMA_signal_2367, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[50]), .O ({new_AGEMA_signal_2368, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[51]), .O ({new_AGEMA_signal_2369, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[52]), .O ({new_AGEMA_signal_2370, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[53]), .O ({new_AGEMA_signal_2371, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[54]), .O ({new_AGEMA_signal_2372, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[55]), .O ({new_AGEMA_signal_2373, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[56]), .O ({new_AGEMA_signal_2374, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[57]), .O ({new_AGEMA_signal_2375, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[58]), .O ({new_AGEMA_signal_2376, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[59]), .O ({new_AGEMA_signal_2377, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0_3 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[60]), .O ({new_AGEMA_signal_2378, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0_2 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[61]), .O ({new_AGEMA_signal_2379, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0_1 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[62]), .O ({new_AGEMA_signal_2380, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0_0 ( .I0 ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }), .I1 ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }), .I2 ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }), .I3 ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }), .I4 ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }), .I5 ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }), .clk (clk), .r (Fresh[63]), .O ({new_AGEMA_signal_2381, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[64]), .O ({new_AGEMA_signal_2388, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[65]), .O ({new_AGEMA_signal_2389, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[66]), .O ({new_AGEMA_signal_2390, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[67]), .O ({new_AGEMA_signal_2391, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[68]), .O ({new_AGEMA_signal_2392, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[69]), .O ({new_AGEMA_signal_2393, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[70]), .O ({new_AGEMA_signal_2394, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[71]), .O ({new_AGEMA_signal_2395, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[72]), .O ({new_AGEMA_signal_2396, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[73]), .O ({new_AGEMA_signal_2397, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[74]), .O ({new_AGEMA_signal_2398, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[75]), .O ({new_AGEMA_signal_2399, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[76]), .O ({new_AGEMA_signal_2400, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[77]), .O ({new_AGEMA_signal_2401, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[78]), .O ({new_AGEMA_signal_2402, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[79]), .O ({new_AGEMA_signal_2403, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[80]), .O ({new_AGEMA_signal_2404, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[81]), .O ({new_AGEMA_signal_2405, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[82]), .O ({new_AGEMA_signal_2406, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[83]), .O ({new_AGEMA_signal_2407, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[84]), .O ({new_AGEMA_signal_2408, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[85]), .O ({new_AGEMA_signal_2409, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[86]), .O ({new_AGEMA_signal_2410, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[87]), .O ({new_AGEMA_signal_2411, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[88]), .O ({new_AGEMA_signal_2412, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[89]), .O ({new_AGEMA_signal_2413, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[90]), .O ({new_AGEMA_signal_2414, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[91]), .O ({new_AGEMA_signal_2415, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0_3 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[92]), .O ({new_AGEMA_signal_2416, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0_2 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[93]), .O ({new_AGEMA_signal_2417, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0_1 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[94]), .O ({new_AGEMA_signal_2418, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0_0 ( .I0 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I1 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I2 ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }), .I3 ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }), .I4 ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }), .I5 ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }), .clk (clk), .r (Fresh[95]), .O ({new_AGEMA_signal_2419, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[96]), .O ({new_AGEMA_signal_2426, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[97]), .O ({new_AGEMA_signal_2427, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[98]), .O ({new_AGEMA_signal_2428, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[99]), .O ({new_AGEMA_signal_2429, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[100]), .O ({new_AGEMA_signal_2430, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[101]), .O ({new_AGEMA_signal_2431, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[102]), .O ({new_AGEMA_signal_2432, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[103]), .O ({new_AGEMA_signal_2433, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[104]), .O ({new_AGEMA_signal_2434, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[105]), .O ({new_AGEMA_signal_2435, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[106]), .O ({new_AGEMA_signal_2436, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[107]), .O ({new_AGEMA_signal_2437, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[108]), .O ({new_AGEMA_signal_2438, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[109]), .O ({new_AGEMA_signal_2439, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[110]), .O ({new_AGEMA_signal_2440, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[111]), .O ({new_AGEMA_signal_2441, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[112]), .O ({new_AGEMA_signal_2442, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[113]), .O ({new_AGEMA_signal_2443, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[114]), .O ({new_AGEMA_signal_2444, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[115]), .O ({new_AGEMA_signal_2445, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[116]), .O ({new_AGEMA_signal_2446, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[117]), .O ({new_AGEMA_signal_2447, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[118]), .O ({new_AGEMA_signal_2448, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[119]), .O ({new_AGEMA_signal_2449, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[120]), .O ({new_AGEMA_signal_2450, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[121]), .O ({new_AGEMA_signal_2451, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[122]), .O ({new_AGEMA_signal_2452, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[123]), .O ({new_AGEMA_signal_2453, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0_3 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[124]), .O ({new_AGEMA_signal_2454, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0_2 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[125]), .O ({new_AGEMA_signal_2455, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0_1 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[126]), .O ({new_AGEMA_signal_2456, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0_0 ( .I0 ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }), .I1 ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }), .I2 ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }), .I3 ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }), .I4 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I5 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .clk (clk), .r (Fresh[127]), .O ({new_AGEMA_signal_2457, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[128]), .O ({new_AGEMA_signal_2898, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[129]), .O ({new_AGEMA_signal_2899, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[130]), .O ({new_AGEMA_signal_2900, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[131]), .O ({new_AGEMA_signal_2901, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[132]), .O ({new_AGEMA_signal_2902, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[133]), .O ({new_AGEMA_signal_2903, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[134]), .O ({new_AGEMA_signal_2904, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[135]), .O ({new_AGEMA_signal_2905, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[136]), .O ({new_AGEMA_signal_2906, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[137]), .O ({new_AGEMA_signal_2907, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[138]), .O ({new_AGEMA_signal_2908, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[139]), .O ({new_AGEMA_signal_2909, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[140]), .O ({new_AGEMA_signal_2910, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[141]), .O ({new_AGEMA_signal_2911, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[142]), .O ({new_AGEMA_signal_2912, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[143]), .O ({new_AGEMA_signal_2913, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[144]), .O ({new_AGEMA_signal_2914, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[145]), .O ({new_AGEMA_signal_2915, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[146]), .O ({new_AGEMA_signal_2916, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[147]), .O ({new_AGEMA_signal_2917, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[148]), .O ({new_AGEMA_signal_2918, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[149]), .O ({new_AGEMA_signal_2919, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[150]), .O ({new_AGEMA_signal_2920, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[151]), .O ({new_AGEMA_signal_2921, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[152]), .O ({new_AGEMA_signal_2922, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[153]), .O ({new_AGEMA_signal_2923, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[154]), .O ({new_AGEMA_signal_2924, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[155]), .O ({new_AGEMA_signal_2925, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[156]), .O ({new_AGEMA_signal_2926, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[157]), .O ({new_AGEMA_signal_2927, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[158]), .O ({new_AGEMA_signal_2928, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[0], ciphertext_s0[0]}), .I1 ({ciphertext_s1[1], ciphertext_s0[1]}), .I2 ({ciphertext_s1[2], ciphertext_s0[2]}), .I3 ({ciphertext_s1[3], ciphertext_s0[3]}), .I4 ({ciphertext_s1[4], ciphertext_s0[4]}), .I5 ({ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r (Fresh[159]), .O ({new_AGEMA_signal_2929, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[160]), .O ({new_AGEMA_signal_2930, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[161]), .O ({new_AGEMA_signal_2931, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[162]), .O ({new_AGEMA_signal_2932, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[163]), .O ({new_AGEMA_signal_2933, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[164]), .O ({new_AGEMA_signal_2934, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[165]), .O ({new_AGEMA_signal_2935, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[166]), .O ({new_AGEMA_signal_2936, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[167]), .O ({new_AGEMA_signal_2937, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[168]), .O ({new_AGEMA_signal_2938, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[169]), .O ({new_AGEMA_signal_2939, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[170]), .O ({new_AGEMA_signal_2940, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[171]), .O ({new_AGEMA_signal_2941, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[172]), .O ({new_AGEMA_signal_2942, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[173]), .O ({new_AGEMA_signal_2943, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[174]), .O ({new_AGEMA_signal_2944, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[175]), .O ({new_AGEMA_signal_2945, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[176]), .O ({new_AGEMA_signal_2946, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[177]), .O ({new_AGEMA_signal_2947, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[178]), .O ({new_AGEMA_signal_2948, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[179]), .O ({new_AGEMA_signal_2949, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[180]), .O ({new_AGEMA_signal_2950, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[181]), .O ({new_AGEMA_signal_2951, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[182]), .O ({new_AGEMA_signal_2952, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[183]), .O ({new_AGEMA_signal_2953, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[184]), .O ({new_AGEMA_signal_2954, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[185]), .O ({new_AGEMA_signal_2955, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[186]), .O ({new_AGEMA_signal_2956, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[187]), .O ({new_AGEMA_signal_2957, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[188]), .O ({new_AGEMA_signal_2958, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[189]), .O ({new_AGEMA_signal_2959, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[190]), .O ({new_AGEMA_signal_2960, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[8], ciphertext_s0[8]}), .I1 ({ciphertext_s1[9], ciphertext_s0[9]}), .I2 ({ciphertext_s1[10], ciphertext_s0[10]}), .I3 ({ciphertext_s1[11], ciphertext_s0[11]}), .I4 ({ciphertext_s1[12], ciphertext_s0[12]}), .I5 ({ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r (Fresh[191]), .O ({new_AGEMA_signal_2961, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[192]), .O ({new_AGEMA_signal_2962, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[193]), .O ({new_AGEMA_signal_2963, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[194]), .O ({new_AGEMA_signal_2964, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[195]), .O ({new_AGEMA_signal_2965, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[196]), .O ({new_AGEMA_signal_2966, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[197]), .O ({new_AGEMA_signal_2967, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[198]), .O ({new_AGEMA_signal_2968, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[199]), .O ({new_AGEMA_signal_2969, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[200]), .O ({new_AGEMA_signal_2970, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[201]), .O ({new_AGEMA_signal_2971, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[202]), .O ({new_AGEMA_signal_2972, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[203]), .O ({new_AGEMA_signal_2973, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[204]), .O ({new_AGEMA_signal_2974, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[205]), .O ({new_AGEMA_signal_2975, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[206]), .O ({new_AGEMA_signal_2976, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[207]), .O ({new_AGEMA_signal_2977, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[208]), .O ({new_AGEMA_signal_2978, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[209]), .O ({new_AGEMA_signal_2979, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[210]), .O ({new_AGEMA_signal_2980, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[211]), .O ({new_AGEMA_signal_2981, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[212]), .O ({new_AGEMA_signal_2982, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[213]), .O ({new_AGEMA_signal_2983, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[214]), .O ({new_AGEMA_signal_2984, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[215]), .O ({new_AGEMA_signal_2985, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[216]), .O ({new_AGEMA_signal_2986, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[217]), .O ({new_AGEMA_signal_2987, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[218]), .O ({new_AGEMA_signal_2988, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[219]), .O ({new_AGEMA_signal_2989, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[220]), .O ({new_AGEMA_signal_2990, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[221]), .O ({new_AGEMA_signal_2991, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[222]), .O ({new_AGEMA_signal_2992, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[16], ciphertext_s0[16]}), .I1 ({ciphertext_s1[17], ciphertext_s0[17]}), .I2 ({ciphertext_s1[18], ciphertext_s0[18]}), .I3 ({ciphertext_s1[19], ciphertext_s0[19]}), .I4 ({ciphertext_s1[20], ciphertext_s0[20]}), .I5 ({ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r (Fresh[223]), .O ({new_AGEMA_signal_2993, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[224]), .O ({new_AGEMA_signal_2994, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[225]), .O ({new_AGEMA_signal_2995, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[226]), .O ({new_AGEMA_signal_2996, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[227]), .O ({new_AGEMA_signal_2997, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[228]), .O ({new_AGEMA_signal_2998, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[229]), .O ({new_AGEMA_signal_2999, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[230]), .O ({new_AGEMA_signal_3000, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[231]), .O ({new_AGEMA_signal_3001, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[232]), .O ({new_AGEMA_signal_3002, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[233]), .O ({new_AGEMA_signal_3003, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[234]), .O ({new_AGEMA_signal_3004, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[235]), .O ({new_AGEMA_signal_3005, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[236]), .O ({new_AGEMA_signal_3006, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[237]), .O ({new_AGEMA_signal_3007, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[238]), .O ({new_AGEMA_signal_3008, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[239]), .O ({new_AGEMA_signal_3009, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[240]), .O ({new_AGEMA_signal_3010, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[241]), .O ({new_AGEMA_signal_3011, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[242]), .O ({new_AGEMA_signal_3012, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[243]), .O ({new_AGEMA_signal_3013, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[244]), .O ({new_AGEMA_signal_3014, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[245]), .O ({new_AGEMA_signal_3015, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[246]), .O ({new_AGEMA_signal_3016, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[247]), .O ({new_AGEMA_signal_3017, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[248]), .O ({new_AGEMA_signal_3018, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[249]), .O ({new_AGEMA_signal_3019, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[250]), .O ({new_AGEMA_signal_3020, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[251]), .O ({new_AGEMA_signal_3021, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[252]), .O ({new_AGEMA_signal_3022, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[253]), .O ({new_AGEMA_signal_3023, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[254]), .O ({new_AGEMA_signal_3024, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[24], ciphertext_s0[24]}), .I1 ({ciphertext_s1[25], ciphertext_s0[25]}), .I2 ({ciphertext_s1[26], ciphertext_s0[26]}), .I3 ({ciphertext_s1[27], ciphertext_s0[27]}), .I4 ({ciphertext_s1[28], ciphertext_s0[28]}), .I5 ({ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r (Fresh[255]), .O ({new_AGEMA_signal_3025, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[256]), .O ({new_AGEMA_signal_3026, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[257]), .O ({new_AGEMA_signal_3027, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[258]), .O ({new_AGEMA_signal_3028, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[259]), .O ({new_AGEMA_signal_3029, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[260]), .O ({new_AGEMA_signal_3030, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[261]), .O ({new_AGEMA_signal_3031, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[262]), .O ({new_AGEMA_signal_3032, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[263]), .O ({new_AGEMA_signal_3033, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[264]), .O ({new_AGEMA_signal_3034, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[265]), .O ({new_AGEMA_signal_3035, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[266]), .O ({new_AGEMA_signal_3036, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[267]), .O ({new_AGEMA_signal_3037, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[268]), .O ({new_AGEMA_signal_3038, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[269]), .O ({new_AGEMA_signal_3039, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[270]), .O ({new_AGEMA_signal_3040, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[271]), .O ({new_AGEMA_signal_3041, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[272]), .O ({new_AGEMA_signal_3042, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[273]), .O ({new_AGEMA_signal_3043, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[274]), .O ({new_AGEMA_signal_3044, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[275]), .O ({new_AGEMA_signal_3045, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[276]), .O ({new_AGEMA_signal_3046, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[277]), .O ({new_AGEMA_signal_3047, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[278]), .O ({new_AGEMA_signal_3048, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[279]), .O ({new_AGEMA_signal_3049, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[280]), .O ({new_AGEMA_signal_3050, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[281]), .O ({new_AGEMA_signal_3051, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[282]), .O ({new_AGEMA_signal_3052, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[283]), .O ({new_AGEMA_signal_3053, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[284]), .O ({new_AGEMA_signal_3054, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[285]), .O ({new_AGEMA_signal_3055, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[286]), .O ({new_AGEMA_signal_3056, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[32], ciphertext_s0[32]}), .I1 ({ciphertext_s1[33], ciphertext_s0[33]}), .I2 ({ciphertext_s1[34], ciphertext_s0[34]}), .I3 ({ciphertext_s1[35], ciphertext_s0[35]}), .I4 ({ciphertext_s1[36], ciphertext_s0[36]}), .I5 ({ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r (Fresh[287]), .O ({new_AGEMA_signal_3057, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[288]), .O ({new_AGEMA_signal_3058, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[289]), .O ({new_AGEMA_signal_3059, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[290]), .O ({new_AGEMA_signal_3060, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[291]), .O ({new_AGEMA_signal_3061, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[292]), .O ({new_AGEMA_signal_3062, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[293]), .O ({new_AGEMA_signal_3063, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[294]), .O ({new_AGEMA_signal_3064, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[295]), .O ({new_AGEMA_signal_3065, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[296]), .O ({new_AGEMA_signal_3066, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[297]), .O ({new_AGEMA_signal_3067, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[298]), .O ({new_AGEMA_signal_3068, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[299]), .O ({new_AGEMA_signal_3069, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[300]), .O ({new_AGEMA_signal_3070, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[301]), .O ({new_AGEMA_signal_3071, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[302]), .O ({new_AGEMA_signal_3072, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[303]), .O ({new_AGEMA_signal_3073, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[304]), .O ({new_AGEMA_signal_3074, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[305]), .O ({new_AGEMA_signal_3075, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[306]), .O ({new_AGEMA_signal_3076, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[307]), .O ({new_AGEMA_signal_3077, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[308]), .O ({new_AGEMA_signal_3078, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[309]), .O ({new_AGEMA_signal_3079, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[310]), .O ({new_AGEMA_signal_3080, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[311]), .O ({new_AGEMA_signal_3081, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[312]), .O ({new_AGEMA_signal_3082, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[313]), .O ({new_AGEMA_signal_3083, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[314]), .O ({new_AGEMA_signal_3084, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[315]), .O ({new_AGEMA_signal_3085, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[316]), .O ({new_AGEMA_signal_3086, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[317]), .O ({new_AGEMA_signal_3087, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[318]), .O ({new_AGEMA_signal_3088, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[40], ciphertext_s0[40]}), .I1 ({ciphertext_s1[41], ciphertext_s0[41]}), .I2 ({ciphertext_s1[42], ciphertext_s0[42]}), .I3 ({ciphertext_s1[43], ciphertext_s0[43]}), .I4 ({ciphertext_s1[44], ciphertext_s0[44]}), .I5 ({ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r (Fresh[319]), .O ({new_AGEMA_signal_3089, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[320]), .O ({new_AGEMA_signal_3090, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[321]), .O ({new_AGEMA_signal_3091, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[322]), .O ({new_AGEMA_signal_3092, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[323]), .O ({new_AGEMA_signal_3093, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[324]), .O ({new_AGEMA_signal_3094, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[325]), .O ({new_AGEMA_signal_3095, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[326]), .O ({new_AGEMA_signal_3096, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[327]), .O ({new_AGEMA_signal_3097, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[328]), .O ({new_AGEMA_signal_3098, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[329]), .O ({new_AGEMA_signal_3099, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[330]), .O ({new_AGEMA_signal_3100, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[331]), .O ({new_AGEMA_signal_3101, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[332]), .O ({new_AGEMA_signal_3102, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[333]), .O ({new_AGEMA_signal_3103, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[334]), .O ({new_AGEMA_signal_3104, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[335]), .O ({new_AGEMA_signal_3105, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[336]), .O ({new_AGEMA_signal_3106, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[337]), .O ({new_AGEMA_signal_3107, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[338]), .O ({new_AGEMA_signal_3108, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[339]), .O ({new_AGEMA_signal_3109, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[340]), .O ({new_AGEMA_signal_3110, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[341]), .O ({new_AGEMA_signal_3111, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[342]), .O ({new_AGEMA_signal_3112, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[343]), .O ({new_AGEMA_signal_3113, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[344]), .O ({new_AGEMA_signal_3114, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[345]), .O ({new_AGEMA_signal_3115, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[346]), .O ({new_AGEMA_signal_3116, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[347]), .O ({new_AGEMA_signal_3117, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[348]), .O ({new_AGEMA_signal_3118, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[349]), .O ({new_AGEMA_signal_3119, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[350]), .O ({new_AGEMA_signal_3120, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[48], ciphertext_s0[48]}), .I1 ({ciphertext_s1[49], ciphertext_s0[49]}), .I2 ({ciphertext_s1[50], ciphertext_s0[50]}), .I3 ({ciphertext_s1[51], ciphertext_s0[51]}), .I4 ({ciphertext_s1[52], ciphertext_s0[52]}), .I5 ({ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r (Fresh[351]), .O ({new_AGEMA_signal_3121, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[352]), .O ({new_AGEMA_signal_3122, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[353]), .O ({new_AGEMA_signal_3123, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[354]), .O ({new_AGEMA_signal_3124, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[355]), .O ({new_AGEMA_signal_3125, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[356]), .O ({new_AGEMA_signal_3126, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[357]), .O ({new_AGEMA_signal_3127, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[358]), .O ({new_AGEMA_signal_3128, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[359]), .O ({new_AGEMA_signal_3129, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[360]), .O ({new_AGEMA_signal_3130, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[361]), .O ({new_AGEMA_signal_3131, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[362]), .O ({new_AGEMA_signal_3132, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[363]), .O ({new_AGEMA_signal_3133, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[364]), .O ({new_AGEMA_signal_3134, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[365]), .O ({new_AGEMA_signal_3135, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[366]), .O ({new_AGEMA_signal_3136, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[367]), .O ({new_AGEMA_signal_3137, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[368]), .O ({new_AGEMA_signal_3138, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[369]), .O ({new_AGEMA_signal_3139, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[370]), .O ({new_AGEMA_signal_3140, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[371]), .O ({new_AGEMA_signal_3141, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[372]), .O ({new_AGEMA_signal_3142, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[373]), .O ({new_AGEMA_signal_3143, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[374]), .O ({new_AGEMA_signal_3144, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[375]), .O ({new_AGEMA_signal_3145, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[376]), .O ({new_AGEMA_signal_3146, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[377]), .O ({new_AGEMA_signal_3147, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[378]), .O ({new_AGEMA_signal_3148, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[379]), .O ({new_AGEMA_signal_3149, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[380]), .O ({new_AGEMA_signal_3150, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[381]), .O ({new_AGEMA_signal_3151, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[382]), .O ({new_AGEMA_signal_3152, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[56], ciphertext_s0[56]}), .I1 ({ciphertext_s1[57], ciphertext_s0[57]}), .I2 ({ciphertext_s1[58], ciphertext_s0[58]}), .I3 ({ciphertext_s1[59], ciphertext_s0[59]}), .I4 ({ciphertext_s1[60], ciphertext_s0[60]}), .I5 ({ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r (Fresh[383]), .O ({new_AGEMA_signal_3153, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[384]), .O ({new_AGEMA_signal_3154, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[385]), .O ({new_AGEMA_signal_3155, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[386]), .O ({new_AGEMA_signal_3156, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[387]), .O ({new_AGEMA_signal_3157, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[388]), .O ({new_AGEMA_signal_3158, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[389]), .O ({new_AGEMA_signal_3159, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[390]), .O ({new_AGEMA_signal_3160, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[391]), .O ({new_AGEMA_signal_3161, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[392]), .O ({new_AGEMA_signal_3162, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[393]), .O ({new_AGEMA_signal_3163, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[394]), .O ({new_AGEMA_signal_3164, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[395]), .O ({new_AGEMA_signal_3165, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[396]), .O ({new_AGEMA_signal_3166, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[397]), .O ({new_AGEMA_signal_3167, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[398]), .O ({new_AGEMA_signal_3168, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[399]), .O ({new_AGEMA_signal_3169, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[400]), .O ({new_AGEMA_signal_3170, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[401]), .O ({new_AGEMA_signal_3171, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[402]), .O ({new_AGEMA_signal_3172, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[403]), .O ({new_AGEMA_signal_3173, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[404]), .O ({new_AGEMA_signal_3174, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[405]), .O ({new_AGEMA_signal_3175, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[406]), .O ({new_AGEMA_signal_3176, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[407]), .O ({new_AGEMA_signal_3177, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[408]), .O ({new_AGEMA_signal_3178, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[409]), .O ({new_AGEMA_signal_3179, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[410]), .O ({new_AGEMA_signal_3180, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[411]), .O ({new_AGEMA_signal_3181, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[412]), .O ({new_AGEMA_signal_3182, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[413]), .O ({new_AGEMA_signal_3183, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[414]), .O ({new_AGEMA_signal_3184, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[64], ciphertext_s0[64]}), .I1 ({ciphertext_s1[65], ciphertext_s0[65]}), .I2 ({ciphertext_s1[66], ciphertext_s0[66]}), .I3 ({ciphertext_s1[67], ciphertext_s0[67]}), .I4 ({ciphertext_s1[68], ciphertext_s0[68]}), .I5 ({ciphertext_s1[69], ciphertext_s0[69]}), .clk (clk), .r (Fresh[415]), .O ({new_AGEMA_signal_3185, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[416]), .O ({new_AGEMA_signal_3186, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[417]), .O ({new_AGEMA_signal_3187, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[418]), .O ({new_AGEMA_signal_3188, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[419]), .O ({new_AGEMA_signal_3189, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[420]), .O ({new_AGEMA_signal_3190, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[421]), .O ({new_AGEMA_signal_3191, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[422]), .O ({new_AGEMA_signal_3192, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[423]), .O ({new_AGEMA_signal_3193, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[424]), .O ({new_AGEMA_signal_3194, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[425]), .O ({new_AGEMA_signal_3195, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[426]), .O ({new_AGEMA_signal_3196, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[427]), .O ({new_AGEMA_signal_3197, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[428]), .O ({new_AGEMA_signal_3198, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[429]), .O ({new_AGEMA_signal_3199, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[430]), .O ({new_AGEMA_signal_3200, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[431]), .O ({new_AGEMA_signal_3201, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[432]), .O ({new_AGEMA_signal_3202, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[433]), .O ({new_AGEMA_signal_3203, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[434]), .O ({new_AGEMA_signal_3204, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[435]), .O ({new_AGEMA_signal_3205, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[436]), .O ({new_AGEMA_signal_3206, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[437]), .O ({new_AGEMA_signal_3207, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[438]), .O ({new_AGEMA_signal_3208, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[439]), .O ({new_AGEMA_signal_3209, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[440]), .O ({new_AGEMA_signal_3210, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[441]), .O ({new_AGEMA_signal_3211, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[442]), .O ({new_AGEMA_signal_3212, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[443]), .O ({new_AGEMA_signal_3213, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[444]), .O ({new_AGEMA_signal_3214, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[445]), .O ({new_AGEMA_signal_3215, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[446]), .O ({new_AGEMA_signal_3216, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[72], ciphertext_s0[72]}), .I1 ({ciphertext_s1[73], ciphertext_s0[73]}), .I2 ({ciphertext_s1[74], ciphertext_s0[74]}), .I3 ({ciphertext_s1[75], ciphertext_s0[75]}), .I4 ({ciphertext_s1[76], ciphertext_s0[76]}), .I5 ({ciphertext_s1[77], ciphertext_s0[77]}), .clk (clk), .r (Fresh[447]), .O ({new_AGEMA_signal_3217, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[448]), .O ({new_AGEMA_signal_3218, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[449]), .O ({new_AGEMA_signal_3219, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[450]), .O ({new_AGEMA_signal_3220, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[451]), .O ({new_AGEMA_signal_3221, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[452]), .O ({new_AGEMA_signal_3222, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[453]), .O ({new_AGEMA_signal_3223, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[454]), .O ({new_AGEMA_signal_3224, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[455]), .O ({new_AGEMA_signal_3225, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[456]), .O ({new_AGEMA_signal_3226, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[457]), .O ({new_AGEMA_signal_3227, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[458]), .O ({new_AGEMA_signal_3228, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[459]), .O ({new_AGEMA_signal_3229, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[460]), .O ({new_AGEMA_signal_3230, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[461]), .O ({new_AGEMA_signal_3231, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[462]), .O ({new_AGEMA_signal_3232, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[463]), .O ({new_AGEMA_signal_3233, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[464]), .O ({new_AGEMA_signal_3234, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[465]), .O ({new_AGEMA_signal_3235, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[466]), .O ({new_AGEMA_signal_3236, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[467]), .O ({new_AGEMA_signal_3237, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[468]), .O ({new_AGEMA_signal_3238, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[469]), .O ({new_AGEMA_signal_3239, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[470]), .O ({new_AGEMA_signal_3240, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[471]), .O ({new_AGEMA_signal_3241, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[472]), .O ({new_AGEMA_signal_3242, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[473]), .O ({new_AGEMA_signal_3243, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[474]), .O ({new_AGEMA_signal_3244, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[475]), .O ({new_AGEMA_signal_3245, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[476]), .O ({new_AGEMA_signal_3246, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[477]), .O ({new_AGEMA_signal_3247, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[478]), .O ({new_AGEMA_signal_3248, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[80], ciphertext_s0[80]}), .I1 ({ciphertext_s1[81], ciphertext_s0[81]}), .I2 ({ciphertext_s1[82], ciphertext_s0[82]}), .I3 ({ciphertext_s1[83], ciphertext_s0[83]}), .I4 ({ciphertext_s1[84], ciphertext_s0[84]}), .I5 ({ciphertext_s1[85], ciphertext_s0[85]}), .clk (clk), .r (Fresh[479]), .O ({new_AGEMA_signal_3249, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[480]), .O ({new_AGEMA_signal_3250, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[481]), .O ({new_AGEMA_signal_3251, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[482]), .O ({new_AGEMA_signal_3252, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[483]), .O ({new_AGEMA_signal_3253, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[484]), .O ({new_AGEMA_signal_3254, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[485]), .O ({new_AGEMA_signal_3255, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[486]), .O ({new_AGEMA_signal_3256, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[487]), .O ({new_AGEMA_signal_3257, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[488]), .O ({new_AGEMA_signal_3258, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[489]), .O ({new_AGEMA_signal_3259, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[490]), .O ({new_AGEMA_signal_3260, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[491]), .O ({new_AGEMA_signal_3261, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[492]), .O ({new_AGEMA_signal_3262, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[493]), .O ({new_AGEMA_signal_3263, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[494]), .O ({new_AGEMA_signal_3264, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[495]), .O ({new_AGEMA_signal_3265, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[496]), .O ({new_AGEMA_signal_3266, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[497]), .O ({new_AGEMA_signal_3267, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[498]), .O ({new_AGEMA_signal_3268, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[499]), .O ({new_AGEMA_signal_3269, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[500]), .O ({new_AGEMA_signal_3270, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[501]), .O ({new_AGEMA_signal_3271, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[502]), .O ({new_AGEMA_signal_3272, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[503]), .O ({new_AGEMA_signal_3273, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[504]), .O ({new_AGEMA_signal_3274, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[505]), .O ({new_AGEMA_signal_3275, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[506]), .O ({new_AGEMA_signal_3276, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[507]), .O ({new_AGEMA_signal_3277, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[508]), .O ({new_AGEMA_signal_3278, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[509]), .O ({new_AGEMA_signal_3279, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[510]), .O ({new_AGEMA_signal_3280, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[88], ciphertext_s0[88]}), .I1 ({ciphertext_s1[89], ciphertext_s0[89]}), .I2 ({ciphertext_s1[90], ciphertext_s0[90]}), .I3 ({ciphertext_s1[91], ciphertext_s0[91]}), .I4 ({ciphertext_s1[92], ciphertext_s0[92]}), .I5 ({ciphertext_s1[93], ciphertext_s0[93]}), .clk (clk), .r (Fresh[511]), .O ({new_AGEMA_signal_3281, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[512]), .O ({new_AGEMA_signal_3282, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[513]), .O ({new_AGEMA_signal_3283, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[514]), .O ({new_AGEMA_signal_3284, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[515]), .O ({new_AGEMA_signal_3285, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[516]), .O ({new_AGEMA_signal_3286, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[517]), .O ({new_AGEMA_signal_3287, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[518]), .O ({new_AGEMA_signal_3288, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[519]), .O ({new_AGEMA_signal_3289, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[520]), .O ({new_AGEMA_signal_3290, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[521]), .O ({new_AGEMA_signal_3291, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[522]), .O ({new_AGEMA_signal_3292, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[523]), .O ({new_AGEMA_signal_3293, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[524]), .O ({new_AGEMA_signal_3294, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[525]), .O ({new_AGEMA_signal_3295, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[526]), .O ({new_AGEMA_signal_3296, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[527]), .O ({new_AGEMA_signal_3297, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[528]), .O ({new_AGEMA_signal_3298, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[529]), .O ({new_AGEMA_signal_3299, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[530]), .O ({new_AGEMA_signal_3300, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[531]), .O ({new_AGEMA_signal_3301, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[532]), .O ({new_AGEMA_signal_3302, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[533]), .O ({new_AGEMA_signal_3303, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[534]), .O ({new_AGEMA_signal_3304, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[535]), .O ({new_AGEMA_signal_3305, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[536]), .O ({new_AGEMA_signal_3306, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[537]), .O ({new_AGEMA_signal_3307, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[538]), .O ({new_AGEMA_signal_3308, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[539]), .O ({new_AGEMA_signal_3309, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[540]), .O ({new_AGEMA_signal_3310, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[541]), .O ({new_AGEMA_signal_3311, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[542]), .O ({new_AGEMA_signal_3312, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[96], ciphertext_s0[96]}), .I1 ({ciphertext_s1[97], ciphertext_s0[97]}), .I2 ({ciphertext_s1[98], ciphertext_s0[98]}), .I3 ({ciphertext_s1[99], ciphertext_s0[99]}), .I4 ({ciphertext_s1[100], ciphertext_s0[100]}), .I5 ({ciphertext_s1[101], ciphertext_s0[101]}), .clk (clk), .r (Fresh[543]), .O ({new_AGEMA_signal_3313, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[544]), .O ({new_AGEMA_signal_3314, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[545]), .O ({new_AGEMA_signal_3315, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[546]), .O ({new_AGEMA_signal_3316, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[547]), .O ({new_AGEMA_signal_3317, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[548]), .O ({new_AGEMA_signal_3318, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[549]), .O ({new_AGEMA_signal_3319, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[550]), .O ({new_AGEMA_signal_3320, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[551]), .O ({new_AGEMA_signal_3321, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[552]), .O ({new_AGEMA_signal_3322, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[553]), .O ({new_AGEMA_signal_3323, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[554]), .O ({new_AGEMA_signal_3324, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[555]), .O ({new_AGEMA_signal_3325, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[556]), .O ({new_AGEMA_signal_3326, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[557]), .O ({new_AGEMA_signal_3327, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[558]), .O ({new_AGEMA_signal_3328, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[559]), .O ({new_AGEMA_signal_3329, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[560]), .O ({new_AGEMA_signal_3330, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[561]), .O ({new_AGEMA_signal_3331, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[562]), .O ({new_AGEMA_signal_3332, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[563]), .O ({new_AGEMA_signal_3333, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[564]), .O ({new_AGEMA_signal_3334, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[565]), .O ({new_AGEMA_signal_3335, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[566]), .O ({new_AGEMA_signal_3336, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[567]), .O ({new_AGEMA_signal_3337, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[568]), .O ({new_AGEMA_signal_3338, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[569]), .O ({new_AGEMA_signal_3339, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[570]), .O ({new_AGEMA_signal_3340, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[571]), .O ({new_AGEMA_signal_3341, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[572]), .O ({new_AGEMA_signal_3342, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[573]), .O ({new_AGEMA_signal_3343, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[574]), .O ({new_AGEMA_signal_3344, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[104], ciphertext_s0[104]}), .I1 ({ciphertext_s1[105], ciphertext_s0[105]}), .I2 ({ciphertext_s1[106], ciphertext_s0[106]}), .I3 ({ciphertext_s1[107], ciphertext_s0[107]}), .I4 ({ciphertext_s1[108], ciphertext_s0[108]}), .I5 ({ciphertext_s1[109], ciphertext_s0[109]}), .clk (clk), .r (Fresh[575]), .O ({new_AGEMA_signal_3345, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[576]), .O ({new_AGEMA_signal_3346, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[577]), .O ({new_AGEMA_signal_3347, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[578]), .O ({new_AGEMA_signal_3348, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[579]), .O ({new_AGEMA_signal_3349, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[580]), .O ({new_AGEMA_signal_3350, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[581]), .O ({new_AGEMA_signal_3351, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[582]), .O ({new_AGEMA_signal_3352, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[583]), .O ({new_AGEMA_signal_3353, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[584]), .O ({new_AGEMA_signal_3354, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[585]), .O ({new_AGEMA_signal_3355, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[586]), .O ({new_AGEMA_signal_3356, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[587]), .O ({new_AGEMA_signal_3357, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[588]), .O ({new_AGEMA_signal_3358, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[589]), .O ({new_AGEMA_signal_3359, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[590]), .O ({new_AGEMA_signal_3360, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[591]), .O ({new_AGEMA_signal_3361, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[592]), .O ({new_AGEMA_signal_3362, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[593]), .O ({new_AGEMA_signal_3363, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[594]), .O ({new_AGEMA_signal_3364, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[595]), .O ({new_AGEMA_signal_3365, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[596]), .O ({new_AGEMA_signal_3366, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[597]), .O ({new_AGEMA_signal_3367, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[598]), .O ({new_AGEMA_signal_3368, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[599]), .O ({new_AGEMA_signal_3369, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[600]), .O ({new_AGEMA_signal_3370, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[601]), .O ({new_AGEMA_signal_3371, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[602]), .O ({new_AGEMA_signal_3372, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[603]), .O ({new_AGEMA_signal_3373, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[604]), .O ({new_AGEMA_signal_3374, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[605]), .O ({new_AGEMA_signal_3375, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[606]), .O ({new_AGEMA_signal_3376, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[112], ciphertext_s0[112]}), .I1 ({ciphertext_s1[113], ciphertext_s0[113]}), .I2 ({ciphertext_s1[114], ciphertext_s0[114]}), .I3 ({ciphertext_s1[115], ciphertext_s0[115]}), .I4 ({ciphertext_s1[116], ciphertext_s0[116]}), .I5 ({ciphertext_s1[117], ciphertext_s0[117]}), .clk (clk), .r (Fresh[607]), .O ({new_AGEMA_signal_3377, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB14EDE67096C6EED ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[608]), .O ({new_AGEMA_signal_3378, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h68AB4BFA8ACB7A13 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[609]), .O ({new_AGEMA_signal_3379, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h10BDB210C006EAB5 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[610]), .O ({new_AGEMA_signal_3380, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4F1EAD396F247A04 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[611]), .O ({new_AGEMA_signal_3381, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7BAE007D4C53FC7D ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[612]), .O ({new_AGEMA_signal_3382, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE61A4C5E97816F7A ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[613]), .O ({new_AGEMA_signal_3383, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6A450B2EF33486B4 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[614]), .O ({new_AGEMA_signal_3384, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC870974094EAD8A9 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[615]), .O ({new_AGEMA_signal_3385, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hA16387FB3B48B4C6 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[616]), .O ({new_AGEMA_signal_3386, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h23A869A2A428C424 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[617]), .O ({new_AGEMA_signal_3387, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h577D64E03B0C3FFB ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[618]), .O ({new_AGEMA_signal_3388, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hAC39B6C0D6CE2EFC ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[619]), .O ({new_AGEMA_signal_3389, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h109020A2193D586A ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[620]), .O ({new_AGEMA_signal_3390, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2568EA2EFFA8527D ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[621]), .O ({new_AGEMA_signal_3391, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE9DA849CF6AC6C1B ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[622]), .O ({new_AGEMA_signal_3392, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4E9DDB76C892FB1B ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[623]), .O ({new_AGEMA_signal_3393, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hC2B0F97752B8B11E ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[624]), .O ({new_AGEMA_signal_3394, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF7F17A494CE30F58 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[625]), .O ({new_AGEMA_signal_3395, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h2624B286BC48ECB4 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[626]), .O ({new_AGEMA_signal_3396, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF210A3AECE472E53 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[627]), .O ({new_AGEMA_signal_3397, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hF8045F7B6D98DD7F ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[628]), .O ({new_AGEMA_signal_3398, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6BC2AA4E0D787AA4 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[629]), .O ({new_AGEMA_signal_3399, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h7D8DCC4706319E08 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[630]), .O ({new_AGEMA_signal_3400, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h54B248130B4F256F ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[631]), .O ({new_AGEMA_signal_3401, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h980A3CC2C2FDB4FF ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[632]), .O ({new_AGEMA_signal_3402, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE4851B3BF3AB2560 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[633]), .O ({new_AGEMA_signal_3403, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h3F6BCB91B30DB559 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[634]), .O ({new_AGEMA_signal_3404, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h21E0B83325591782 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[635]), .O ({new_AGEMA_signal_3405, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<3> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5CAA2EC7BF977090 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7_0 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[636]), .O ({new_AGEMA_signal_3406, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<0> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hE7BAC28F866AAC82 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7_1 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[637]), .O ({new_AGEMA_signal_3407, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<1> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4CB3770196CA0329 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7_2 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[638]), .O ({new_AGEMA_signal_3408, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<2> }) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'h52379DE7B844E3E1 ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7_3 ( .I0 ({ciphertext_s1[120], ciphertext_s0[120]}), .I1 ({ciphertext_s1[121], ciphertext_s0[121]}), .I2 ({ciphertext_s1[122], ciphertext_s0[122]}), .I3 ({ciphertext_s1[123], ciphertext_s0[123]}), .I4 ({ciphertext_s1[124], ciphertext_s0[124]}), .I5 ({ciphertext_s1[125], ciphertext_s0[125]}), .clk (clk), .r (Fresh[639]), .O ({new_AGEMA_signal_3409, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<3> }) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2315, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2314, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2313, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2312, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b7<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[640]), .O ({new_AGEMA_signal_2866, \KeyExpansionIns/tmp [7]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2319, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2318, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2317, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2316, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b6<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[641]), .O ({new_AGEMA_signal_2867, \KeyExpansionIns/tmp [6]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2323, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2322, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2321, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2320, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b5<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[642]), .O ({new_AGEMA_signal_2868, \KeyExpansionIns/tmp [5]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2327, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2326, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2325, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2324, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b4<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[643]), .O ({new_AGEMA_signal_2869, \KeyExpansionIns/tmp [4]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2331, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2330, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2329, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2328, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b3<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[644]), .O ({new_AGEMA_signal_2870, \KeyExpansionIns/tmp [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2335, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2334, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2333, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2332, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b2<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[645]), .O ({new_AGEMA_signal_2871, \KeyExpansionIns/tmp [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2339, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2338, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2337, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2336, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b1<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[646]), .O ({new_AGEMA_signal_2872, \KeyExpansionIns/tmp [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2343, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2342, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2341, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2340, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[3].Inst_Sbox/b0<3> }), .I4 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I5 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .clk (clk), .r (Fresh[647]), .O ({new_AGEMA_signal_2873, \KeyExpansionIns/tmp [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2353, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2352, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2351, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2350, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b7<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[648]), .O ({new_AGEMA_signal_2874, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [7]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2357, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2356, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2355, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2354, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b6<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[649]), .O ({new_AGEMA_signal_2875, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [6]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2361, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2360, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2359, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2358, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b5<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[650]), .O ({new_AGEMA_signal_2876, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [5]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2365, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2364, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2363, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2362, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b4<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[651]), .O ({new_AGEMA_signal_2877, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [4]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2369, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2368, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2367, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2366, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b3<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[652]), .O ({new_AGEMA_signal_2878, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2373, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2372, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2371, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2370, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b2<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[653]), .O ({new_AGEMA_signal_2879, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2377, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2376, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2375, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2374, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b1<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[654]), .O ({new_AGEMA_signal_2880, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2381, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2380, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2379, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2378, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[0].Inst_Sbox/b0<3> }), .I4 ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }), .I5 ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }), .clk (clk), .r (Fresh[655]), .O ({new_AGEMA_signal_2881, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2391, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2390, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2389, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2388, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b7<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[656]), .O ({new_AGEMA_signal_2882, \KeyExpansionIns/tmp [23]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2395, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2394, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2393, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2392, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b6<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[657]), .O ({new_AGEMA_signal_2883, \KeyExpansionIns/tmp [22]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2399, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2398, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2397, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2396, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b5<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[658]), .O ({new_AGEMA_signal_2884, \KeyExpansionIns/tmp [21]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2403, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2402, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2401, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2400, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b4<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[659]), .O ({new_AGEMA_signal_2885, \KeyExpansionIns/tmp [20]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2407, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2406, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2405, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2404, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b3<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[660]), .O ({new_AGEMA_signal_2886, \KeyExpansionIns/tmp [19]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2411, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2410, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2409, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2408, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b2<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[661]), .O ({new_AGEMA_signal_2887, \KeyExpansionIns/tmp [18]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2415, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2414, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2413, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2412, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b1<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[662]), .O ({new_AGEMA_signal_2888, \KeyExpansionIns/tmp [17]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2419, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2418, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2417, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2416, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[1].Inst_Sbox/b0<3> }), .I4 ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }), .I5 ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }), .clk (clk), .r (Fresh[663]), .O ({new_AGEMA_signal_2889, \KeyExpansionIns/tmp [16]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2429, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2428, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2427, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2426, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b7<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[664]), .O ({new_AGEMA_signal_2890, \KeyExpansionIns/tmp [15]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2433, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2432, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2431, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2430, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b6<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[665]), .O ({new_AGEMA_signal_2891, \KeyExpansionIns/tmp [14]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2437, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2436, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2435, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2434, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b5<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[666]), .O ({new_AGEMA_signal_2892, \KeyExpansionIns/tmp [13]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2441, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2440, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2439, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2438, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b4<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[667]), .O ({new_AGEMA_signal_2893, \KeyExpansionIns/tmp [12]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2445, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2444, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2443, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2442, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b3<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[668]), .O ({new_AGEMA_signal_2894, \KeyExpansionIns/tmp [11]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2449, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2448, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2447, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2446, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b2<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[669]), .O ({new_AGEMA_signal_2895, \KeyExpansionIns/tmp [10]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2453, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2452, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2451, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2450, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b1<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[670]), .O ({new_AGEMA_signal_2896, \KeyExpansionIns/tmp [9]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2457, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2456, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2455, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2454, \KeyExpansionIns/KeySchedCoreInst/GenSubBytes[2].Inst_Sbox/b0<3> }), .I4 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I5 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .clk (clk), .r (Fresh[671]), .O ({new_AGEMA_signal_2897, \KeyExpansionIns/tmp [8]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2898, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2899, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2900, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2901, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[672]), .O ({new_AGEMA_signal_3410, ShiftRowsInput[0]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2902, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2903, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2904, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2905, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[673]), .O ({new_AGEMA_signal_3411, ShiftRowsInput[1]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2906, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2907, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2908, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2909, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[674]), .O ({new_AGEMA_signal_3412, ShiftRowsInput[2]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2910, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2911, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2912, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2913, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[675]), .O ({new_AGEMA_signal_3413, ShiftRowsInput[3]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2914, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2915, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2916, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2917, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[676]), .O ({new_AGEMA_signal_3414, ShiftRowsInput[4]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2918, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2919, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2920, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2921, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[677]), .O ({new_AGEMA_signal_3415, ShiftRowsInput[5]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2922, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2923, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2924, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2925, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[678]), .O ({new_AGEMA_signal_3416, ShiftRowsInput[6]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2926, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2927, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2928, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2929, \SubBytesIns/GenSubBytes[0].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[6], ciphertext_s0[6]}), .I5 ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[679]), .O ({new_AGEMA_signal_3417, ShiftRowsInput[7]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2930, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2931, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2932, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2933, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[680]), .O ({new_AGEMA_signal_3418, ShiftRowsInput[8]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2934, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2935, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2936, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2937, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[681]), .O ({new_AGEMA_signal_3419, ShiftRowsInput[9]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2938, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2939, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2940, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2941, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[682]), .O ({new_AGEMA_signal_3420, ShiftRowsInput[10]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2942, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2943, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2944, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2945, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[683]), .O ({new_AGEMA_signal_3421, ShiftRowsInput[11]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2946, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2947, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2948, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2949, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[684]), .O ({new_AGEMA_signal_3422, ShiftRowsInput[12]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2950, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2951, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2952, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2953, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[685]), .O ({new_AGEMA_signal_3423, ShiftRowsInput[13]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2954, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2955, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2956, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2957, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[686]), .O ({new_AGEMA_signal_3424, ShiftRowsInput[14]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2958, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2959, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2960, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2961, \SubBytesIns/GenSubBytes[1].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[14], ciphertext_s0[14]}), .I5 ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[687]), .O ({new_AGEMA_signal_3425, ShiftRowsInput[15]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2962, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2963, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2964, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2965, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[688]), .O ({new_AGEMA_signal_3426, ShiftRowsInput[16]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2966, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2967, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_2968, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_2969, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[689]), .O ({new_AGEMA_signal_3427, ShiftRowsInput[17]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_2970, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_2971, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_2972, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_2973, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[690]), .O ({new_AGEMA_signal_3428, ShiftRowsInput[18]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_2974, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_2975, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_2976, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_2977, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[691]), .O ({new_AGEMA_signal_3429, ShiftRowsInput[19]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_2978, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_2979, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_2980, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_2981, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[692]), .O ({new_AGEMA_signal_3430, ShiftRowsInput[20]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_2982, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_2983, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_2984, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_2985, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[693]), .O ({new_AGEMA_signal_3431, ShiftRowsInput[21]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_2986, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_2987, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_2988, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_2989, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[694]), .O ({new_AGEMA_signal_3432, ShiftRowsInput[22]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_2990, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_2991, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_2992, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_2993, \SubBytesIns/GenSubBytes[2].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[22], ciphertext_s0[22]}), .I5 ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[695]), .O ({new_AGEMA_signal_3433, ShiftRowsInput[23]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_2994, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_2995, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_2996, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_2997, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[696]), .O ({new_AGEMA_signal_3434, ShiftRowsInput[24]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_2998, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_2999, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3000, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3001, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[697]), .O ({new_AGEMA_signal_3435, ShiftRowsInput[25]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3002, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3003, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3004, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3005, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[698]), .O ({new_AGEMA_signal_3436, ShiftRowsInput[26]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3006, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3007, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3008, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3009, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[699]), .O ({new_AGEMA_signal_3437, ShiftRowsInput[27]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3010, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3011, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3012, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3013, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[700]), .O ({new_AGEMA_signal_3438, ShiftRowsInput[28]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3014, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3015, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3016, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3017, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[701]), .O ({new_AGEMA_signal_3439, ShiftRowsInput[29]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3018, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3019, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3020, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3021, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[702]), .O ({new_AGEMA_signal_3440, ShiftRowsInput[30]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3022, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3023, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3024, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3025, \SubBytesIns/GenSubBytes[3].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[30], ciphertext_s0[30]}), .I5 ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[703]), .O ({new_AGEMA_signal_3441, ShiftRowsInput[31]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3026, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3027, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3028, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3029, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[704]), .O ({new_AGEMA_signal_3442, ShiftRowsInput[32]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3030, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3031, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3032, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3033, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[705]), .O ({new_AGEMA_signal_3443, ShiftRowsInput[33]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3034, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3035, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3036, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3037, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[706]), .O ({new_AGEMA_signal_3444, ShiftRowsInput[34]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3038, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3039, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3040, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3041, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[707]), .O ({new_AGEMA_signal_3445, ShiftRowsInput[35]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3042, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3043, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3044, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3045, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[708]), .O ({new_AGEMA_signal_3446, ShiftRowsInput[36]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3046, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3047, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3048, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3049, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[709]), .O ({new_AGEMA_signal_3447, ShiftRowsInput[37]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3050, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3051, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3052, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3053, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[710]), .O ({new_AGEMA_signal_3448, ShiftRowsInput[38]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3054, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3055, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3056, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3057, \SubBytesIns/GenSubBytes[4].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[38], ciphertext_s0[38]}), .I5 ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[711]), .O ({new_AGEMA_signal_3449, ShiftRowsInput[39]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3058, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3059, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3060, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3061, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[712]), .O ({new_AGEMA_signal_3450, ShiftRowsInput[40]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3062, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3063, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3064, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3065, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[713]), .O ({new_AGEMA_signal_3451, ShiftRowsInput[41]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3066, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3067, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3068, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3069, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[714]), .O ({new_AGEMA_signal_3452, ShiftRowsInput[42]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3070, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3071, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3072, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3073, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[715]), .O ({new_AGEMA_signal_3453, ShiftRowsInput[43]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3074, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3075, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3076, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3077, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[716]), .O ({new_AGEMA_signal_3454, ShiftRowsInput[44]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3078, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3079, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3080, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3081, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[717]), .O ({new_AGEMA_signal_3455, ShiftRowsInput[45]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3082, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3083, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3084, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3085, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[718]), .O ({new_AGEMA_signal_3456, ShiftRowsInput[46]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3086, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3087, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3088, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3089, \SubBytesIns/GenSubBytes[5].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[46], ciphertext_s0[46]}), .I5 ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[719]), .O ({new_AGEMA_signal_3457, ShiftRowsInput[47]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3090, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3091, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3092, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3093, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[720]), .O ({new_AGEMA_signal_3458, ShiftRowsInput[48]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3094, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3095, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3096, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3097, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[721]), .O ({new_AGEMA_signal_3459, ShiftRowsInput[49]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3098, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3099, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3100, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3101, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[722]), .O ({new_AGEMA_signal_3460, ShiftRowsInput[50]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3102, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3103, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3104, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3105, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[723]), .O ({new_AGEMA_signal_3461, ShiftRowsInput[51]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3106, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3107, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3108, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3109, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[724]), .O ({new_AGEMA_signal_3462, ShiftRowsInput[52]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3110, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3111, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3112, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3113, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[725]), .O ({new_AGEMA_signal_3463, ShiftRowsInput[53]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3114, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3115, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3116, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3117, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[726]), .O ({new_AGEMA_signal_3464, ShiftRowsInput[54]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3118, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3119, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3120, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3121, \SubBytesIns/GenSubBytes[6].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[54], ciphertext_s0[54]}), .I5 ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[727]), .O ({new_AGEMA_signal_3465, ShiftRowsInput[55]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3122, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3123, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3124, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3125, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[728]), .O ({new_AGEMA_signal_3466, ShiftRowsInput[56]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3126, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3127, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3128, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3129, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[729]), .O ({new_AGEMA_signal_3467, ShiftRowsInput[57]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3130, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3131, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3132, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3133, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[730]), .O ({new_AGEMA_signal_3468, ShiftRowsInput[58]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3134, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3135, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3136, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3137, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[731]), .O ({new_AGEMA_signal_3469, ShiftRowsInput[59]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3138, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3139, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3140, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3141, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[732]), .O ({new_AGEMA_signal_3470, ShiftRowsInput[60]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3142, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3143, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3144, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3145, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[733]), .O ({new_AGEMA_signal_3471, ShiftRowsInput[61]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3146, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3147, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3148, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3149, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[734]), .O ({new_AGEMA_signal_3472, ShiftRowsInput[62]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3150, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3151, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3152, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3153, \SubBytesIns/GenSubBytes[7].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[62], ciphertext_s0[62]}), .I5 ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[735]), .O ({new_AGEMA_signal_3473, ShiftRowsInput[63]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3154, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3155, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3156, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3157, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[736]), .O ({new_AGEMA_signal_3474, ShiftRowsInput[64]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3158, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3159, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3160, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3161, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[737]), .O ({new_AGEMA_signal_3475, ShiftRowsInput[65]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3162, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3163, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3164, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3165, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[738]), .O ({new_AGEMA_signal_3476, ShiftRowsInput[66]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3166, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3167, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3168, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3169, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[739]), .O ({new_AGEMA_signal_3477, ShiftRowsInput[67]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3170, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3171, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3172, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3173, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[740]), .O ({new_AGEMA_signal_3478, ShiftRowsInput[68]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3174, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3175, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3176, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3177, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[741]), .O ({new_AGEMA_signal_3479, ShiftRowsInput[69]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3178, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3179, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3180, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3181, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[742]), .O ({new_AGEMA_signal_3480, ShiftRowsInput[70]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3182, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3183, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3184, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3185, \SubBytesIns/GenSubBytes[8].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[70], ciphertext_s0[70]}), .I5 ({ciphertext_s1[71], ciphertext_s0[71]}), .clk (clk), .r (Fresh[743]), .O ({new_AGEMA_signal_3481, ShiftRowsInput[71]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3186, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3187, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3188, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3189, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[744]), .O ({new_AGEMA_signal_3482, ShiftRowsInput[72]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3190, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3191, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3192, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3193, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[745]), .O ({new_AGEMA_signal_3483, ShiftRowsInput[73]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3194, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3195, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3196, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3197, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[746]), .O ({new_AGEMA_signal_3484, ShiftRowsInput[74]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3198, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3199, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3200, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3201, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[747]), .O ({new_AGEMA_signal_3485, ShiftRowsInput[75]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3202, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3203, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3204, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3205, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[748]), .O ({new_AGEMA_signal_3486, ShiftRowsInput[76]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3206, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3207, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3208, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3209, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[749]), .O ({new_AGEMA_signal_3487, ShiftRowsInput[77]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3210, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3211, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3212, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3213, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[750]), .O ({new_AGEMA_signal_3488, ShiftRowsInput[78]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3214, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3215, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3216, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3217, \SubBytesIns/GenSubBytes[9].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[78], ciphertext_s0[78]}), .I5 ({ciphertext_s1[79], ciphertext_s0[79]}), .clk (clk), .r (Fresh[751]), .O ({new_AGEMA_signal_3489, ShiftRowsInput[79]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3218, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3219, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3220, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3221, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[752]), .O ({new_AGEMA_signal_3490, ShiftRowsInput[80]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3222, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3223, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3224, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3225, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[753]), .O ({new_AGEMA_signal_3491, ShiftRowsInput[81]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3226, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3227, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3228, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3229, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[754]), .O ({new_AGEMA_signal_3492, ShiftRowsInput[82]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3230, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3231, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3232, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3233, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[755]), .O ({new_AGEMA_signal_3493, ShiftRowsInput[83]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3234, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3235, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3236, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3237, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[756]), .O ({new_AGEMA_signal_3494, ShiftRowsInput[84]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3238, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3239, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3240, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3241, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[757]), .O ({new_AGEMA_signal_3495, ShiftRowsInput[85]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3242, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3243, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3244, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3245, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[758]), .O ({new_AGEMA_signal_3496, ShiftRowsInput[86]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3246, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3247, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3248, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3249, \SubBytesIns/GenSubBytes[10].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[86], ciphertext_s0[86]}), .I5 ({ciphertext_s1[87], ciphertext_s0[87]}), .clk (clk), .r (Fresh[759]), .O ({new_AGEMA_signal_3497, ShiftRowsInput[87]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3250, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3251, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3252, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3253, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[760]), .O ({new_AGEMA_signal_3498, ShiftRowsInput[88]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3254, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3255, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3256, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3257, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[761]), .O ({new_AGEMA_signal_3499, ShiftRowsInput[89]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3258, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3259, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3260, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3261, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[762]), .O ({new_AGEMA_signal_3500, ShiftRowsInput[90]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3262, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3263, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3264, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3265, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[763]), .O ({new_AGEMA_signal_3501, ShiftRowsInput[91]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3266, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3267, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3268, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3269, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[764]), .O ({new_AGEMA_signal_3502, ShiftRowsInput[92]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3270, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3271, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3272, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3273, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[765]), .O ({new_AGEMA_signal_3503, ShiftRowsInput[93]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3274, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3275, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3276, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3277, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[766]), .O ({new_AGEMA_signal_3504, ShiftRowsInput[94]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3278, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3279, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3280, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3281, \SubBytesIns/GenSubBytes[11].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[94], ciphertext_s0[94]}), .I5 ({ciphertext_s1[95], ciphertext_s0[95]}), .clk (clk), .r (Fresh[767]), .O ({new_AGEMA_signal_3505, ShiftRowsInput[95]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3282, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3283, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3284, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3285, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[768]), .O ({new_AGEMA_signal_3506, ShiftRowsInput[96]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3286, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3287, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3288, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3289, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[769]), .O ({new_AGEMA_signal_3507, ShiftRowsInput[97]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3290, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3291, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3292, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3293, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[770]), .O ({new_AGEMA_signal_3508, ShiftRowsInput[98]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3294, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3295, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3296, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3297, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[771]), .O ({new_AGEMA_signal_3509, ShiftRowsInput[99]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3298, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3299, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3300, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3301, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[772]), .O ({new_AGEMA_signal_3510, ShiftRowsInput[100]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3302, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3303, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3304, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3305, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[773]), .O ({new_AGEMA_signal_3511, ShiftRowsInput[101]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3306, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3307, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3308, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3309, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[774]), .O ({new_AGEMA_signal_3512, ShiftRowsInput[102]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3310, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3311, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3312, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3313, \SubBytesIns/GenSubBytes[12].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[102], ciphertext_s0[102]}), .I5 ({ciphertext_s1[103], ciphertext_s0[103]}), .clk (clk), .r (Fresh[775]), .O ({new_AGEMA_signal_3513, ShiftRowsInput[103]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3314, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3315, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3316, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3317, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[776]), .O ({new_AGEMA_signal_3514, ShiftRowsInput[104]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3318, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3319, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3320, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3321, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[777]), .O ({new_AGEMA_signal_3515, ShiftRowsInput[105]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3322, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3323, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3324, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3325, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[778]), .O ({new_AGEMA_signal_3516, ShiftRowsInput[106]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3326, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3327, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3328, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3329, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[779]), .O ({new_AGEMA_signal_3517, ShiftRowsInput[107]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3330, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3331, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3332, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3333, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[780]), .O ({new_AGEMA_signal_3518, ShiftRowsInput[108]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3334, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3335, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3336, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3337, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[781]), .O ({new_AGEMA_signal_3519, ShiftRowsInput[109]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3338, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3339, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3340, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3341, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[782]), .O ({new_AGEMA_signal_3520, ShiftRowsInput[110]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3342, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3343, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3344, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3345, \SubBytesIns/GenSubBytes[13].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[110], ciphertext_s0[110]}), .I5 ({ciphertext_s1[111], ciphertext_s0[111]}), .clk (clk), .r (Fresh[783]), .O ({new_AGEMA_signal_3521, ShiftRowsInput[111]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3346, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3347, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3348, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3349, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[784]), .O ({new_AGEMA_signal_3522, ShiftRowsInput[112]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3350, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3351, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3352, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3353, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[785]), .O ({new_AGEMA_signal_3523, ShiftRowsInput[113]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3354, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3355, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3356, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3357, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[786]), .O ({new_AGEMA_signal_3524, ShiftRowsInput[114]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3358, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3359, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3360, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3361, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[787]), .O ({new_AGEMA_signal_3525, ShiftRowsInput[115]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3362, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3363, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3364, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3365, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[788]), .O ({new_AGEMA_signal_3526, ShiftRowsInput[116]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3366, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3367, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3368, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3369, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[789]), .O ({new_AGEMA_signal_3527, ShiftRowsInput[117]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3370, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3371, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3372, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3373, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[790]), .O ({new_AGEMA_signal_3528, ShiftRowsInput[118]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3374, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3375, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3376, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3377, \SubBytesIns/GenSubBytes[14].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[118], ciphertext_s0[118]}), .I5 ({ciphertext_s1[119], ciphertext_s0[119]}), .clk (clk), .r (Fresh[791]), .O ({new_AGEMA_signal_3529, ShiftRowsInput[119]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0_4 ( .I0 ({new_AGEMA_signal_3378, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<0> }), .I1 ({new_AGEMA_signal_3379, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<1> }), .I2 ({new_AGEMA_signal_3380, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<2> }), .I3 ({new_AGEMA_signal_3381, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b0<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[792]), .O ({new_AGEMA_signal_3530, ShiftRowsInput[120]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1_4 ( .I0 ({new_AGEMA_signal_3382, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<0> }), .I1 ({new_AGEMA_signal_3383, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<1> }), .I2 ({new_AGEMA_signal_3384, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<2> }), .I3 ({new_AGEMA_signal_3385, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b1<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[793]), .O ({new_AGEMA_signal_3531, ShiftRowsInput[121]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2_4 ( .I0 ({new_AGEMA_signal_3386, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<0> }), .I1 ({new_AGEMA_signal_3387, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<1> }), .I2 ({new_AGEMA_signal_3388, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<2> }), .I3 ({new_AGEMA_signal_3389, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b2<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[794]), .O ({new_AGEMA_signal_3532, ShiftRowsInput[122]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3_4 ( .I0 ({new_AGEMA_signal_3390, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<0> }), .I1 ({new_AGEMA_signal_3391, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<1> }), .I2 ({new_AGEMA_signal_3392, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<2> }), .I3 ({new_AGEMA_signal_3393, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b3<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[795]), .O ({new_AGEMA_signal_3533, ShiftRowsInput[123]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4_4 ( .I0 ({new_AGEMA_signal_3394, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<0> }), .I1 ({new_AGEMA_signal_3395, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<1> }), .I2 ({new_AGEMA_signal_3396, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<2> }), .I3 ({new_AGEMA_signal_3397, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b4<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[796]), .O ({new_AGEMA_signal_3534, ShiftRowsInput[124]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5_4 ( .I0 ({new_AGEMA_signal_3398, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<0> }), .I1 ({new_AGEMA_signal_3399, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<1> }), .I2 ({new_AGEMA_signal_3400, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<2> }), .I3 ({new_AGEMA_signal_3401, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b5<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[797]), .O ({new_AGEMA_signal_3535, ShiftRowsInput[125]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6_4 ( .I0 ({new_AGEMA_signal_3402, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<0> }), .I1 ({new_AGEMA_signal_3403, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<1> }), .I2 ({new_AGEMA_signal_3404, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<2> }), .I3 ({new_AGEMA_signal_3405, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b6<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[798]), .O ({new_AGEMA_signal_3536, ShiftRowsInput[126]}) ) ;
    LUT6_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 64'hFF00F0F0CCCCAAAA ) ) \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7_4 ( .I0 ({new_AGEMA_signal_3406, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<0> }), .I1 ({new_AGEMA_signal_3407, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<1> }), .I2 ({new_AGEMA_signal_3408, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<2> }), .I3 ({new_AGEMA_signal_3409, \SubBytesIns/GenSubBytes[15].Inst_Sbox/b7<3> }), .I4 ({ciphertext_s1[126], ciphertext_s0[126]}), .I5 ({ciphertext_s1[127], ciphertext_s0[127]}), .clk (clk), .r (Fresh[799]), .O ({new_AGEMA_signal_3537, ShiftRowsInput[127]}) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_4_xo<0>1 ( .I0 ({new_AGEMA_signal_3413, ShiftRowsInput[3]}), .I1 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3754, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><4> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_1_xo<0>1 ( .I0 ({new_AGEMA_signal_3442, ShiftRowsInput[32]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .O ({new_AGEMA_signal_3755, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><1> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_3_xo<0>1 ( .I0 ({new_AGEMA_signal_3444, ShiftRowsInput[34]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .O ({new_AGEMA_signal_3756, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><3> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_1_xo<0>1 ( .I0 ({new_AGEMA_signal_3474, ShiftRowsInput[64]}), .I1 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .O ({new_AGEMA_signal_3757, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><1> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_3_xo<0>1 ( .I0 ({new_AGEMA_signal_3476, ShiftRowsInput[66]}), .I1 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .O ({new_AGEMA_signal_3758, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><3> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_4_xo<0>1 ( .I0 ({new_AGEMA_signal_3477, ShiftRowsInput[67]}), .I1 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .O ({new_AGEMA_signal_3759, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><4> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_4_xo<0>1 ( .I0 ({new_AGEMA_signal_3445, ShiftRowsInput[35]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .O ({new_AGEMA_signal_3760, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><4> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_1_xo<0>1 ( .I0 ({new_AGEMA_signal_3506, ShiftRowsInput[96]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .O ({new_AGEMA_signal_3761, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><1> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_3_xo<0>1 ( .I0 ({new_AGEMA_signal_3508, ShiftRowsInput[98]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .O ({new_AGEMA_signal_3762, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><3> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_4_xo<0>1 ( .I0 ({new_AGEMA_signal_3509, ShiftRowsInput[99]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .O ({new_AGEMA_signal_3763, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><4> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_1_xo<0>1 ( .I0 ({new_AGEMA_signal_3410, ShiftRowsInput[0]}), .I1 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3764, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><1> }) ) ;
    LUT2_masked #(.low_latency(0), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/GenMul2[3].Mul2Inst/Mxor_output_3_xo<0>1 ( .I0 ({new_AGEMA_signal_3412, ShiftRowsInput[2]}), .I1 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3765, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><3> }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h5556AAA9 ) , .MASK ( 5'b01110 ), .INIT2 ( 32'h5555AAAA ) ) \KeyExpansionOutput<24>31 ( .I0 ({new_AGEMA_signal_2480, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_393 }), .I1 ({1'b0, \RoundCounterIns/count [2]}), .I2 ({1'b0, \RoundCounterIns/count [1]}), .I3 ({1'b0, \RoundCounterIns/count [0]}), .I4 ({new_AGEMA_signal_2881, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [0]}), .O ({new_AGEMA_signal_3538, \KeyExpansionOutput<24>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h56555559A9AAAAA6 ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<27>31 ( .I0 ({new_AGEMA_signal_2471, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_390 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2878, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [3]}), .O ({new_AGEMA_signal_3539, \KeyExpansionOutput<27>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h655555559AAAAAAA ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<31>31 ( .I0 ({new_AGEMA_signal_2459, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_386 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2874, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [7]}), .O ({new_AGEMA_signal_3540, \KeyExpansionOutput<31>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h55556555AAAA9AAA ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<30>31 ( .I0 ({new_AGEMA_signal_2462, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_387 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2875, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [6]}), .O ({new_AGEMA_signal_3541, \KeyExpansionOutput<30>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h55595569AAA6AA96 ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<28>31 ( .I0 ({new_AGEMA_signal_2468, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_389 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2877, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [4]}), .O ({new_AGEMA_signal_3542, \KeyExpansionOutput<28>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h55695555AA96AAAA ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<29>31 ( .I0 ({new_AGEMA_signal_2465, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_388 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2876, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [5]}), .O ({new_AGEMA_signal_3543, \KeyExpansionOutput<29>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h555A5559AAA5AAA6 ) , .MASK ( 6'b011110 ), .INIT2 ( 64'h55555555AAAAAAAA ) ) \KeyExpansionOutput<25>31 ( .I0 ({new_AGEMA_signal_2477, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_392 }), .I1 ({1'b0, \RoundCounterIns/count [3]}), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, \RoundCounterIns/count [0]}), .I5 ({new_AGEMA_signal_2880, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [1]}), .O ({new_AGEMA_signal_3544, \KeyExpansionOutput<25>_bdd4 }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[24], key_s0[24]}), .I2 ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }), .I3 ({new_AGEMA_signal_2672, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_457 }), .I4 ({new_AGEMA_signal_2576, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 }), .I5 ({new_AGEMA_signal_3538, \KeyExpansionOutput<24>_bdd4 }), .O ({new_AGEMA_signal_3767, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[25], key_s0[25]}), .I2 ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }), .I3 ({new_AGEMA_signal_2669, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_456 }), .I4 ({new_AGEMA_signal_2573, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 }), .I5 ({new_AGEMA_signal_3544, \KeyExpansionOutput<25>_bdd4 }), .O ({new_AGEMA_signal_3769, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[27], key_s0[27]}), .I2 ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }), .I3 ({new_AGEMA_signal_2663, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_454 }), .I4 ({new_AGEMA_signal_2567, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 }), .I5 ({new_AGEMA_signal_3539, \KeyExpansionOutput<27>_bdd4 }), .O ({new_AGEMA_signal_3771, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[28], key_s0[28]}), .I2 ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }), .I3 ({new_AGEMA_signal_2660, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_453 }), .I4 ({new_AGEMA_signal_2564, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 }), .I5 ({new_AGEMA_signal_3542, \KeyExpansionOutput<28>_bdd4 }), .O ({new_AGEMA_signal_3773, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[29], key_s0[29]}), .I2 ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }), .I3 ({new_AGEMA_signal_2657, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_452 }), .I4 ({new_AGEMA_signal_2561, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 }), .I5 ({new_AGEMA_signal_3543, \KeyExpansionOutput<29>_bdd4 }), .O ({new_AGEMA_signal_3775, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[30], key_s0[30]}), .I2 ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }), .I3 ({new_AGEMA_signal_2654, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_451 }), .I4 ({new_AGEMA_signal_2558, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 }), .I5 ({new_AGEMA_signal_3541, \KeyExpansionOutput<30>_bdd4 }), .O ({new_AGEMA_signal_3777, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[31], key_s0[31]}), .I2 ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }), .I3 ({new_AGEMA_signal_2651, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_450 }), .I4 ({new_AGEMA_signal_2555, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 }), .I5 ({new_AGEMA_signal_3540, \KeyExpansionOutput<31>_bdd4 }), .O ({new_AGEMA_signal_3779, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[32], key_s0[32]}), .I2 ({new_AGEMA_signal_2744, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_481 }), .I3 ({new_AGEMA_signal_2648, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 }), .I4 ({new_AGEMA_signal_2873, \KeyExpansionIns/tmp [0]}), .I5 ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }), .O ({new_AGEMA_signal_3546, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[33], key_s0[33]}), .I2 ({new_AGEMA_signal_2741, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_480 }), .I3 ({new_AGEMA_signal_2645, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 }), .I4 ({new_AGEMA_signal_2872, \KeyExpansionIns/tmp [1]}), .I5 ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }), .O ({new_AGEMA_signal_3548, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[34], key_s0[34]}), .I2 ({new_AGEMA_signal_2738, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_479 }), .I3 ({new_AGEMA_signal_2642, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 }), .I4 ({new_AGEMA_signal_2871, \KeyExpansionIns/tmp [2]}), .I5 ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }), .O ({new_AGEMA_signal_3550, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[35], key_s0[35]}), .I2 ({new_AGEMA_signal_2735, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_478 }), .I3 ({new_AGEMA_signal_2639, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 }), .I4 ({new_AGEMA_signal_2870, \KeyExpansionIns/tmp [3]}), .I5 ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }), .O ({new_AGEMA_signal_3552, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[36], key_s0[36]}), .I2 ({new_AGEMA_signal_2732, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_477 }), .I3 ({new_AGEMA_signal_2636, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 }), .I4 ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }), .I5 ({new_AGEMA_signal_2869, \KeyExpansionIns/tmp [4]}), .O ({new_AGEMA_signal_3554, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[37], key_s0[37]}), .I2 ({new_AGEMA_signal_2729, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_476 }), .I3 ({new_AGEMA_signal_2633, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 }), .I4 ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }), .I5 ({new_AGEMA_signal_2868, \KeyExpansionIns/tmp [5]}), .O ({new_AGEMA_signal_3556, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[38], key_s0[38]}), .I2 ({new_AGEMA_signal_2726, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_475 }), .I3 ({new_AGEMA_signal_2630, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 }), .I4 ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }), .I5 ({new_AGEMA_signal_2867, \KeyExpansionIns/tmp [6]}), .O ({new_AGEMA_signal_3558, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[39], key_s0[39]}), .I2 ({new_AGEMA_signal_2723, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_474 }), .I3 ({new_AGEMA_signal_2627, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 }), .I4 ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }), .I5 ({new_AGEMA_signal_2866, \KeyExpansionIns/tmp [7]}), .O ({new_AGEMA_signal_3560, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[40], key_s0[40]}), .I2 ({new_AGEMA_signal_2720, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_473 }), .I3 ({new_AGEMA_signal_2624, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 }), .I4 ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }), .I5 ({new_AGEMA_signal_2897, \KeyExpansionIns/tmp [8]}), .O ({new_AGEMA_signal_3562, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[41], key_s0[41]}), .I2 ({new_AGEMA_signal_2717, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_472 }), .I3 ({new_AGEMA_signal_2621, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 }), .I4 ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }), .I5 ({new_AGEMA_signal_2896, \KeyExpansionIns/tmp [9]}), .O ({new_AGEMA_signal_3564, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[42], key_s0[42]}), .I2 ({new_AGEMA_signal_2714, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_471 }), .I3 ({new_AGEMA_signal_2618, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 }), .I4 ({new_AGEMA_signal_2895, \KeyExpansionIns/tmp [10]}), .I5 ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }), .O ({new_AGEMA_signal_3566, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[43], key_s0[43]}), .I2 ({new_AGEMA_signal_2711, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_470 }), .I3 ({new_AGEMA_signal_2615, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 }), .I4 ({new_AGEMA_signal_2894, \KeyExpansionIns/tmp [11]}), .I5 ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }), .O ({new_AGEMA_signal_3568, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[44], key_s0[44]}), .I2 ({new_AGEMA_signal_2708, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_469 }), .I3 ({new_AGEMA_signal_2612, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 }), .I4 ({new_AGEMA_signal_2893, \KeyExpansionIns/tmp [12]}), .I5 ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }), .O ({new_AGEMA_signal_3570, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[45], key_s0[45]}), .I2 ({new_AGEMA_signal_2705, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_468 }), .I3 ({new_AGEMA_signal_2609, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 }), .I4 ({new_AGEMA_signal_2892, \KeyExpansionIns/tmp [13]}), .I5 ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }), .O ({new_AGEMA_signal_3572, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[46], key_s0[46]}), .I2 ({new_AGEMA_signal_2702, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_467 }), .I3 ({new_AGEMA_signal_2606, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 }), .I4 ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }), .I5 ({new_AGEMA_signal_2891, \KeyExpansionIns/tmp [14]}), .O ({new_AGEMA_signal_3574, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[47], key_s0[47]}), .I2 ({new_AGEMA_signal_2699, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_466 }), .I3 ({new_AGEMA_signal_2603, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 }), .I4 ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }), .I5 ({new_AGEMA_signal_2890, \KeyExpansionIns/tmp [15]}), .O ({new_AGEMA_signal_3576, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[48], key_s0[48]}), .I2 ({new_AGEMA_signal_2696, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_465 }), .I3 ({new_AGEMA_signal_2600, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 }), .I4 ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }), .I5 ({new_AGEMA_signal_2889, \KeyExpansionIns/tmp [16]}), .O ({new_AGEMA_signal_3578, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[49], key_s0[49]}), .I2 ({new_AGEMA_signal_2693, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_464 }), .I3 ({new_AGEMA_signal_2597, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 }), .I4 ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }), .I5 ({new_AGEMA_signal_2888, \KeyExpansionIns/tmp [17]}), .O ({new_AGEMA_signal_3580, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[50], key_s0[50]}), .I2 ({new_AGEMA_signal_2690, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_463 }), .I3 ({new_AGEMA_signal_2594, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 }), .I4 ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }), .I5 ({new_AGEMA_signal_2887, \KeyExpansionIns/tmp [18]}), .O ({new_AGEMA_signal_3582, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[51], key_s0[51]}), .I2 ({new_AGEMA_signal_2687, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_462 }), .I3 ({new_AGEMA_signal_2591, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 }), .I4 ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }), .I5 ({new_AGEMA_signal_2886, \KeyExpansionIns/tmp [19]}), .O ({new_AGEMA_signal_3584, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[52], key_s0[52]}), .I2 ({new_AGEMA_signal_2684, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_461 }), .I3 ({new_AGEMA_signal_2588, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 }), .I4 ({new_AGEMA_signal_2885, \KeyExpansionIns/tmp [20]}), .I5 ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }), .O ({new_AGEMA_signal_3586, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[53], key_s0[53]}), .I2 ({new_AGEMA_signal_2681, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_460 }), .I3 ({new_AGEMA_signal_2585, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 }), .I4 ({new_AGEMA_signal_2884, \KeyExpansionIns/tmp [21]}), .I5 ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }), .O ({new_AGEMA_signal_3588, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[54], key_s0[54]}), .I2 ({new_AGEMA_signal_2678, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_459 }), .I3 ({new_AGEMA_signal_2582, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 }), .I4 ({new_AGEMA_signal_2883, \KeyExpansionIns/tmp [22]}), .I5 ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }), .O ({new_AGEMA_signal_3590, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[55], key_s0[55]}), .I2 ({new_AGEMA_signal_2675, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_458 }), .I3 ({new_AGEMA_signal_2579, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 }), .I4 ({new_AGEMA_signal_2882, \KeyExpansionIns/tmp [23]}), .I5 ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }), .O ({new_AGEMA_signal_3592, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[56], key_s0[56]}), .I2 ({new_AGEMA_signal_2672, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_457 }), .I3 ({new_AGEMA_signal_2576, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 }), .I4 ({new_AGEMA_signal_3538, \KeyExpansionOutput<24>_bdd4 }), .O ({new_AGEMA_signal_3781, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[57], key_s0[57]}), .I2 ({new_AGEMA_signal_2669, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_456 }), .I3 ({new_AGEMA_signal_2573, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 }), .I4 ({new_AGEMA_signal_3544, \KeyExpansionOutput<25>_bdd4 }), .O ({new_AGEMA_signal_3783, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[59], key_s0[59]}), .I2 ({new_AGEMA_signal_2663, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_454 }), .I3 ({new_AGEMA_signal_2567, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 }), .I4 ({new_AGEMA_signal_3539, \KeyExpansionOutput<27>_bdd4 }), .O ({new_AGEMA_signal_3785, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[60], key_s0[60]}), .I2 ({new_AGEMA_signal_2660, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_453 }), .I3 ({new_AGEMA_signal_2564, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 }), .I4 ({new_AGEMA_signal_3542, \KeyExpansionOutput<28>_bdd4 }), .O ({new_AGEMA_signal_3787, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[61], key_s0[61]}), .I2 ({new_AGEMA_signal_2657, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_452 }), .I3 ({new_AGEMA_signal_2561, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 }), .I4 ({new_AGEMA_signal_3543, \KeyExpansionOutput<29>_bdd4 }), .O ({new_AGEMA_signal_3789, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[62], key_s0[62]}), .I2 ({new_AGEMA_signal_2654, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_451 }), .I3 ({new_AGEMA_signal_2558, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 }), .I4 ({new_AGEMA_signal_3541, \KeyExpansionOutput<30>_bdd4 }), .O ({new_AGEMA_signal_3791, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[63], key_s0[63]}), .I2 ({new_AGEMA_signal_2651, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_450 }), .I3 ({new_AGEMA_signal_2555, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 }), .I4 ({new_AGEMA_signal_3540, \KeyExpansionOutput<31>_bdd4 }), .O ({new_AGEMA_signal_3793, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[64], key_s0[64]}), .I2 ({new_AGEMA_signal_2648, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 }), .I3 ({new_AGEMA_signal_2873, \KeyExpansionIns/tmp [0]}), .I4 ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }), .O ({new_AGEMA_signal_3594, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[65], key_s0[65]}), .I2 ({new_AGEMA_signal_2645, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 }), .I3 ({new_AGEMA_signal_2872, \KeyExpansionIns/tmp [1]}), .I4 ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }), .O ({new_AGEMA_signal_3596, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[66], key_s0[66]}), .I2 ({new_AGEMA_signal_2642, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 }), .I3 ({new_AGEMA_signal_2871, \KeyExpansionIns/tmp [2]}), .I4 ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }), .O ({new_AGEMA_signal_3598, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[67], key_s0[67]}), .I2 ({new_AGEMA_signal_2639, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 }), .I3 ({new_AGEMA_signal_2870, \KeyExpansionIns/tmp [3]}), .I4 ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }), .O ({new_AGEMA_signal_3600, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[68], key_s0[68]}), .I2 ({new_AGEMA_signal_2636, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 }), .I3 ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }), .I4 ({new_AGEMA_signal_2869, \KeyExpansionIns/tmp [4]}), .O ({new_AGEMA_signal_3602, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[69], key_s0[69]}), .I2 ({new_AGEMA_signal_2633, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 }), .I3 ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }), .I4 ({new_AGEMA_signal_2868, \KeyExpansionIns/tmp [5]}), .O ({new_AGEMA_signal_3604, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[70], key_s0[70]}), .I2 ({new_AGEMA_signal_2630, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 }), .I3 ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }), .I4 ({new_AGEMA_signal_2867, \KeyExpansionIns/tmp [6]}), .O ({new_AGEMA_signal_3606, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[71], key_s0[71]}), .I2 ({new_AGEMA_signal_2627, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 }), .I3 ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }), .I4 ({new_AGEMA_signal_2866, \KeyExpansionIns/tmp [7]}), .O ({new_AGEMA_signal_3608, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[72], key_s0[72]}), .I2 ({new_AGEMA_signal_2624, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 }), .I3 ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }), .I4 ({new_AGEMA_signal_2897, \KeyExpansionIns/tmp [8]}), .O ({new_AGEMA_signal_3610, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[73], key_s0[73]}), .I2 ({new_AGEMA_signal_2621, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 }), .I3 ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }), .I4 ({new_AGEMA_signal_2896, \KeyExpansionIns/tmp [9]}), .O ({new_AGEMA_signal_3612, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[74], key_s0[74]}), .I2 ({new_AGEMA_signal_2618, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 }), .I3 ({new_AGEMA_signal_2895, \KeyExpansionIns/tmp [10]}), .I4 ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }), .O ({new_AGEMA_signal_3614, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[75], key_s0[75]}), .I2 ({new_AGEMA_signal_2615, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 }), .I3 ({new_AGEMA_signal_2894, \KeyExpansionIns/tmp [11]}), .I4 ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }), .O ({new_AGEMA_signal_3616, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[76], key_s0[76]}), .I2 ({new_AGEMA_signal_2612, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 }), .I3 ({new_AGEMA_signal_2893, \KeyExpansionIns/tmp [12]}), .I4 ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }), .O ({new_AGEMA_signal_3618, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[77], key_s0[77]}), .I2 ({new_AGEMA_signal_2609, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 }), .I3 ({new_AGEMA_signal_2892, \KeyExpansionIns/tmp [13]}), .I4 ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }), .O ({new_AGEMA_signal_3620, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[78], key_s0[78]}), .I2 ({new_AGEMA_signal_2606, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 }), .I3 ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }), .I4 ({new_AGEMA_signal_2891, \KeyExpansionIns/tmp [14]}), .O ({new_AGEMA_signal_3622, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[79], key_s0[79]}), .I2 ({new_AGEMA_signal_2603, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 }), .I3 ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }), .I4 ({new_AGEMA_signal_2890, \KeyExpansionIns/tmp [15]}), .O ({new_AGEMA_signal_3624, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[80], key_s0[80]}), .I2 ({new_AGEMA_signal_2600, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 }), .I3 ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }), .I4 ({new_AGEMA_signal_2889, \KeyExpansionIns/tmp [16]}), .O ({new_AGEMA_signal_3626, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[81], key_s0[81]}), .I2 ({new_AGEMA_signal_2597, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 }), .I3 ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }), .I4 ({new_AGEMA_signal_2888, \KeyExpansionIns/tmp [17]}), .O ({new_AGEMA_signal_3628, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[82], key_s0[82]}), .I2 ({new_AGEMA_signal_2594, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 }), .I3 ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }), .I4 ({new_AGEMA_signal_2887, \KeyExpansionIns/tmp [18]}), .O ({new_AGEMA_signal_3630, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[83], key_s0[83]}), .I2 ({new_AGEMA_signal_2591, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 }), .I3 ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }), .I4 ({new_AGEMA_signal_2886, \KeyExpansionIns/tmp [19]}), .O ({new_AGEMA_signal_3632, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[84], key_s0[84]}), .I2 ({new_AGEMA_signal_2588, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 }), .I3 ({new_AGEMA_signal_2885, \KeyExpansionIns/tmp [20]}), .I4 ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }), .O ({new_AGEMA_signal_3634, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[85], key_s0[85]}), .I2 ({new_AGEMA_signal_2585, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 }), .I3 ({new_AGEMA_signal_2884, \KeyExpansionIns/tmp [21]}), .I4 ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }), .O ({new_AGEMA_signal_3636, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[86], key_s0[86]}), .I2 ({new_AGEMA_signal_2582, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 }), .I3 ({new_AGEMA_signal_2883, \KeyExpansionIns/tmp [22]}), .I4 ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }), .O ({new_AGEMA_signal_3638, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hD88D8DD8 ) , .MASK ( 5'b00001 ), .INIT2 ( 32'hD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({key_s1[87], key_s0[87]}), .I2 ({new_AGEMA_signal_2579, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 }), .I3 ({new_AGEMA_signal_2882, \KeyExpansionIns/tmp [23]}), .I4 ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }), .O ({new_AGEMA_signal_3640, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[88], key_s0[88]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2576, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 }), .I3 ({new_AGEMA_signal_3538, \KeyExpansionOutput<24>_bdd4 }), .O ({new_AGEMA_signal_3795, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[89], key_s0[89]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2573, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 }), .I3 ({new_AGEMA_signal_3544, \KeyExpansionOutput<25>_bdd4 }), .O ({new_AGEMA_signal_3797, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state }) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hB8 ) , .MASK ( 3'b010 ), .INIT2 ( 8'hB8 ) ) \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[90], key_s0[90]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_3751, KeyExpansionOutput[90]}), .O ({new_AGEMA_signal_3799, \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[91], key_s0[91]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2567, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 }), .I3 ({new_AGEMA_signal_3539, \KeyExpansionOutput<27>_bdd4 }), .O ({new_AGEMA_signal_3801, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[92], key_s0[92]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2564, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 }), .I3 ({new_AGEMA_signal_3542, \KeyExpansionOutput<28>_bdd4 }), .O ({new_AGEMA_signal_3803, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[93], key_s0[93]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2561, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 }), .I3 ({new_AGEMA_signal_3543, \KeyExpansionOutput<29>_bdd4 }), .O ({new_AGEMA_signal_3805, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[94], key_s0[94]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2558, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 }), .I3 ({new_AGEMA_signal_3541, \KeyExpansionOutput<30>_bdd4 }), .O ({new_AGEMA_signal_3807, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[95], key_s0[95]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2555, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 }), .I3 ({new_AGEMA_signal_3540, \KeyExpansionOutput<31>_bdd4 }), .O ({new_AGEMA_signal_3809, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2873, \KeyExpansionIns/tmp [0]}), .I2 ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }), .I3 ({key_s1[96], key_s0[96]}), .O ({new_AGEMA_signal_3642, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2872, \KeyExpansionIns/tmp [1]}), .I2 ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }), .I3 ({key_s1[97], key_s0[97]}), .O ({new_AGEMA_signal_3644, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2871, \KeyExpansionIns/tmp [2]}), .I2 ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }), .I3 ({key_s1[98], key_s0[98]}), .O ({new_AGEMA_signal_3646, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2870, \KeyExpansionIns/tmp [3]}), .I2 ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }), .I3 ({key_s1[99], key_s0[99]}), .O ({new_AGEMA_signal_3648, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }), .I2 ({new_AGEMA_signal_2869, \KeyExpansionIns/tmp [4]}), .I3 ({key_s1[100], key_s0[100]}), .O ({new_AGEMA_signal_3650, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }), .I2 ({new_AGEMA_signal_2868, \KeyExpansionIns/tmp [5]}), .I3 ({key_s1[101], key_s0[101]}), .O ({new_AGEMA_signal_3652, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }), .I2 ({new_AGEMA_signal_2867, \KeyExpansionIns/tmp [6]}), .I3 ({key_s1[102], key_s0[102]}), .O ({new_AGEMA_signal_3654, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }), .I2 ({new_AGEMA_signal_2866, \KeyExpansionIns/tmp [7]}), .I3 ({key_s1[103], key_s0[103]}), .O ({new_AGEMA_signal_3656, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }), .I2 ({new_AGEMA_signal_2897, \KeyExpansionIns/tmp [8]}), .I3 ({key_s1[104], key_s0[104]}), .O ({new_AGEMA_signal_3658, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }), .I2 ({new_AGEMA_signal_2896, \KeyExpansionIns/tmp [9]}), .I3 ({key_s1[105], key_s0[105]}), .O ({new_AGEMA_signal_3660, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2895, \KeyExpansionIns/tmp [10]}), .I2 ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }), .I3 ({key_s1[106], key_s0[106]}), .O ({new_AGEMA_signal_3662, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2894, \KeyExpansionIns/tmp [11]}), .I2 ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }), .I3 ({key_s1[107], key_s0[107]}), .O ({new_AGEMA_signal_3664, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2893, \KeyExpansionIns/tmp [12]}), .I2 ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }), .I3 ({key_s1[108], key_s0[108]}), .O ({new_AGEMA_signal_3666, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2892, \KeyExpansionIns/tmp [13]}), .I2 ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }), .I3 ({key_s1[109], key_s0[109]}), .O ({new_AGEMA_signal_3668, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }), .I2 ({new_AGEMA_signal_2891, \KeyExpansionIns/tmp [14]}), .I3 ({key_s1[110], key_s0[110]}), .O ({new_AGEMA_signal_3670, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }), .I2 ({new_AGEMA_signal_2890, \KeyExpansionIns/tmp [15]}), .I3 ({key_s1[111], key_s0[111]}), .O ({new_AGEMA_signal_3672, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }), .I2 ({new_AGEMA_signal_2889, \KeyExpansionIns/tmp [16]}), .I3 ({key_s1[112], key_s0[112]}), .O ({new_AGEMA_signal_3674, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }), .I2 ({new_AGEMA_signal_2888, \KeyExpansionIns/tmp [17]}), .I3 ({key_s1[113], key_s0[113]}), .O ({new_AGEMA_signal_3676, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }), .I2 ({new_AGEMA_signal_2887, \KeyExpansionIns/tmp [18]}), .I3 ({key_s1[114], key_s0[114]}), .O ({new_AGEMA_signal_3678, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }), .I2 ({new_AGEMA_signal_2886, \KeyExpansionIns/tmp [19]}), .I3 ({key_s1[115], key_s0[115]}), .O ({new_AGEMA_signal_3680, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2885, \KeyExpansionIns/tmp [20]}), .I2 ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }), .I3 ({key_s1[116], key_s0[116]}), .O ({new_AGEMA_signal_3682, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2884, \KeyExpansionIns/tmp [21]}), .I2 ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }), .I3 ({key_s1[117], key_s0[117]}), .O ({new_AGEMA_signal_3684, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2883, \KeyExpansionIns/tmp [22]}), .I2 ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }), .I3 ({key_s1[118], key_s0[118]}), .O ({new_AGEMA_signal_3686, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'hBE14 ) , .MASK ( 4'b0001 ), .INIT2 ( 16'hBE14 ) ) \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2882, \KeyExpansionIns/tmp [23]}), .I2 ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }), .I3 ({key_s1[119], key_s0[119]}), .O ({new_AGEMA_signal_3688, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[0], key_s0[0]}), .I2 ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }), .I3 ({new_AGEMA_signal_2648, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 }), .I4 ({new_AGEMA_signal_2873, \KeyExpansionIns/tmp [0]}), .I5 ({new_AGEMA_signal_2842, N01}), .O ({new_AGEMA_signal_3690, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[1], key_s0[1]}), .I2 ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }), .I3 ({new_AGEMA_signal_2645, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 }), .I4 ({new_AGEMA_signal_2872, \KeyExpansionIns/tmp [1]}), .I5 ({new_AGEMA_signal_2843, N2}), .O ({new_AGEMA_signal_3692, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[2], key_s0[2]}), .I2 ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }), .I3 ({new_AGEMA_signal_2642, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 }), .I4 ({new_AGEMA_signal_2871, \KeyExpansionIns/tmp [2]}), .I5 ({new_AGEMA_signal_2844, N4}), .O ({new_AGEMA_signal_3694, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[3], key_s0[3]}), .I2 ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }), .I3 ({new_AGEMA_signal_2639, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 }), .I4 ({new_AGEMA_signal_2870, \KeyExpansionIns/tmp [3]}), .I5 ({new_AGEMA_signal_2845, N6}), .O ({new_AGEMA_signal_3696, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[4], key_s0[4]}), .I2 ({new_AGEMA_signal_2636, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 }), .I3 ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }), .I4 ({new_AGEMA_signal_2869, \KeyExpansionIns/tmp [4]}), .I5 ({new_AGEMA_signal_2846, N8}), .O ({new_AGEMA_signal_3698, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[5], key_s0[5]}), .I2 ({new_AGEMA_signal_2633, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 }), .I3 ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }), .I4 ({new_AGEMA_signal_2868, \KeyExpansionIns/tmp [5]}), .I5 ({new_AGEMA_signal_2847, N10}), .O ({new_AGEMA_signal_3700, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[6], key_s0[6]}), .I2 ({new_AGEMA_signal_2630, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 }), .I3 ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }), .I4 ({new_AGEMA_signal_2867, \KeyExpansionIns/tmp [6]}), .I5 ({new_AGEMA_signal_2848, N12}), .O ({new_AGEMA_signal_3702, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[7], key_s0[7]}), .I2 ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }), .I3 ({new_AGEMA_signal_2627, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 }), .I4 ({new_AGEMA_signal_2866, \KeyExpansionIns/tmp [7]}), .I5 ({new_AGEMA_signal_2849, N14}), .O ({new_AGEMA_signal_3704, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[8], key_s0[8]}), .I2 ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }), .I3 ({new_AGEMA_signal_2624, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 }), .I4 ({new_AGEMA_signal_2897, \KeyExpansionIns/tmp [8]}), .I5 ({new_AGEMA_signal_2850, N16}), .O ({new_AGEMA_signal_3706, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[9], key_s0[9]}), .I2 ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }), .I3 ({new_AGEMA_signal_2621, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 }), .I4 ({new_AGEMA_signal_2896, \KeyExpansionIns/tmp [9]}), .I5 ({new_AGEMA_signal_2851, N18}), .O ({new_AGEMA_signal_3708, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[10], key_s0[10]}), .I2 ({new_AGEMA_signal_2618, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 }), .I3 ({new_AGEMA_signal_2714, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_471 }), .I4 ({new_AGEMA_signal_2895, \KeyExpansionIns/tmp [10]}), .I5 ({new_AGEMA_signal_2852, N20}), .O ({new_AGEMA_signal_3710, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[11], key_s0[11]}), .I2 ({new_AGEMA_signal_2615, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 }), .I3 ({new_AGEMA_signal_2711, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_470 }), .I4 ({new_AGEMA_signal_2894, \KeyExpansionIns/tmp [11]}), .I5 ({new_AGEMA_signal_2853, N22}), .O ({new_AGEMA_signal_3712, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[12], key_s0[12]}), .I2 ({new_AGEMA_signal_2612, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 }), .I3 ({new_AGEMA_signal_2708, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_469 }), .I4 ({new_AGEMA_signal_2893, \KeyExpansionIns/tmp [12]}), .I5 ({new_AGEMA_signal_2854, N24}), .O ({new_AGEMA_signal_3714, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[13], key_s0[13]}), .I2 ({new_AGEMA_signal_2609, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 }), .I3 ({new_AGEMA_signal_2705, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_468 }), .I4 ({new_AGEMA_signal_2892, \KeyExpansionIns/tmp [13]}), .I5 ({new_AGEMA_signal_2855, N26}), .O ({new_AGEMA_signal_3716, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[14], key_s0[14]}), .I2 ({new_AGEMA_signal_2606, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 }), .I3 ({new_AGEMA_signal_2702, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_467 }), .I4 ({new_AGEMA_signal_2891, \KeyExpansionIns/tmp [14]}), .I5 ({new_AGEMA_signal_2856, N28}), .O ({new_AGEMA_signal_3718, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[15], key_s0[15]}), .I2 ({new_AGEMA_signal_2603, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 }), .I3 ({new_AGEMA_signal_2699, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_466 }), .I4 ({new_AGEMA_signal_2890, \KeyExpansionIns/tmp [15]}), .I5 ({new_AGEMA_signal_2857, N30}), .O ({new_AGEMA_signal_3720, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[16], key_s0[16]}), .I2 ({new_AGEMA_signal_2600, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 }), .I3 ({new_AGEMA_signal_2696, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_465 }), .I4 ({new_AGEMA_signal_2889, \KeyExpansionIns/tmp [16]}), .I5 ({new_AGEMA_signal_2858, N32}), .O ({new_AGEMA_signal_3722, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[17], key_s0[17]}), .I2 ({new_AGEMA_signal_2597, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 }), .I3 ({new_AGEMA_signal_2693, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_464 }), .I4 ({new_AGEMA_signal_2888, \KeyExpansionIns/tmp [17]}), .I5 ({new_AGEMA_signal_2859, N34}), .O ({new_AGEMA_signal_3724, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[18], key_s0[18]}), .I2 ({new_AGEMA_signal_2594, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 }), .I3 ({new_AGEMA_signal_2690, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_463 }), .I4 ({new_AGEMA_signal_2887, \KeyExpansionIns/tmp [18]}), .I5 ({new_AGEMA_signal_2860, N36}), .O ({new_AGEMA_signal_3726, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[19], key_s0[19]}), .I2 ({new_AGEMA_signal_2591, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 }), .I3 ({new_AGEMA_signal_2687, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_462 }), .I4 ({new_AGEMA_signal_2886, \KeyExpansionIns/tmp [19]}), .I5 ({new_AGEMA_signal_2861, N38}), .O ({new_AGEMA_signal_3728, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[20], key_s0[20]}), .I2 ({new_AGEMA_signal_2588, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 }), .I3 ({new_AGEMA_signal_2684, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_461 }), .I4 ({new_AGEMA_signal_2885, \KeyExpansionIns/tmp [20]}), .I5 ({new_AGEMA_signal_2862, N40}), .O ({new_AGEMA_signal_3730, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[21], key_s0[21]}), .I2 ({new_AGEMA_signal_2585, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 }), .I3 ({new_AGEMA_signal_2681, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_460 }), .I4 ({new_AGEMA_signal_2884, \KeyExpansionIns/tmp [21]}), .I5 ({new_AGEMA_signal_2863, N42}), .O ({new_AGEMA_signal_3732, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[22], key_s0[22]}), .I2 ({new_AGEMA_signal_2582, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 }), .I3 ({new_AGEMA_signal_2678, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_459 }), .I4 ({new_AGEMA_signal_2883, \KeyExpansionIns/tmp [22]}), .I5 ({new_AGEMA_signal_2864, N44}), .O ({new_AGEMA_signal_3734, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8DD8D88DD88D8DD8 ) , .MASK ( 6'b000001 ), .INIT2 ( 64'h8DD8D88DD88D8DD8 ) ) \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({key_s1[23], key_s0[23]}), .I2 ({new_AGEMA_signal_2579, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 }), .I3 ({new_AGEMA_signal_2675, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_458 }), .I4 ({new_AGEMA_signal_2882, \KeyExpansionIns/tmp [23]}), .I5 ({new_AGEMA_signal_2865, N46}), .O ({new_AGEMA_signal_3736, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2480, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_393 }), .I2 ({new_AGEMA_signal_2881, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [0]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, N48}), .I5 ({key_s1[120], key_s0[120]}), .O ({new_AGEMA_signal_3738, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2477, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_392 }), .I2 ({new_AGEMA_signal_2880, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [1]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, N50}), .I5 ({key_s1[121], key_s0[121]}), .O ({new_AGEMA_signal_3740, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2471, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_390 }), .I2 ({new_AGEMA_signal_2878, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [3]}), .I3 ({1'b0, \RoundCounterIns/count [2]}), .I4 ({1'b0, N52}), .I5 ({key_s1[123], key_s0[123]}), .O ({new_AGEMA_signal_3742, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2468, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_389 }), .I2 ({new_AGEMA_signal_2877, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [4]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, N54}), .I5 ({key_s1[124], key_s0[124]}), .O ({new_AGEMA_signal_3744, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2465, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_388 }), .I2 ({new_AGEMA_signal_2876, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [5]}), .I3 ({1'b0, \RoundCounterIns/count [1]}), .I4 ({1'b0, N56}), .I5 ({key_s1[125], key_s0[125]}), .O ({new_AGEMA_signal_3746, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2462, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_387 }), .I2 ({new_AGEMA_signal_2875, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [6]}), .I3 ({1'b0, \RoundCounterIns/count [3]}), .I4 ({1'b0, N58}), .I5 ({key_s1[126], key_s0[126]}), .O ({new_AGEMA_signal_3748, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2459, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_386 }), .I2 ({new_AGEMA_signal_2874, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [7]}), .I3 ({1'b0, \RoundCounterIns/count [3]}), .I4 ({1'b0, N60}), .I5 ({key_s1[127], key_s0[127]}), .O ({new_AGEMA_signal_3750, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I2 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .I3 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3810, N62}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[0], plaintext_s0[0]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3442, ShiftRowsInput[32]}), .I4 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I5 ({new_AGEMA_signal_3810, N62}), .O ({new_AGEMA_signal_3943, \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I1 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .I2 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .I3 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .I4 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .O ({new_AGEMA_signal_3811, N64}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[1], plaintext_s0[1]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I4 ({new_AGEMA_signal_3755, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3811, N64}), .O ({new_AGEMA_signal_3945, \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .I1 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .I2 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .I3 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .O ({new_AGEMA_signal_3812, N66}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[2], plaintext_s0[2]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3444, ShiftRowsInput[34]}), .I4 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I5 ({new_AGEMA_signal_3812, N66}), .O ({new_AGEMA_signal_3947, \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .I1 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I2 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .I3 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .I4 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3813, N68}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[3], plaintext_s0[3]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3445, ShiftRowsInput[35]}), .I4 ({new_AGEMA_signal_3756, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3813, N68}), .O ({new_AGEMA_signal_3949, \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I1 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I2 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .I3 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .I4 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3814, N70}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[4], plaintext_s0[4]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I4 ({new_AGEMA_signal_3760, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3814, N70}), .O ({new_AGEMA_signal_3951, \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I1 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I2 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .I3 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .O ({new_AGEMA_signal_3815, N72}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[5], plaintext_s0[5]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .I4 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I5 ({new_AGEMA_signal_3815, N72}), .O ({new_AGEMA_signal_3953, \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .I1 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I2 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .I3 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .O ({new_AGEMA_signal_3816, N74}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[6], plaintext_s0[6]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I4 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I5 ({new_AGEMA_signal_3816, N74}), .O ({new_AGEMA_signal_3955, \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I1 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I2 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .I3 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3817, N76}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[7], plaintext_s0[7]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3817, N76}), .O ({new_AGEMA_signal_3957, \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3442, ShiftRowsInput[32]}), .I1 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I2 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I3 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .O ({new_AGEMA_signal_3818, N78}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[8], plaintext_s0[8]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3818, N78}), .O ({new_AGEMA_signal_3959, \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I1 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .I2 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I3 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I4 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .O ({new_AGEMA_signal_3819, N80}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[9], plaintext_s0[9]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I4 ({new_AGEMA_signal_3755, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3819, N80}), .O ({new_AGEMA_signal_3961, \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3444, ShiftRowsInput[34]}), .I1 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .I2 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I3 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .O ({new_AGEMA_signal_3820, N82}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[10], plaintext_s0[10]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .I4 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I5 ({new_AGEMA_signal_3820, N82}), .O ({new_AGEMA_signal_3963, \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3445, ShiftRowsInput[35]}), .I1 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .I2 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I3 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I4 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .O ({new_AGEMA_signal_3821, N84}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[11], plaintext_s0[11]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .I4 ({new_AGEMA_signal_3756, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3821, N84}), .O ({new_AGEMA_signal_3965, \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I1 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .I2 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I3 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I4 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .O ({new_AGEMA_signal_3822, N86}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[12], plaintext_s0[12]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I4 ({new_AGEMA_signal_3760, \MixColumnsIns/GenMixColumns[3].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3822, N86}), .O ({new_AGEMA_signal_3967, \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .I1 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I2 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I3 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .O ({new_AGEMA_signal_3823, N88}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[13], plaintext_s0[13]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I4 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I5 ({new_AGEMA_signal_3823, N88}), .O ({new_AGEMA_signal_3969, \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .I1 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I2 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I3 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .O ({new_AGEMA_signal_3824, N90}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[14], plaintext_s0[14]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I4 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I5 ({new_AGEMA_signal_3824, N90}), .O ({new_AGEMA_signal_3971, \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I2 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I3 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3825, N92}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[15], plaintext_s0[15]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3825, N92}), .O ({new_AGEMA_signal_3973, \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3442, ShiftRowsInput[32]}), .I1 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I2 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I3 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .O ({new_AGEMA_signal_3826, N94}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[16], plaintext_s0[16]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3826, N94}), .O ({new_AGEMA_signal_3975, \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I1 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I2 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .O ({new_AGEMA_signal_3827, N96}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[17], plaintext_s0[17]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .I4 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I5 ({new_AGEMA_signal_3827, N96}), .O ({new_AGEMA_signal_3977, \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3444, ShiftRowsInput[34]}), .I1 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .I2 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .I3 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .O ({new_AGEMA_signal_3828, N98}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[18], plaintext_s0[18]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .I4 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I5 ({new_AGEMA_signal_3828, N98}), .O ({new_AGEMA_signal_3979, \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .I1 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .I2 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .O ({new_AGEMA_signal_3829, N100}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[19], plaintext_s0[19]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3445, ShiftRowsInput[35]}), .I4 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I5 ({new_AGEMA_signal_3829, N100}), .O ({new_AGEMA_signal_3981, \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .I1 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I2 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .O ({new_AGEMA_signal_3830, N102}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[20], plaintext_s0[20]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I4 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I5 ({new_AGEMA_signal_3830, N102}), .O ({new_AGEMA_signal_3983, \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I1 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I2 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .I3 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .O ({new_AGEMA_signal_3831, N104}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[21], plaintext_s0[21]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I4 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I5 ({new_AGEMA_signal_3831, N104}), .O ({new_AGEMA_signal_3985, \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I1 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I2 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I3 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .O ({new_AGEMA_signal_3832, N106}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[22], plaintext_s0[22]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I4 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I5 ({new_AGEMA_signal_3832, N106}), .O ({new_AGEMA_signal_3987, \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I1 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I2 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I3 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3833, N108}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[23], plaintext_s0[23]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I5 ({new_AGEMA_signal_3833, N108}), .O ({new_AGEMA_signal_3989, \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3442, ShiftRowsInput[32]}), .I1 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I2 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I3 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3834, N110}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[24], plaintext_s0[24]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3482, ShiftRowsInput[72]}), .I4 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .I5 ({new_AGEMA_signal_3834, N110}), .O ({new_AGEMA_signal_3991, \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3522, ShiftRowsInput[112]}), .I1 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .I2 ({new_AGEMA_signal_3443, ShiftRowsInput[33]}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3434, ShiftRowsInput[24]}), .I5 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3835, N112}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[25], plaintext_s0[25]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3483, ShiftRowsInput[73]}), .I4 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .I5 ({new_AGEMA_signal_3835, N112}), .O ({new_AGEMA_signal_3993, \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3484, ShiftRowsInput[74]}), .I1 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .I2 ({new_AGEMA_signal_3523, ShiftRowsInput[113]}), .I3 ({new_AGEMA_signal_3444, ShiftRowsInput[34]}), .O ({new_AGEMA_signal_3836, N114}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[26], plaintext_s0[26]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .I4 ({new_AGEMA_signal_3435, ShiftRowsInput[25]}), .I5 ({new_AGEMA_signal_3836, N114}), .O ({new_AGEMA_signal_3995, \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I1 ({new_AGEMA_signal_3485, ShiftRowsInput[75]}), .I2 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .I3 ({new_AGEMA_signal_3436, ShiftRowsInput[26]}), .I4 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I5 ({new_AGEMA_signal_3524, ShiftRowsInput[114]}), .O ({new_AGEMA_signal_3837, N116}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[27], plaintext_s0[27]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3445, ShiftRowsInput[35]}), .I4 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .I5 ({new_AGEMA_signal_3837, N116}), .O ({new_AGEMA_signal_3997, \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3486, ShiftRowsInput[76]}), .I1 ({new_AGEMA_signal_3525, ShiftRowsInput[115]}), .I2 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I3 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I4 ({new_AGEMA_signal_3437, ShiftRowsInput[27]}), .I5 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .O ({new_AGEMA_signal_3838, N118}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[28], plaintext_s0[28]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3446, ShiftRowsInput[36]}), .I4 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .I5 ({new_AGEMA_signal_3838, N118}), .O ({new_AGEMA_signal_3999, \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3526, ShiftRowsInput[116]}), .I1 ({new_AGEMA_signal_3487, ShiftRowsInput[77]}), .I2 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I3 ({new_AGEMA_signal_3447, ShiftRowsInput[37]}), .O ({new_AGEMA_signal_3839, N120}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[29], plaintext_s0[29]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .I4 ({new_AGEMA_signal_3438, ShiftRowsInput[28]}), .I5 ({new_AGEMA_signal_3839, N120}), .O ({new_AGEMA_signal_4001, \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3448, ShiftRowsInput[38]}), .I1 ({new_AGEMA_signal_3527, ShiftRowsInput[117]}), .I2 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I3 ({new_AGEMA_signal_3439, ShiftRowsInput[29]}), .O ({new_AGEMA_signal_3840, N122}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[30], plaintext_s0[30]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3488, ShiftRowsInput[78]}), .I4 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .I5 ({new_AGEMA_signal_3840, N122}), .O ({new_AGEMA_signal_4003, \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3528, ShiftRowsInput[118]}), .I1 ({new_AGEMA_signal_3449, ShiftRowsInput[39]}), .I2 ({new_AGEMA_signal_3529, ShiftRowsInput[119]}), .I3 ({new_AGEMA_signal_3440, ShiftRowsInput[30]}), .O ({new_AGEMA_signal_3841, N124}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[31], plaintext_s0[31]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3489, ShiftRowsInput[79]}), .I4 ({new_AGEMA_signal_3441, ShiftRowsInput[31]}), .I5 ({new_AGEMA_signal_3841, N124}), .O ({new_AGEMA_signal_4005, \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .I1 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I2 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I3 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .O ({new_AGEMA_signal_3842, N126}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[32], plaintext_s0[32]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3474, ShiftRowsInput[64]}), .I4 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I5 ({new_AGEMA_signal_3842, N126}), .O ({new_AGEMA_signal_4007, \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I1 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I2 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I3 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I4 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .O ({new_AGEMA_signal_3843, N128}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[33], plaintext_s0[33]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I4 ({new_AGEMA_signal_3757, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3843, N128}), .O ({new_AGEMA_signal_4009, \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I1 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I2 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .I3 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .O ({new_AGEMA_signal_3844, N130}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[34], plaintext_s0[34]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3476, ShiftRowsInput[66]}), .I4 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I5 ({new_AGEMA_signal_3844, N130}), .O ({new_AGEMA_signal_4011, \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I1 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I2 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I3 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I4 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .O ({new_AGEMA_signal_3845, N132}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[35], plaintext_s0[35]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3477, ShiftRowsInput[67]}), .I4 ({new_AGEMA_signal_3758, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3845, N132}), .O ({new_AGEMA_signal_4013, \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I1 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I2 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .I3 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I4 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .O ({new_AGEMA_signal_3846, N134}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[36], plaintext_s0[36]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I4 ({new_AGEMA_signal_3759, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3846, N134}), .O ({new_AGEMA_signal_4015, \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I1 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I2 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .I3 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .O ({new_AGEMA_signal_3847, N136}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[37], plaintext_s0[37]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .I4 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I5 ({new_AGEMA_signal_3847, N136}), .O ({new_AGEMA_signal_4017, \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .I1 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I2 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I3 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .O ({new_AGEMA_signal_3848, N138}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[38], plaintext_s0[38]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I4 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I5 ({new_AGEMA_signal_3848, N138}), .O ({new_AGEMA_signal_4019, \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I1 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I2 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I3 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3849, N140}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[39], plaintext_s0[39]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I4 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I5 ({new_AGEMA_signal_3849, N140}), .O ({new_AGEMA_signal_4021, \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3474, ShiftRowsInput[64]}), .I1 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I2 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I3 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .O ({new_AGEMA_signal_3850, N142}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[40], plaintext_s0[40]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .I4 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I5 ({new_AGEMA_signal_3850, N142}), .O ({new_AGEMA_signal_4023, \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I1 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I2 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .O ({new_AGEMA_signal_3851, N144}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[41], plaintext_s0[41]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I4 ({new_AGEMA_signal_3757, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3851, N144}), .O ({new_AGEMA_signal_4025, \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I1 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I2 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .I3 ({new_AGEMA_signal_3476, ShiftRowsInput[66]}), .O ({new_AGEMA_signal_3852, N146}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[42], plaintext_s0[42]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .I4 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I5 ({new_AGEMA_signal_3852, N146}), .O ({new_AGEMA_signal_4027, \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3477, ShiftRowsInput[67]}), .I1 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I2 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .O ({new_AGEMA_signal_3853, N148}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[43], plaintext_s0[43]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .I4 ({new_AGEMA_signal_3758, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3853, N148}), .O ({new_AGEMA_signal_4029, \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I1 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I2 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .O ({new_AGEMA_signal_3854, N150}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[44], plaintext_s0[44]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .I4 ({new_AGEMA_signal_3759, \MixColumnsIns/GenMixColumns[2].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3854, N150}), .O ({new_AGEMA_signal_4031, \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .I1 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .I2 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I3 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .O ({new_AGEMA_signal_3855, N152}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[45], plaintext_s0[45]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .I4 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I5 ({new_AGEMA_signal_3855, N152}), .O ({new_AGEMA_signal_4033, \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .I1 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I2 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .I3 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .O ({new_AGEMA_signal_3856, N154}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[46], plaintext_s0[46]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I4 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I5 ({new_AGEMA_signal_3856, N154}), .O ({new_AGEMA_signal_4035, \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I1 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I2 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I3 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3857, N156}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[47], plaintext_s0[47]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I5 ({new_AGEMA_signal_3857, N156}), .O ({new_AGEMA_signal_4037, \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3474, ShiftRowsInput[64]}), .I1 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .I2 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I3 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3858, N158}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[48], plaintext_s0[48]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I4 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .I5 ({new_AGEMA_signal_3858, N158}), .O ({new_AGEMA_signal_4039, \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I1 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I2 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .I3 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .I4 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I5 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .O ({new_AGEMA_signal_3859, N160}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[49], plaintext_s0[49]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I4 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .I5 ({new_AGEMA_signal_3859, N160}), .O ({new_AGEMA_signal_4041, \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3476, ShiftRowsInput[66]}), .I1 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .I2 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I3 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .O ({new_AGEMA_signal_3860, N162}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[50], plaintext_s0[50]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I4 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .I5 ({new_AGEMA_signal_3860, N162}), .O ({new_AGEMA_signal_4043, \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .I1 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .I2 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .I5 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3861, N164}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[51], plaintext_s0[51]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3477, ShiftRowsInput[67]}), .I4 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I5 ({new_AGEMA_signal_3861, N164}), .O ({new_AGEMA_signal_4045, \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .I1 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .I2 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I3 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I4 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I5 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3862, N166}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[52], plaintext_s0[52]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I4 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .I5 ({new_AGEMA_signal_3862, N166}), .O ({new_AGEMA_signal_4047, \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I1 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .I2 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .I3 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .O ({new_AGEMA_signal_3863, N168}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[53], plaintext_s0[53]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .I4 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .I5 ({new_AGEMA_signal_3863, N168}), .O ({new_AGEMA_signal_4049, \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I1 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .I2 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I3 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .O ({new_AGEMA_signal_3864, N170}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[54], plaintext_s0[54]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I4 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .I5 ({new_AGEMA_signal_3864, N170}), .O ({new_AGEMA_signal_4051, \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I1 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I2 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I3 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .O ({new_AGEMA_signal_3865, N172}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[55], plaintext_s0[55]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I4 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .I5 ({new_AGEMA_signal_3865, N172}), .O ({new_AGEMA_signal_4053, \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3474, ShiftRowsInput[64]}), .I1 ({new_AGEMA_signal_3514, ShiftRowsInput[104]}), .I2 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .I3 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3866, N174}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[56], plaintext_s0[56]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I4 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I5 ({new_AGEMA_signal_3866, N174}), .O ({new_AGEMA_signal_4055, \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3466, ShiftRowsInput[56]}), .I1 ({new_AGEMA_signal_3515, ShiftRowsInput[105]}), .I2 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I3 ({new_AGEMA_signal_3426, ShiftRowsInput[16]}), .I4 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .I5 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3867, N176}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[57], plaintext_s0[57]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I4 ({new_AGEMA_signal_3475, ShiftRowsInput[65]}), .I5 ({new_AGEMA_signal_3867, N176}), .O ({new_AGEMA_signal_4057, \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3476, ShiftRowsInput[66]}), .I1 ({new_AGEMA_signal_3516, ShiftRowsInput[106]}), .I2 ({new_AGEMA_signal_3427, ShiftRowsInput[17]}), .I3 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .O ({new_AGEMA_signal_3868, N178}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[58], plaintext_s0[58]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I4 ({new_AGEMA_signal_3467, ShiftRowsInput[57]}), .I5 ({new_AGEMA_signal_3868, N178}), .O ({new_AGEMA_signal_4059, \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3517, ShiftRowsInput[107]}), .I1 ({new_AGEMA_signal_3468, ShiftRowsInput[58]}), .I2 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I3 ({new_AGEMA_signal_3428, ShiftRowsInput[18]}), .I4 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I5 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3869, N180}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[59], plaintext_s0[59]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3477, ShiftRowsInput[67]}), .I4 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I5 ({new_AGEMA_signal_3869, N180}), .O ({new_AGEMA_signal_4061, \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3518, ShiftRowsInput[108]}), .I1 ({new_AGEMA_signal_3469, ShiftRowsInput[59]}), .I2 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I3 ({new_AGEMA_signal_3429, ShiftRowsInput[19]}), .I4 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .I5 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3870, N182}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[60], plaintext_s0[60]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I4 ({new_AGEMA_signal_3478, ShiftRowsInput[68]}), .I5 ({new_AGEMA_signal_3870, N182}), .O ({new_AGEMA_signal_4063, \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3479, ShiftRowsInput[69]}), .I1 ({new_AGEMA_signal_3519, ShiftRowsInput[109]}), .I2 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .I3 ({new_AGEMA_signal_3430, ShiftRowsInput[20]}), .O ({new_AGEMA_signal_3871, N184}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[61], plaintext_s0[61]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I4 ({new_AGEMA_signal_3470, ShiftRowsInput[60]}), .I5 ({new_AGEMA_signal_3871, N184}), .O ({new_AGEMA_signal_4065, \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3480, ShiftRowsInput[70]}), .I1 ({new_AGEMA_signal_3520, ShiftRowsInput[110]}), .I2 ({new_AGEMA_signal_3431, ShiftRowsInput[21]}), .I3 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .O ({new_AGEMA_signal_3872, N186}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[62], plaintext_s0[62]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I4 ({new_AGEMA_signal_3471, ShiftRowsInput[61]}), .I5 ({new_AGEMA_signal_3872, N186}), .O ({new_AGEMA_signal_4067, \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3481, ShiftRowsInput[71]}), .I1 ({new_AGEMA_signal_3521, ShiftRowsInput[111]}), .I2 ({new_AGEMA_signal_3432, ShiftRowsInput[22]}), .I3 ({new_AGEMA_signal_3433, ShiftRowsInput[23]}), .O ({new_AGEMA_signal_3873, N188}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[63], plaintext_s0[63]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3472, ShiftRowsInput[62]}), .I4 ({new_AGEMA_signal_3473, ShiftRowsInput[63]}), .I5 ({new_AGEMA_signal_3873, N188}), .O ({new_AGEMA_signal_4069, \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I1 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I2 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I3 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .O ({new_AGEMA_signal_3874, N190}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[64], plaintext_s0[64]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3506, ShiftRowsInput[96]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3874, N190}), .O ({new_AGEMA_signal_4071, \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I1 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I2 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I3 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I4 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .O ({new_AGEMA_signal_3875, N192}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[65], plaintext_s0[65]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I4 ({new_AGEMA_signal_3761, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3875, N192}), .O ({new_AGEMA_signal_4073, \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I1 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I2 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I3 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .O ({new_AGEMA_signal_3876, N194}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[66], plaintext_s0[66]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3508, ShiftRowsInput[98]}), .I4 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I5 ({new_AGEMA_signal_3876, N194}), .O ({new_AGEMA_signal_4075, \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I1 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I2 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I3 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I4 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .O ({new_AGEMA_signal_3877, N196}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[67], plaintext_s0[67]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3509, ShiftRowsInput[99]}), .I4 ({new_AGEMA_signal_3762, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3877, N196}), .O ({new_AGEMA_signal_4077, \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I1 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I2 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I3 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I4 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .O ({new_AGEMA_signal_3878, N198}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[68], plaintext_s0[68]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I4 ({new_AGEMA_signal_3763, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3878, N198}), .O ({new_AGEMA_signal_4079, \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I1 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I2 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I3 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .O ({new_AGEMA_signal_3879, N200}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[69], plaintext_s0[69]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .I4 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I5 ({new_AGEMA_signal_3879, N200}), .O ({new_AGEMA_signal_4081, \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I1 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I2 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .I3 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .O ({new_AGEMA_signal_3880, N202}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[70], plaintext_s0[70]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .I4 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I5 ({new_AGEMA_signal_3880, N202}), .O ({new_AGEMA_signal_4083, \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I1 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I2 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I3 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .O ({new_AGEMA_signal_3881, N204}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[71], plaintext_s0[71]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3881, N204}), .O ({new_AGEMA_signal_4085, \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3506, ShiftRowsInput[96]}), .I1 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I2 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3882, N206}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[72], plaintext_s0[72]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I4 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .I5 ({new_AGEMA_signal_3882, N206}), .O ({new_AGEMA_signal_4087, \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I1 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I2 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .I3 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I4 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3883, N208}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[73], plaintext_s0[73]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .I4 ({new_AGEMA_signal_3761, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3883, N208}), .O ({new_AGEMA_signal_4089, \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I1 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I2 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I3 ({new_AGEMA_signal_3508, ShiftRowsInput[98]}), .O ({new_AGEMA_signal_3884, N210}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[74], plaintext_s0[74]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .I4 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .I5 ({new_AGEMA_signal_3884, N210}), .O ({new_AGEMA_signal_4091, \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3509, ShiftRowsInput[99]}), .I1 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I2 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I4 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .O ({new_AGEMA_signal_3885, N212}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[75], plaintext_s0[75]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .I4 ({new_AGEMA_signal_3762, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3885, N212}), .O ({new_AGEMA_signal_4093, \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I1 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I2 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I4 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .O ({new_AGEMA_signal_3886, N214}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[76], plaintext_s0[76]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .I4 ({new_AGEMA_signal_3763, \MixColumnsIns/GenMixColumns[1].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3886, N214}), .O ({new_AGEMA_signal_4095, \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I1 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I2 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .I3 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .O ({new_AGEMA_signal_3887, N216}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[77], plaintext_s0[77]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I4 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .I5 ({new_AGEMA_signal_3887, N216}), .O ({new_AGEMA_signal_4097, \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .I1 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .I2 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I3 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .O ({new_AGEMA_signal_3888, N218}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[78], plaintext_s0[78]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I4 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .I5 ({new_AGEMA_signal_3888, N218}), .O ({new_AGEMA_signal_4099, \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I2 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I3 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .O ({new_AGEMA_signal_3889, N220}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[79], plaintext_s0[79]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I4 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I5 ({new_AGEMA_signal_3889, N220}), .O ({new_AGEMA_signal_4101, \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I1 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I2 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I3 ({new_AGEMA_signal_3506, ShiftRowsInput[96]}), .O ({new_AGEMA_signal_3890, N222}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[80], plaintext_s0[80]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I4 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .I5 ({new_AGEMA_signal_3890, N222}), .O ({new_AGEMA_signal_4103, \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I1 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I2 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .I3 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I4 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I5 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3891, N224}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[81], plaintext_s0[81]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I4 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .I5 ({new_AGEMA_signal_3891, N224}), .O ({new_AGEMA_signal_4105, \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I1 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I2 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .I3 ({new_AGEMA_signal_3508, ShiftRowsInput[98]}), .O ({new_AGEMA_signal_3892, N226}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[82], plaintext_s0[82]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I4 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .I5 ({new_AGEMA_signal_3892, N226}), .O ({new_AGEMA_signal_4107, \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I1 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I2 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I3 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .I4 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .I5 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3893, N228}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[83], plaintext_s0[83]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3509, ShiftRowsInput[99]}), .I4 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I5 ({new_AGEMA_signal_3893, N228}), .O ({new_AGEMA_signal_4109, \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I1 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I2 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .I4 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .I5 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .O ({new_AGEMA_signal_3894, N230}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[84], plaintext_s0[84]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I4 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I5 ({new_AGEMA_signal_3894, N230}), .O ({new_AGEMA_signal_4111, \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .I1 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I2 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .I3 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .O ({new_AGEMA_signal_3895, N232}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[85], plaintext_s0[85]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I4 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I5 ({new_AGEMA_signal_3895, N232}), .O ({new_AGEMA_signal_4113, \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .I1 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I2 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .I3 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .O ({new_AGEMA_signal_3896, N234}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[86], plaintext_s0[86]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I4 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I5 ({new_AGEMA_signal_3896, N234}), .O ({new_AGEMA_signal_4115, \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I2 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3897, N236}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[87], plaintext_s0[87]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3897, N236}), .O ({new_AGEMA_signal_4117, \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3506, ShiftRowsInput[96]}), .I1 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I2 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I3 ({new_AGEMA_signal_3418, ShiftRowsInput[8]}), .O ({new_AGEMA_signal_3898, N238}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[88], plaintext_s0[88]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3898, N238}), .O ({new_AGEMA_signal_4119, \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3458, ShiftRowsInput[48]}), .I1 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I2 ({new_AGEMA_signal_3498, ShiftRowsInput[88]}), .I3 ({new_AGEMA_signal_3507, ShiftRowsInput[97]}), .I4 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I5 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .O ({new_AGEMA_signal_3899, N240}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[89], plaintext_s0[89]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I4 ({new_AGEMA_signal_3419, ShiftRowsInput[9]}), .I5 ({new_AGEMA_signal_3899, N240}), .O ({new_AGEMA_signal_4121, \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I1 ({new_AGEMA_signal_3459, ShiftRowsInput[49]}), .I2 ({new_AGEMA_signal_3420, ShiftRowsInput[10]}), .I3 ({new_AGEMA_signal_3508, ShiftRowsInput[98]}), .O ({new_AGEMA_signal_3900, N242}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[90], plaintext_s0[90]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I4 ({new_AGEMA_signal_3499, ShiftRowsInput[89]}), .I5 ({new_AGEMA_signal_3900, N242}), .O ({new_AGEMA_signal_4123, \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3460, ShiftRowsInput[50]}), .I1 ({new_AGEMA_signal_3500, ShiftRowsInput[90]}), .I2 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I3 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3421, ShiftRowsInput[11]}), .O ({new_AGEMA_signal_3901, N244}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[91], plaintext_s0[91]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3509, ShiftRowsInput[99]}), .I4 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I5 ({new_AGEMA_signal_3901, N244}), .O ({new_AGEMA_signal_4125, \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I1 ({new_AGEMA_signal_3461, ShiftRowsInput[51]}), .I2 ({new_AGEMA_signal_3510, ShiftRowsInput[100]}), .I3 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I4 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I5 ({new_AGEMA_signal_3422, ShiftRowsInput[12]}), .O ({new_AGEMA_signal_3902, N246}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[92], plaintext_s0[92]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I4 ({new_AGEMA_signal_3501, ShiftRowsInput[91]}), .I5 ({new_AGEMA_signal_3902, N246}), .O ({new_AGEMA_signal_4127, \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3462, ShiftRowsInput[52]}), .I1 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I2 ({new_AGEMA_signal_3423, ShiftRowsInput[13]}), .I3 ({new_AGEMA_signal_3511, ShiftRowsInput[101]}), .O ({new_AGEMA_signal_3903, N248}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[93], plaintext_s0[93]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I4 ({new_AGEMA_signal_3502, ShiftRowsInput[92]}), .I5 ({new_AGEMA_signal_3903, N248}), .O ({new_AGEMA_signal_4129, \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I1 ({new_AGEMA_signal_3463, ShiftRowsInput[53]}), .I2 ({new_AGEMA_signal_3424, ShiftRowsInput[14]}), .I3 ({new_AGEMA_signal_3512, ShiftRowsInput[102]}), .O ({new_AGEMA_signal_3904, N250}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[94], plaintext_s0[94]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I4 ({new_AGEMA_signal_3503, ShiftRowsInput[93]}), .I5 ({new_AGEMA_signal_3904, N250}), .O ({new_AGEMA_signal_4131, \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3464, ShiftRowsInput[54]}), .I1 ({new_AGEMA_signal_3513, ShiftRowsInput[103]}), .I2 ({new_AGEMA_signal_3465, ShiftRowsInput[55]}), .I3 ({new_AGEMA_signal_3425, ShiftRowsInput[15]}), .O ({new_AGEMA_signal_3905, N252}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[95], plaintext_s0[95]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3504, ShiftRowsInput[94]}), .I4 ({new_AGEMA_signal_3505, ShiftRowsInput[95]}), .I5 ({new_AGEMA_signal_3905, N252}), .O ({new_AGEMA_signal_4133, \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I1 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I2 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .I3 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3906, N254}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[96], plaintext_s0[96]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I4 ({new_AGEMA_signal_3410, ShiftRowsInput[0]}), .I5 ({new_AGEMA_signal_3906, N254}), .O ({new_AGEMA_signal_4135, \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I1 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I2 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .O ({new_AGEMA_signal_3907, N256}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[97], plaintext_s0[97]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .I4 ({new_AGEMA_signal_3764, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3907, N256}), .O ({new_AGEMA_signal_4137, \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I1 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I2 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .I3 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .O ({new_AGEMA_signal_3908, N258}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[98], plaintext_s0[98]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3412, ShiftRowsInput[2]}), .I4 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .I5 ({new_AGEMA_signal_3908, N258}), .O ({new_AGEMA_signal_4139, \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I1 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I2 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .O ({new_AGEMA_signal_3909, N260}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[99], plaintext_s0[99]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3413, ShiftRowsInput[3]}), .I4 ({new_AGEMA_signal_3765, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3909, N260}), .O ({new_AGEMA_signal_4141, \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I1 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I2 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I3 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I4 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .O ({new_AGEMA_signal_3910, N262}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[100], plaintext_s0[100]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .I4 ({new_AGEMA_signal_3754, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3910, N262}), .O ({new_AGEMA_signal_4143, \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I1 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I2 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I3 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .O ({new_AGEMA_signal_3911, N264}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[101], plaintext_s0[101]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .I4 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .I5 ({new_AGEMA_signal_3911, N264}), .O ({new_AGEMA_signal_4145, \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I1 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I2 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .O ({new_AGEMA_signal_3912, N266}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[102], plaintext_s0[102]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I4 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .I5 ({new_AGEMA_signal_3912, N266}), .O ({new_AGEMA_signal_4147, \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I1 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I2 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I3 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .O ({new_AGEMA_signal_3913, N268}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[103], plaintext_s0[103]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I4 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .I5 ({new_AGEMA_signal_3913, N268}), .O ({new_AGEMA_signal_4149, \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .I1 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I2 ({new_AGEMA_signal_3410, ShiftRowsInput[0]}), .I3 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3914, N270}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[104], plaintext_s0[104]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I4 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I5 ({new_AGEMA_signal_3914, N270}), .O ({new_AGEMA_signal_4151, \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I1 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I2 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .O ({new_AGEMA_signal_3915, N272}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[105], plaintext_s0[105]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I4 ({new_AGEMA_signal_3764, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><1> }), .I5 ({new_AGEMA_signal_3915, N272}), .O ({new_AGEMA_signal_4153, \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .I1 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I2 ({new_AGEMA_signal_3412, ShiftRowsInput[2]}), .I3 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .O ({new_AGEMA_signal_3916, N274}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[106], plaintext_s0[106]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .I4 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I5 ({new_AGEMA_signal_3916, N274}), .O ({new_AGEMA_signal_4155, \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I1 ({new_AGEMA_signal_3413, ShiftRowsInput[3]}), .I2 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .O ({new_AGEMA_signal_3917, N276}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[107], plaintext_s0[107]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .I4 ({new_AGEMA_signal_3765, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><3> }), .I5 ({new_AGEMA_signal_3917, N276}), .O ({new_AGEMA_signal_4157, \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I1 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .I2 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .O ({new_AGEMA_signal_3918, N278}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[108], plaintext_s0[108]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I4 ({new_AGEMA_signal_3754, \MixColumnsIns/GenMixColumns[0].MixOneColumnInst/DoubleBytes<3><4> }), .I5 ({new_AGEMA_signal_3918, N278}), .O ({new_AGEMA_signal_4159, \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I1 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I2 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .O ({new_AGEMA_signal_3919, N280}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[109], plaintext_s0[109]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I4 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .I5 ({new_AGEMA_signal_3919, N280}), .O ({new_AGEMA_signal_4161, \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I1 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I2 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .O ({new_AGEMA_signal_3920, N282}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[110], plaintext_s0[110]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I4 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I5 ({new_AGEMA_signal_3920, N282}), .O ({new_AGEMA_signal_4163, \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I1 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I2 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .I3 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .O ({new_AGEMA_signal_3921, N284}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[111], plaintext_s0[111]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3921, N284}), .O ({new_AGEMA_signal_4165, \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .I1 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I2 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I3 ({new_AGEMA_signal_3410, ShiftRowsInput[0]}), .O ({new_AGEMA_signal_3922, N286}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[112], plaintext_s0[112]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3922, N286}), .O ({new_AGEMA_signal_4167, \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I1 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I2 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .O ({new_AGEMA_signal_3923, N288}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[113], plaintext_s0[113]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I4 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I5 ({new_AGEMA_signal_3923, N288}), .O ({new_AGEMA_signal_4169, \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I1 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .I2 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .I3 ({new_AGEMA_signal_3412, ShiftRowsInput[2]}), .O ({new_AGEMA_signal_3924, N290}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[114], plaintext_s0[114]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I4 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I5 ({new_AGEMA_signal_3924, N290}), .O ({new_AGEMA_signal_4171, \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .I1 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .I2 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I3 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I4 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I5 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .O ({new_AGEMA_signal_3925, N292}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[115], plaintext_s0[115]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I4 ({new_AGEMA_signal_3413, ShiftRowsInput[3]}), .I5 ({new_AGEMA_signal_3925, N292}), .O ({new_AGEMA_signal_4173, \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .I1 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I2 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I3 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .O ({new_AGEMA_signal_3926, N294}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[116], plaintext_s0[116]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I4 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I5 ({new_AGEMA_signal_3926, N294}), .O ({new_AGEMA_signal_4175, \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I1 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I2 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .O ({new_AGEMA_signal_3927, N296}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[117], plaintext_s0[117]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I4 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I5 ({new_AGEMA_signal_3927, N296}), .O ({new_AGEMA_signal_4177, \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I1 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I2 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I3 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .O ({new_AGEMA_signal_3928, N298}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[118], plaintext_s0[118]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I4 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I5 ({new_AGEMA_signal_3928, N298}), .O ({new_AGEMA_signal_4179, \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I1 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I2 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I3 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3929, N300}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB8BB888BBBB88B88 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB8BB888BBBB88B88 ) ) \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[119], plaintext_s0[119]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3929, N300}), .O ({new_AGEMA_signal_4181, \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I1 ({new_AGEMA_signal_3450, ShiftRowsInput[40]}), .I2 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I3 ({new_AGEMA_signal_3410, ShiftRowsInput[0]}), .O ({new_AGEMA_signal_3930, N302}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[120], plaintext_s0[120]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3930, N302}), .O ({new_AGEMA_signal_4183, \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3530, ShiftRowsInput[120]}), .I1 ({new_AGEMA_signal_3490, ShiftRowsInput[80]}), .I2 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3411, ShiftRowsInput[1]}), .O ({new_AGEMA_signal_3931, N304}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[121], plaintext_s0[121]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I4 ({new_AGEMA_signal_3451, ShiftRowsInput[41]}), .I5 ({new_AGEMA_signal_3931, N304}), .O ({new_AGEMA_signal_4185, \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I1 ({new_AGEMA_signal_3491, ShiftRowsInput[81]}), .I2 ({new_AGEMA_signal_3452, ShiftRowsInput[42]}), .I3 ({new_AGEMA_signal_3412, ShiftRowsInput[2]}), .O ({new_AGEMA_signal_3932, N306}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[122], plaintext_s0[122]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .I4 ({new_AGEMA_signal_3531, ShiftRowsInput[121]}), .I5 ({new_AGEMA_signal_3932, N306}), .O ({new_AGEMA_signal_4187, \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3532, ShiftRowsInput[122]}), .I1 ({new_AGEMA_signal_3453, ShiftRowsInput[43]}), .I2 ({new_AGEMA_signal_3492, ShiftRowsInput[82]}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3413, ShiftRowsInput[3]}), .O ({new_AGEMA_signal_3933, N308}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[123], plaintext_s0[123]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I4 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I5 ({new_AGEMA_signal_3933, N308}), .O ({new_AGEMA_signal_4189, \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state }) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3454, ShiftRowsInput[44]}), .I1 ({new_AGEMA_signal_3533, ShiftRowsInput[123]}), .I2 ({new_AGEMA_signal_3493, ShiftRowsInput[83]}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3414, ShiftRowsInput[4]}), .O ({new_AGEMA_signal_3934, N310}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[124], plaintext_s0[124]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I4 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I5 ({new_AGEMA_signal_3934, N310}), .O ({new_AGEMA_signal_4191, \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3534, ShiftRowsInput[124]}), .I1 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I2 ({new_AGEMA_signal_3455, ShiftRowsInput[45]}), .I3 ({new_AGEMA_signal_3415, ShiftRowsInput[5]}), .O ({new_AGEMA_signal_3935, N312}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[125], plaintext_s0[125]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .I4 ({new_AGEMA_signal_3494, ShiftRowsInput[84]}), .I5 ({new_AGEMA_signal_3935, N312}), .O ({new_AGEMA_signal_4193, \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3495, ShiftRowsInput[85]}), .I1 ({new_AGEMA_signal_3456, ShiftRowsInput[46]}), .I2 ({new_AGEMA_signal_3535, ShiftRowsInput[125]}), .I3 ({new_AGEMA_signal_3416, ShiftRowsInput[6]}), .O ({new_AGEMA_signal_3936, N314}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[126], plaintext_s0[126]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I4 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I5 ({new_AGEMA_signal_3936, N314}), .O ({new_AGEMA_signal_4195, \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/MUX_inst/Mmux_Q1_SW0 ( .I0 ({new_AGEMA_signal_3496, ShiftRowsInput[86]}), .I1 ({new_AGEMA_signal_3457, ShiftRowsInput[47]}), .I2 ({new_AGEMA_signal_3536, ShiftRowsInput[126]}), .I3 ({new_AGEMA_signal_3417, ShiftRowsInput[7]}), .O ({new_AGEMA_signal_3937, N316}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB888BB8BBB8BB888 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hB888BB8BBB8BB888 ) ) \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/MUX_inst/Mmux_Q1 ( .I0 ({plaintext_s1[127], plaintext_s0[127]}), .I1 ({1'b0, reset}), .I2 ({1'b0, LastRound}), .I3 ({new_AGEMA_signal_3537, ShiftRowsInput[127]}), .I4 ({new_AGEMA_signal_3497, ShiftRowsInput[87]}), .I5 ({new_AGEMA_signal_3937, N316}), .O ({new_AGEMA_signal_4197, \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'hB88B8BB8 ) , .MASK ( 5'b00010 ), .INIT2 ( 32'hB88B8BB8 ) ) \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[26], key_s0[26]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2666, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_455 }), .I3 ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }), .I4 ({new_AGEMA_signal_3751, KeyExpansionOutput[90]}), .O ({new_AGEMA_signal_3939, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state }) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h8BB8 ) , .MASK ( 4'b0010 ), .INIT2 ( 16'h8BB8 ) ) \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({key_s1[58], key_s0[58]}), .I1 ({1'b0, reset}), .I2 ({new_AGEMA_signal_2666, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_455 }), .I3 ({new_AGEMA_signal_3751, KeyExpansionOutput[90]}), .O ({new_AGEMA_signal_3941, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state }) ) ;
    LUT5_masked #(.low_latency(0), .pipeline(0),  .INIT ( 32'h99966669 ) , .MASK ( 5'b01100 ), .INIT2 ( 32'h99996666 ) ) \KeyExpansionIns/Mxor_OutWords<1>_26_xo<0>1 ( .I0 ({new_AGEMA_signal_2570, \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_423 }), .I1 ({new_AGEMA_signal_2474, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_391 }), .I2 ({1'b0, \RoundCounterIns/count [2]}), .I3 ({1'b0, N318}), .I4 ({new_AGEMA_signal_2879, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [2]}), .O ({new_AGEMA_signal_3751, KeyExpansionOutput[90]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hBEEBBEBE14411414 ) , .MASK ( 6'b011001 ), .INIT2 ( 64'hBEBEBEBE14141414 ) ) \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/MUX_inst/Mmux_Q11 ( .I0 ({1'b0, reset}), .I1 ({new_AGEMA_signal_2474, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_391 }), .I2 ({new_AGEMA_signal_2879, \KeyExpansionIns/KeySchedCoreInst/OutBytes<0> [2]}), .I3 ({1'b0, \RoundCounterIns/count [2]}), .I4 ({1'b0, N320}), .I5 ({key_s1[122], key_s0[122]}), .O ({new_AGEMA_signal_3753, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state }) ) ;

    /* register cells */
    FDR \RoundCounterIns/count_0 ( .D (Result[0]), .C (clk_gated), .R (reset), .Q (\RoundCounterIns/count [0]) ) ;
    FDR \RoundCounterIns/count_1 ( .D (Result[1]), .C (clk_gated), .R (reset), .Q (\RoundCounterIns/count [1]) ) ;
    FDR \RoundCounterIns/count_2 ( .D (Result[2]), .C (clk_gated), .R (reset), .Q (\RoundCounterIns/count [2]) ) ;
    FDR \RoundCounterIns/count_3 ( .D (Result[3]), .C (clk_gated), .R (reset), .Q (\RoundCounterIns/count [3]) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3690, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2420, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_513 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3692, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2421, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_512 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3694, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2422, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_511 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3696, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2423, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_510 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3698, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2424, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_509 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3700, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2425, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_508 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3702, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2822, \KeyReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_507 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3704, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2819, \KeyReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_506 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3706, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2382, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_505 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3708, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2383, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_504 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3710, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2384, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_503 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3712, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2385, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_502 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3714, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2386, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_501 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3716, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2387, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_500 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3718, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2798, \KeyReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_499 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3720, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2795, \KeyReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_498 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3722, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2344, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_497 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3724, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2345, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_496 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3726, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2346, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_495 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3728, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2347, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_494 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3730, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2348, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_493 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3732, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2349, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_492 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3734, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2774, \KeyReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_491 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3736, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2771, \KeyReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_490 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3767, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2306, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_489 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3769, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2307, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_488 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3939, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2308, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_487 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3771, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2309, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_486 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3773, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2310, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_485 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3775, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2311, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_484 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3777, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2750, \KeyReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_483 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3779, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2747, \KeyReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_482 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3546, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2744, \KeyReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_481 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3548, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2741, \KeyReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_480 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3550, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2738, \KeyReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_479 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3552, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2735, \KeyReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_478 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3554, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2732, \KeyReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_477 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3556, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2729, \KeyReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_476 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3558, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2726, \KeyReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_475 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3560, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2723, \KeyReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_474 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3562, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2720, \KeyReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_473 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3564, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2717, \KeyReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_472 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3566, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2714, \KeyReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_471 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3568, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2711, \KeyReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_470 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3570, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2708, \KeyReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_469 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3572, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2705, \KeyReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_468 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3574, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2702, \KeyReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_467 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3576, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2699, \KeyReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_466 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3578, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2696, \KeyReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_465 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3580, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2693, \KeyReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_464 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3582, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2690, \KeyReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_463 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3584, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2687, \KeyReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_462 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3586, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2684, \KeyReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_461 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3588, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2681, \KeyReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_460 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3590, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2678, \KeyReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_459 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3592, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2675, \KeyReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_458 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3781, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2672, \KeyReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_457 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3783, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2669, \KeyReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_456 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3941, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2666, \KeyReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_455 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3785, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2663, \KeyReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_454 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3787, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2660, \KeyReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_453 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3789, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2657, \KeyReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_452 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3791, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2654, \KeyReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_451 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3793, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2651, \KeyReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_450 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3594, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2648, \KeyReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_449 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3596, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2645, \KeyReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_448 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3598, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2642, \KeyReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_447 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3600, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2639, \KeyReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_446 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3602, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2636, \KeyReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_445 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3604, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2633, \KeyReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_444 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3606, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2630, \KeyReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_443 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3608, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2627, \KeyReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_442 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3610, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2624, \KeyReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_441 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3612, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2621, \KeyReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_440 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3614, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2618, \KeyReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_439 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3616, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2615, \KeyReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_438 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3618, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2612, \KeyReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_437 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3620, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2609, \KeyReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_436 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3622, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2606, \KeyReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_435 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3624, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2603, \KeyReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_434 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3626, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2600, \KeyReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_433 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3628, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2597, \KeyReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_432 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3630, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2594, \KeyReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_431 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3632, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2591, \KeyReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_430 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3634, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2588, \KeyReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_429 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3636, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2585, \KeyReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_428 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3638, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2582, \KeyReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_427 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3640, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2579, \KeyReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_426 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3795, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2576, \KeyReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_425 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3797, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2573, \KeyReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_424 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3799, \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2570, \KeyReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_423 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3801, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2567, \KeyReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_422 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3803, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2564, \KeyReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_421 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3805, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2561, \KeyReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_420 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3807, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2558, \KeyReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_419 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3809, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2555, \KeyReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_418 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3642, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2552, \KeyReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_417 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3644, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2549, \KeyReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_416 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3646, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2546, \KeyReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_415 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3648, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2543, \KeyReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_414 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3650, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2540, \KeyReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_413 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3652, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2537, \KeyReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_412 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3654, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2534, \KeyReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_411 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3656, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2531, \KeyReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_410 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3658, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2528, \KeyReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_409 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3660, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2525, \KeyReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_408 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3662, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2522, \KeyReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_407 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3664, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2519, \KeyReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_406 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3666, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2516, \KeyReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_405 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3668, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2513, \KeyReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_404 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3670, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2510, \KeyReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_403 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3672, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2507, \KeyReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_402 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3674, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2504, \KeyReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_401 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3676, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2501, \KeyReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_400 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3678, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2498, \KeyReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_399 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3680, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2495, \KeyReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_398 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3682, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2492, \KeyReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_397 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3684, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2489, \KeyReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_396 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3686, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2486, \KeyReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_395 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3688, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2483, \KeyReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_394 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3738, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2480, \KeyReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_393 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3740, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2477, \KeyReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_392 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3753, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2474, \KeyReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_391 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3742, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2471, \KeyReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_390 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3744, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2468, \KeyReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_389 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3746, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2465, \KeyReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_388 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3748, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2462, \KeyReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_387 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3750, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2459, \KeyReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_386 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3943, \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2839, \RoundReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_385 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3945, \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2836, \RoundReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_384 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3947, \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2833, \RoundReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_383 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3949, \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2830, \RoundReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_382 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3951, \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2827, \RoundReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_381 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3953, \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2824, \RoundReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_380 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3955, \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2821, \RoundReg/gen_Reg_SDE[6].Inst_ff_SDE/current_state_379 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3957, \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2818, \RoundReg/gen_Reg_SDE[7].Inst_ff_SDE/current_state_378 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3959, \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2815, \RoundReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_377 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3961, \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2812, \RoundReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_376 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3963, \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2809, \RoundReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_375 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3965, \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2806, \RoundReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_374 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3967, \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2803, \RoundReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_373 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3969, \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2800, \RoundReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_372 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3971, \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2797, \RoundReg/gen_Reg_SDE[14].Inst_ff_SDE/current_state_371 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3973, \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2794, \RoundReg/gen_Reg_SDE[15].Inst_ff_SDE/current_state_370 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3975, \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2791, \RoundReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_369 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3977, \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2788, \RoundReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_368 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3979, \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2785, \RoundReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_367 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3981, \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2782, \RoundReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_366 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3983, \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2779, \RoundReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_365 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3985, \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2776, \RoundReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_364 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3987, \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2773, \RoundReg/gen_Reg_SDE[22].Inst_ff_SDE/current_state_363 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3989, \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2770, \RoundReg/gen_Reg_SDE[23].Inst_ff_SDE/current_state_362 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3991, \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2767, \RoundReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_361 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3993, \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2764, \RoundReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_360 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3995, \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2761, \RoundReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_359 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3997, \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2758, \RoundReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_358 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_3999, \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2755, \RoundReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_357 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4001, \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2752, \RoundReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_356 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4003, \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2749, \RoundReg/gen_Reg_SDE[30].Inst_ff_SDE/current_state_355 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4005, \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2746, \RoundReg/gen_Reg_SDE[31].Inst_ff_SDE/current_state_354 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4007, \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2743, \RoundReg/gen_Reg_SDE[32].Inst_ff_SDE/current_state_353 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4009, \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2740, \RoundReg/gen_Reg_SDE[33].Inst_ff_SDE/current_state_352 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4011, \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2737, \RoundReg/gen_Reg_SDE[34].Inst_ff_SDE/current_state_351 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4013, \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2734, \RoundReg/gen_Reg_SDE[35].Inst_ff_SDE/current_state_350 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4015, \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2731, \RoundReg/gen_Reg_SDE[36].Inst_ff_SDE/current_state_349 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4017, \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2728, \RoundReg/gen_Reg_SDE[37].Inst_ff_SDE/current_state_348 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4019, \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2725, \RoundReg/gen_Reg_SDE[38].Inst_ff_SDE/current_state_347 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4021, \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2722, \RoundReg/gen_Reg_SDE[39].Inst_ff_SDE/current_state_346 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4023, \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2719, \RoundReg/gen_Reg_SDE[40].Inst_ff_SDE/current_state_345 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4025, \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2716, \RoundReg/gen_Reg_SDE[41].Inst_ff_SDE/current_state_344 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4027, \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2713, \RoundReg/gen_Reg_SDE[42].Inst_ff_SDE/current_state_343 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4029, \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2710, \RoundReg/gen_Reg_SDE[43].Inst_ff_SDE/current_state_342 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4031, \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2707, \RoundReg/gen_Reg_SDE[44].Inst_ff_SDE/current_state_341 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4033, \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2704, \RoundReg/gen_Reg_SDE[45].Inst_ff_SDE/current_state_340 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4035, \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2701, \RoundReg/gen_Reg_SDE[46].Inst_ff_SDE/current_state_339 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4037, \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2698, \RoundReg/gen_Reg_SDE[47].Inst_ff_SDE/current_state_338 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4039, \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2695, \RoundReg/gen_Reg_SDE[48].Inst_ff_SDE/current_state_337 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4041, \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2692, \RoundReg/gen_Reg_SDE[49].Inst_ff_SDE/current_state_336 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4043, \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2689, \RoundReg/gen_Reg_SDE[50].Inst_ff_SDE/current_state_335 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4045, \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2686, \RoundReg/gen_Reg_SDE[51].Inst_ff_SDE/current_state_334 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4047, \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2683, \RoundReg/gen_Reg_SDE[52].Inst_ff_SDE/current_state_333 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4049, \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2680, \RoundReg/gen_Reg_SDE[53].Inst_ff_SDE/current_state_332 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4051, \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2677, \RoundReg/gen_Reg_SDE[54].Inst_ff_SDE/current_state_331 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4053, \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2674, \RoundReg/gen_Reg_SDE[55].Inst_ff_SDE/current_state_330 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4055, \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2671, \RoundReg/gen_Reg_SDE[56].Inst_ff_SDE/current_state_329 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4057, \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2668, \RoundReg/gen_Reg_SDE[57].Inst_ff_SDE/current_state_328 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4059, \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2665, \RoundReg/gen_Reg_SDE[58].Inst_ff_SDE/current_state_327 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4061, \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2662, \RoundReg/gen_Reg_SDE[59].Inst_ff_SDE/current_state_326 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4063, \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2659, \RoundReg/gen_Reg_SDE[60].Inst_ff_SDE/current_state_325 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4065, \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2656, \RoundReg/gen_Reg_SDE[61].Inst_ff_SDE/current_state_324 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4067, \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2653, \RoundReg/gen_Reg_SDE[62].Inst_ff_SDE/current_state_323 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4069, \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2650, \RoundReg/gen_Reg_SDE[63].Inst_ff_SDE/current_state_322 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4071, \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2647, \RoundReg/gen_Reg_SDE[64].Inst_ff_SDE/current_state_321 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4073, \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2644, \RoundReg/gen_Reg_SDE[65].Inst_ff_SDE/current_state_320 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4075, \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2641, \RoundReg/gen_Reg_SDE[66].Inst_ff_SDE/current_state_319 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4077, \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2638, \RoundReg/gen_Reg_SDE[67].Inst_ff_SDE/current_state_318 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4079, \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2635, \RoundReg/gen_Reg_SDE[68].Inst_ff_SDE/current_state_317 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4081, \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2632, \RoundReg/gen_Reg_SDE[69].Inst_ff_SDE/current_state_316 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4083, \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2629, \RoundReg/gen_Reg_SDE[70].Inst_ff_SDE/current_state_315 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4085, \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2626, \RoundReg/gen_Reg_SDE[71].Inst_ff_SDE/current_state_314 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4087, \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2623, \RoundReg/gen_Reg_SDE[72].Inst_ff_SDE/current_state_313 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4089, \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2620, \RoundReg/gen_Reg_SDE[73].Inst_ff_SDE/current_state_312 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4091, \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2617, \RoundReg/gen_Reg_SDE[74].Inst_ff_SDE/current_state_311 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4093, \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2614, \RoundReg/gen_Reg_SDE[75].Inst_ff_SDE/current_state_310 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4095, \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2611, \RoundReg/gen_Reg_SDE[76].Inst_ff_SDE/current_state_309 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4097, \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2608, \RoundReg/gen_Reg_SDE[77].Inst_ff_SDE/current_state_308 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4099, \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2605, \RoundReg/gen_Reg_SDE[78].Inst_ff_SDE/current_state_307 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4101, \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2602, \RoundReg/gen_Reg_SDE[79].Inst_ff_SDE/current_state_306 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4103, \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2599, \RoundReg/gen_Reg_SDE[80].Inst_ff_SDE/current_state_305 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4105, \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2596, \RoundReg/gen_Reg_SDE[81].Inst_ff_SDE/current_state_304 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4107, \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2593, \RoundReg/gen_Reg_SDE[82].Inst_ff_SDE/current_state_303 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4109, \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2590, \RoundReg/gen_Reg_SDE[83].Inst_ff_SDE/current_state_302 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4111, \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2587, \RoundReg/gen_Reg_SDE[84].Inst_ff_SDE/current_state_301 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4113, \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2584, \RoundReg/gen_Reg_SDE[85].Inst_ff_SDE/current_state_300 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4115, \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2581, \RoundReg/gen_Reg_SDE[86].Inst_ff_SDE/current_state_299 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4117, \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2578, \RoundReg/gen_Reg_SDE[87].Inst_ff_SDE/current_state_298 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4119, \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2575, \RoundReg/gen_Reg_SDE[88].Inst_ff_SDE/current_state_297 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4121, \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2572, \RoundReg/gen_Reg_SDE[89].Inst_ff_SDE/current_state_296 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4123, \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2569, \RoundReg/gen_Reg_SDE[90].Inst_ff_SDE/current_state_295 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4125, \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2566, \RoundReg/gen_Reg_SDE[91].Inst_ff_SDE/current_state_294 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4127, \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2563, \RoundReg/gen_Reg_SDE[92].Inst_ff_SDE/current_state_293 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4129, \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2560, \RoundReg/gen_Reg_SDE[93].Inst_ff_SDE/current_state_292 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4131, \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2557, \RoundReg/gen_Reg_SDE[94].Inst_ff_SDE/current_state_291 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4133, \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2554, \RoundReg/gen_Reg_SDE[95].Inst_ff_SDE/current_state_290 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4135, \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2551, \RoundReg/gen_Reg_SDE[96].Inst_ff_SDE/current_state_289 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4137, \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2548, \RoundReg/gen_Reg_SDE[97].Inst_ff_SDE/current_state_288 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4139, \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2545, \RoundReg/gen_Reg_SDE[98].Inst_ff_SDE/current_state_287 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4141, \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2542, \RoundReg/gen_Reg_SDE[99].Inst_ff_SDE/current_state_286 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4143, \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2539, \RoundReg/gen_Reg_SDE[100].Inst_ff_SDE/current_state_285 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4145, \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2536, \RoundReg/gen_Reg_SDE[101].Inst_ff_SDE/current_state_284 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4147, \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2533, \RoundReg/gen_Reg_SDE[102].Inst_ff_SDE/current_state_283 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4149, \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2530, \RoundReg/gen_Reg_SDE[103].Inst_ff_SDE/current_state_282 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4151, \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2527, \RoundReg/gen_Reg_SDE[104].Inst_ff_SDE/current_state_281 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4153, \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2524, \RoundReg/gen_Reg_SDE[105].Inst_ff_SDE/current_state_280 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4155, \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2521, \RoundReg/gen_Reg_SDE[106].Inst_ff_SDE/current_state_279 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4157, \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2518, \RoundReg/gen_Reg_SDE[107].Inst_ff_SDE/current_state_278 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4159, \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2515, \RoundReg/gen_Reg_SDE[108].Inst_ff_SDE/current_state_277 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4161, \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2512, \RoundReg/gen_Reg_SDE[109].Inst_ff_SDE/current_state_276 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4163, \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2509, \RoundReg/gen_Reg_SDE[110].Inst_ff_SDE/current_state_275 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4165, \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2506, \RoundReg/gen_Reg_SDE[111].Inst_ff_SDE/current_state_274 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4167, \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2503, \RoundReg/gen_Reg_SDE[112].Inst_ff_SDE/current_state_273 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4169, \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2500, \RoundReg/gen_Reg_SDE[113].Inst_ff_SDE/current_state_272 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4171, \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2497, \RoundReg/gen_Reg_SDE[114].Inst_ff_SDE/current_state_271 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4173, \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2494, \RoundReg/gen_Reg_SDE[115].Inst_ff_SDE/current_state_270 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4175, \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2491, \RoundReg/gen_Reg_SDE[116].Inst_ff_SDE/current_state_269 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4177, \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2488, \RoundReg/gen_Reg_SDE[117].Inst_ff_SDE/current_state_268 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4179, \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2485, \RoundReg/gen_Reg_SDE[118].Inst_ff_SDE/current_state_267 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4181, \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2482, \RoundReg/gen_Reg_SDE[119].Inst_ff_SDE/current_state_266 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4183, \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2479, \RoundReg/gen_Reg_SDE[120].Inst_ff_SDE/current_state_265 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4185, \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2476, \RoundReg/gen_Reg_SDE[121].Inst_ff_SDE/current_state_264 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4187, \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2473, \RoundReg/gen_Reg_SDE[122].Inst_ff_SDE/current_state_263 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4189, \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2470, \RoundReg/gen_Reg_SDE[123].Inst_ff_SDE/current_state_262 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4191, \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2467, \RoundReg/gen_Reg_SDE[124].Inst_ff_SDE/current_state_261 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4193, \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2464, \RoundReg/gen_Reg_SDE[125].Inst_ff_SDE/current_state_260 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4195, \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2461, \RoundReg/gen_Reg_SDE[126].Inst_ff_SDE/current_state_259 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state ( .D ({new_AGEMA_signal_4197, \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2458, \RoundReg/gen_Reg_SDE[127].Inst_ff_SDE/current_state_258 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3722, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2792, \KeyReg/gen_Reg_SDE[16].Inst_ff_SDE/current_state_1_2276 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3724, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2789, \KeyReg/gen_Reg_SDE[17].Inst_ff_SDE/current_state_1_2277 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3726, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2786, \KeyReg/gen_Reg_SDE[18].Inst_ff_SDE/current_state_1_2278 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3728, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2783, \KeyReg/gen_Reg_SDE[19].Inst_ff_SDE/current_state_1_2279 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3730, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2780, \KeyReg/gen_Reg_SDE[20].Inst_ff_SDE/current_state_1_2280 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3732, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2777, \KeyReg/gen_Reg_SDE[21].Inst_ff_SDE/current_state_1_2281 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3767, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2768, \KeyReg/gen_Reg_SDE[24].Inst_ff_SDE/current_state_1_2282 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3769, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2765, \KeyReg/gen_Reg_SDE[25].Inst_ff_SDE/current_state_1_2283 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3771, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2759, \KeyReg/gen_Reg_SDE[27].Inst_ff_SDE/current_state_1_2284 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3773, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2756, \KeyReg/gen_Reg_SDE[28].Inst_ff_SDE/current_state_1_2285 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3775, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2753, \KeyReg/gen_Reg_SDE[29].Inst_ff_SDE/current_state_1_2286 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3690, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2840, \KeyReg/gen_Reg_SDE[0].Inst_ff_SDE/current_state_1_2287 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3692, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2837, \KeyReg/gen_Reg_SDE[1].Inst_ff_SDE/current_state_1_2288 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3694, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2834, \KeyReg/gen_Reg_SDE[2].Inst_ff_SDE/current_state_1_2289 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3696, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2831, \KeyReg/gen_Reg_SDE[3].Inst_ff_SDE/current_state_1_2290 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3698, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2828, \KeyReg/gen_Reg_SDE[4].Inst_ff_SDE/current_state_1_2291 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3700, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2825, \KeyReg/gen_Reg_SDE[5].Inst_ff_SDE/current_state_1_2292 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3706, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2816, \KeyReg/gen_Reg_SDE[8].Inst_ff_SDE/current_state_1_2293 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3708, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2813, \KeyReg/gen_Reg_SDE[9].Inst_ff_SDE/current_state_1_2294 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3710, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2810, \KeyReg/gen_Reg_SDE[10].Inst_ff_SDE/current_state_1_2295 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3712, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2807, \KeyReg/gen_Reg_SDE[11].Inst_ff_SDE/current_state_1_2296 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3714, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2804, \KeyReg/gen_Reg_SDE[12].Inst_ff_SDE/current_state_1_2297 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3716, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2801, \KeyReg/gen_Reg_SDE[13].Inst_ff_SDE/current_state_1_2298 }) ) ;
    FD_masked #(.low_latency(0), .pipeline(0)) \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_1 ( .D ({new_AGEMA_signal_3939, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/next_state }), .clk (clk_gated), .Q ({new_AGEMA_signal_2762, \KeyReg/gen_Reg_SDE[26].Inst_ff_SDE/current_state_1_2299 }) ) ;
endmodule
