/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module AES_HPC2_AIG_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [679:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_423 ;
    wire signal_425 ;
    wire signal_427 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_443 ;
    wire signal_445 ;
    wire signal_447 ;
    wire signal_449 ;
    wire signal_451 ;
    wire signal_453 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_459 ;
    wire signal_461 ;
    wire signal_463 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3874 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3882 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3890 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3898 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3906 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3914 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3922 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3930 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3938 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3946 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3954 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3962 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3970 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3978 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3986 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4394 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4402 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4410 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4474 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4482 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4490 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4498 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4506 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4514 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;
    wire signal_8952 ;
    wire signal_8953 ;
    wire signal_8954 ;
    wire signal_8955 ;
    wire signal_8956 ;
    wire signal_8957 ;
    wire signal_8958 ;
    wire signal_8959 ;
    wire signal_8960 ;
    wire signal_8961 ;
    wire signal_8962 ;
    wire signal_8963 ;
    wire signal_8964 ;
    wire signal_8965 ;
    wire signal_8966 ;
    wire signal_8967 ;
    wire signal_8968 ;
    wire signal_8969 ;
    wire signal_8970 ;
    wire signal_8971 ;
    wire signal_8972 ;
    wire signal_8973 ;
    wire signal_8974 ;
    wire signal_8975 ;
    wire signal_8976 ;
    wire signal_8977 ;
    wire signal_8978 ;
    wire signal_8979 ;
    wire signal_8980 ;
    wire signal_8981 ;
    wire signal_8982 ;
    wire signal_8983 ;
    wire signal_8984 ;
    wire signal_8985 ;
    wire signal_8986 ;
    wire signal_8987 ;
    wire signal_8988 ;
    wire signal_8989 ;
    wire signal_8990 ;
    wire signal_8991 ;
    wire signal_8992 ;
    wire signal_8993 ;
    wire signal_8994 ;
    wire signal_8995 ;
    wire signal_8996 ;
    wire signal_8997 ;
    wire signal_8998 ;
    wire signal_8999 ;
    wire signal_9000 ;
    wire signal_9001 ;
    wire signal_9002 ;
    wire signal_9003 ;
    wire signal_9004 ;
    wire signal_9005 ;
    wire signal_9006 ;
    wire signal_9007 ;
    wire signal_9008 ;
    wire signal_9009 ;
    wire signal_9010 ;
    wire signal_9011 ;
    wire signal_9012 ;
    wire signal_9013 ;
    wire signal_9014 ;
    wire signal_9015 ;
    wire signal_9016 ;
    wire signal_9017 ;
    wire signal_9018 ;
    wire signal_9019 ;
    wire signal_9020 ;
    wire signal_9021 ;
    wire signal_9022 ;
    wire signal_9023 ;
    wire signal_9024 ;
    wire signal_9025 ;
    wire signal_9026 ;
    wire signal_9027 ;
    wire signal_9028 ;
    wire signal_9029 ;
    wire signal_9030 ;
    wire signal_9031 ;
    wire signal_9032 ;
    wire signal_9033 ;
    wire signal_9034 ;
    wire signal_9035 ;
    wire signal_9036 ;
    wire signal_9037 ;
    wire signal_9038 ;
    wire signal_9039 ;
    wire signal_9040 ;
    wire signal_9041 ;
    wire signal_9042 ;
    wire signal_9043 ;
    wire signal_9044 ;
    wire signal_9045 ;
    wire signal_9046 ;
    wire signal_9047 ;
    wire signal_9048 ;
    wire signal_9049 ;
    wire signal_9050 ;
    wire signal_9051 ;
    wire signal_9052 ;
    wire signal_9053 ;
    wire signal_9054 ;
    wire signal_9055 ;
    wire signal_9056 ;
    wire signal_9057 ;
    wire signal_9058 ;
    wire signal_9059 ;
    wire signal_9060 ;
    wire signal_9061 ;
    wire signal_9062 ;
    wire signal_9063 ;
    wire signal_9064 ;
    wire signal_9065 ;
    wire signal_9066 ;
    wire signal_9067 ;
    wire signal_9068 ;
    wire signal_9069 ;
    wire signal_9070 ;
    wire signal_9071 ;
    wire signal_9072 ;
    wire signal_9073 ;
    wire signal_9074 ;
    wire signal_9075 ;
    wire signal_9076 ;
    wire signal_9077 ;
    wire signal_9078 ;
    wire signal_9079 ;
    wire signal_9080 ;
    wire signal_9081 ;
    wire signal_9082 ;
    wire signal_9083 ;
    wire signal_9084 ;
    wire signal_9085 ;
    wire signal_9086 ;
    wire signal_9087 ;
    wire signal_9088 ;
    wire signal_9089 ;
    wire signal_9090 ;
    wire signal_9091 ;
    wire signal_9092 ;
    wire signal_9093 ;
    wire signal_9094 ;
    wire signal_9095 ;
    wire signal_9096 ;
    wire signal_9097 ;
    wire signal_9098 ;
    wire signal_9099 ;
    wire signal_9100 ;
    wire signal_9101 ;
    wire signal_9102 ;
    wire signal_9103 ;
    wire signal_9104 ;
    wire signal_9105 ;
    wire signal_9106 ;
    wire signal_9107 ;
    wire signal_9108 ;
    wire signal_9109 ;
    wire signal_9110 ;
    wire signal_9111 ;
    wire signal_9112 ;
    wire signal_9113 ;
    wire signal_9114 ;
    wire signal_9115 ;
    wire signal_9116 ;
    wire signal_9117 ;
    wire signal_9118 ;
    wire signal_9119 ;
    wire signal_9120 ;
    wire signal_9121 ;
    wire signal_9122 ;
    wire signal_9123 ;
    wire signal_9124 ;
    wire signal_9125 ;
    wire signal_9126 ;
    wire signal_9127 ;
    wire signal_9128 ;
    wire signal_9129 ;
    wire signal_9130 ;
    wire signal_9131 ;
    wire signal_9132 ;
    wire signal_9133 ;
    wire signal_9134 ;
    wire signal_9135 ;
    wire signal_9136 ;
    wire signal_9137 ;
    wire signal_9138 ;
    wire signal_9139 ;
    wire signal_9140 ;
    wire signal_9141 ;
    wire signal_9142 ;
    wire signal_9143 ;
    wire signal_9144 ;
    wire signal_9145 ;
    wire signal_9146 ;
    wire signal_9147 ;
    wire signal_9148 ;
    wire signal_9149 ;
    wire signal_9150 ;
    wire signal_9151 ;
    wire signal_9152 ;
    wire signal_9153 ;
    wire signal_9154 ;
    wire signal_9155 ;
    wire signal_9156 ;
    wire signal_9157 ;
    wire signal_9158 ;
    wire signal_9159 ;
    wire signal_9160 ;
    wire signal_9161 ;
    wire signal_9162 ;
    wire signal_9163 ;
    wire signal_9164 ;
    wire signal_9165 ;
    wire signal_9166 ;
    wire signal_9167 ;
    wire signal_9168 ;
    wire signal_9169 ;
    wire signal_9170 ;
    wire signal_9171 ;
    wire signal_9172 ;
    wire signal_9173 ;
    wire signal_9174 ;
    wire signal_9175 ;
    wire signal_9176 ;
    wire signal_9177 ;
    wire signal_9178 ;
    wire signal_9179 ;
    wire signal_9180 ;
    wire signal_9181 ;
    wire signal_9182 ;
    wire signal_9183 ;
    wire signal_9184 ;
    wire signal_9185 ;
    wire signal_9186 ;
    wire signal_9187 ;
    wire signal_9188 ;
    wire signal_9189 ;
    wire signal_9190 ;
    wire signal_9191 ;
    wire signal_9192 ;
    wire signal_9193 ;
    wire signal_9194 ;
    wire signal_9195 ;
    wire signal_9196 ;
    wire signal_9197 ;
    wire signal_9198 ;
    wire signal_9199 ;
    wire signal_9200 ;
    wire signal_9201 ;
    wire signal_9202 ;
    wire signal_9203 ;
    wire signal_9204 ;
    wire signal_9205 ;
    wire signal_9206 ;
    wire signal_9207 ;
    wire signal_9208 ;
    wire signal_9209 ;
    wire signal_9210 ;
    wire signal_9211 ;
    wire signal_9212 ;
    wire signal_9213 ;
    wire signal_9214 ;
    wire signal_9215 ;
    wire signal_9216 ;
    wire signal_9217 ;
    wire signal_9218 ;
    wire signal_9219 ;
    wire signal_9220 ;
    wire signal_9221 ;
    wire signal_9222 ;
    wire signal_9223 ;
    wire signal_9224 ;
    wire signal_9225 ;
    wire signal_9226 ;
    wire signal_9227 ;
    wire signal_9228 ;
    wire signal_9229 ;
    wire signal_9230 ;
    wire signal_9231 ;
    wire signal_9232 ;
    wire signal_9233 ;
    wire signal_9234 ;
    wire signal_9235 ;
    wire signal_9236 ;
    wire signal_9237 ;
    wire signal_9238 ;
    wire signal_9239 ;
    wire signal_9240 ;
    wire signal_9241 ;
    wire signal_9242 ;
    wire signal_9243 ;
    wire signal_9244 ;
    wire signal_9245 ;
    wire signal_9246 ;
    wire signal_9247 ;
    wire signal_9248 ;
    wire signal_9249 ;
    wire signal_9250 ;
    wire signal_9251 ;
    wire signal_9252 ;
    wire signal_9253 ;
    wire signal_9254 ;
    wire signal_9255 ;
    wire signal_9256 ;
    wire signal_9257 ;
    wire signal_9258 ;
    wire signal_9259 ;
    wire signal_9260 ;
    wire signal_9261 ;
    wire signal_9262 ;
    wire signal_9263 ;
    wire signal_9264 ;
    wire signal_9265 ;
    wire signal_9266 ;
    wire signal_9267 ;
    wire signal_9268 ;
    wire signal_9269 ;
    wire signal_9270 ;
    wire signal_9271 ;
    wire signal_9272 ;
    wire signal_9273 ;
    wire signal_9274 ;
    wire signal_9275 ;
    wire signal_9276 ;
    wire signal_9277 ;
    wire signal_9278 ;
    wire signal_9279 ;
    wire signal_9280 ;
    wire signal_9281 ;
    wire signal_9282 ;
    wire signal_9283 ;
    wire signal_9284 ;
    wire signal_9285 ;
    wire signal_9286 ;
    wire signal_9287 ;
    wire signal_9288 ;
    wire signal_9289 ;
    wire signal_9290 ;
    wire signal_9291 ;
    wire signal_9292 ;
    wire signal_9293 ;
    wire signal_9294 ;
    wire signal_9295 ;
    wire signal_9296 ;
    wire signal_9297 ;
    wire signal_9298 ;
    wire signal_9299 ;
    wire signal_9300 ;
    wire signal_9301 ;
    wire signal_9302 ;
    wire signal_9303 ;
    wire signal_9304 ;
    wire signal_9305 ;
    wire signal_9306 ;
    wire signal_9307 ;
    wire signal_9308 ;
    wire signal_9309 ;
    wire signal_9310 ;
    wire signal_9311 ;
    wire signal_9312 ;
    wire signal_9313 ;
    wire signal_9314 ;
    wire signal_9315 ;
    wire signal_9316 ;
    wire signal_9317 ;
    wire signal_9318 ;
    wire signal_9319 ;
    wire signal_9320 ;
    wire signal_9321 ;
    wire signal_9322 ;
    wire signal_9323 ;
    wire signal_9324 ;
    wire signal_9325 ;
    wire signal_9326 ;
    wire signal_9327 ;
    wire signal_9328 ;
    wire signal_9329 ;
    wire signal_9330 ;
    wire signal_9331 ;
    wire signal_9332 ;
    wire signal_9333 ;
    wire signal_9334 ;
    wire signal_9335 ;
    wire signal_9336 ;
    wire signal_9337 ;
    wire signal_9338 ;
    wire signal_9339 ;
    wire signal_9340 ;
    wire signal_9341 ;
    wire signal_9342 ;
    wire signal_9343 ;
    wire signal_9344 ;
    wire signal_9345 ;
    wire signal_9346 ;
    wire signal_9347 ;
    wire signal_9348 ;
    wire signal_9349 ;
    wire signal_9350 ;
    wire signal_9351 ;
    wire signal_9352 ;
    wire signal_9353 ;
    wire signal_9354 ;
    wire signal_9355 ;
    wire signal_9356 ;
    wire signal_9357 ;
    wire signal_9358 ;
    wire signal_9359 ;
    wire signal_9360 ;
    wire signal_9361 ;
    wire signal_9362 ;
    wire signal_9363 ;
    wire signal_9364 ;
    wire signal_9365 ;
    wire signal_9366 ;
    wire signal_9367 ;
    wire signal_9368 ;
    wire signal_9369 ;
    wire signal_9370 ;
    wire signal_9371 ;
    wire signal_9372 ;
    wire signal_9373 ;
    wire signal_9374 ;
    wire signal_9375 ;
    wire signal_9376 ;
    wire signal_9377 ;
    wire signal_9378 ;
    wire signal_9379 ;
    wire signal_9380 ;
    wire signal_9381 ;
    wire signal_9382 ;
    wire signal_9383 ;
    wire signal_9384 ;
    wire signal_9385 ;
    wire signal_9386 ;
    wire signal_9387 ;
    wire signal_9388 ;
    wire signal_9389 ;
    wire signal_9390 ;
    wire signal_9391 ;
    wire signal_9392 ;
    wire signal_9393 ;
    wire signal_9394 ;
    wire signal_9395 ;
    wire signal_9396 ;
    wire signal_9397 ;
    wire signal_9398 ;
    wire signal_9399 ;
    wire signal_9400 ;
    wire signal_9401 ;
    wire signal_9402 ;
    wire signal_9403 ;
    wire signal_9404 ;
    wire signal_9405 ;
    wire signal_9406 ;
    wire signal_9407 ;
    wire signal_9408 ;
    wire signal_9409 ;
    wire signal_9410 ;
    wire signal_9411 ;
    wire signal_9412 ;
    wire signal_9413 ;
    wire signal_9414 ;
    wire signal_9415 ;
    wire signal_9416 ;
    wire signal_9417 ;
    wire signal_9418 ;
    wire signal_9419 ;
    wire signal_9420 ;
    wire signal_9421 ;
    wire signal_9422 ;
    wire signal_9423 ;
    wire signal_9424 ;
    wire signal_9425 ;
    wire signal_9426 ;
    wire signal_9427 ;
    wire signal_9428 ;
    wire signal_9429 ;
    wire signal_9430 ;
    wire signal_9431 ;
    wire signal_9432 ;
    wire signal_9433 ;
    wire signal_9434 ;
    wire signal_9435 ;
    wire signal_9436 ;
    wire signal_9437 ;
    wire signal_9438 ;
    wire signal_9439 ;
    wire signal_9440 ;
    wire signal_9441 ;
    wire signal_9442 ;
    wire signal_9443 ;
    wire signal_9444 ;
    wire signal_9445 ;
    wire signal_9446 ;
    wire signal_9447 ;
    wire signal_9448 ;
    wire signal_9449 ;
    wire signal_9450 ;
    wire signal_9451 ;
    wire signal_9452 ;
    wire signal_9453 ;
    wire signal_9454 ;
    wire signal_9455 ;
    wire signal_9456 ;
    wire signal_9457 ;
    wire signal_9458 ;
    wire signal_9459 ;
    wire signal_9460 ;
    wire signal_9461 ;
    wire signal_9462 ;
    wire signal_9463 ;
    wire signal_9464 ;
    wire signal_9465 ;
    wire signal_9466 ;
    wire signal_9467 ;
    wire signal_9468 ;
    wire signal_9469 ;
    wire signal_9470 ;
    wire signal_9471 ;
    wire signal_9472 ;
    wire signal_9473 ;
    wire signal_9474 ;
    wire signal_9475 ;
    wire signal_9476 ;
    wire signal_9477 ;
    wire signal_9478 ;
    wire signal_9479 ;
    wire signal_9480 ;
    wire signal_9481 ;
    wire signal_9482 ;
    wire signal_9483 ;
    wire signal_9484 ;
    wire signal_9485 ;
    wire signal_9486 ;
    wire signal_9487 ;
    wire signal_9488 ;
    wire signal_9489 ;
    wire signal_9490 ;
    wire signal_9491 ;
    wire signal_9492 ;
    wire signal_9493 ;
    wire signal_9494 ;
    wire signal_9495 ;
    wire signal_9496 ;
    wire signal_9497 ;
    wire signal_9498 ;
    wire signal_9499 ;
    wire signal_9500 ;
    wire signal_9501 ;
    wire signal_9502 ;
    wire signal_9503 ;
    wire signal_9504 ;
    wire signal_9505 ;
    wire signal_9506 ;
    wire signal_9507 ;
    wire signal_9508 ;
    wire signal_9509 ;
    wire signal_9510 ;
    wire signal_9511 ;
    wire signal_9512 ;
    wire signal_9513 ;
    wire signal_9514 ;
    wire signal_9515 ;
    wire signal_9516 ;
    wire signal_9517 ;
    wire signal_9518 ;
    wire signal_9519 ;
    wire signal_9520 ;
    wire signal_9521 ;
    wire signal_9522 ;
    wire signal_9523 ;
    wire signal_9524 ;
    wire signal_9525 ;
    wire signal_9526 ;
    wire signal_9527 ;
    wire signal_9528 ;
    wire signal_9529 ;
    wire signal_9530 ;
    wire signal_9531 ;
    wire signal_9532 ;
    wire signal_9533 ;
    wire signal_9534 ;
    wire signal_9535 ;
    wire signal_9536 ;
    wire signal_9537 ;
    wire signal_9538 ;
    wire signal_9539 ;
    wire signal_9540 ;
    wire signal_9541 ;
    wire signal_9542 ;
    wire signal_9543 ;
    wire signal_9544 ;
    wire signal_9545 ;
    wire signal_9546 ;
    wire signal_9547 ;
    wire signal_9548 ;
    wire signal_9549 ;
    wire signal_9550 ;
    wire signal_9551 ;
    wire signal_9552 ;
    wire signal_9553 ;
    wire signal_9554 ;
    wire signal_9555 ;
    wire signal_9556 ;
    wire signal_9557 ;
    wire signal_9558 ;
    wire signal_9559 ;
    wire signal_9560 ;
    wire signal_9561 ;
    wire signal_9562 ;
    wire signal_9563 ;
    wire signal_9564 ;
    wire signal_9565 ;
    wire signal_9566 ;
    wire signal_9567 ;
    wire signal_9568 ;
    wire signal_9569 ;
    wire signal_9570 ;
    wire signal_9571 ;
    wire signal_9572 ;
    wire signal_9573 ;
    wire signal_9574 ;
    wire signal_9575 ;
    wire signal_9576 ;
    wire signal_9577 ;
    wire signal_9578 ;
    wire signal_9579 ;
    wire signal_9580 ;
    wire signal_9581 ;
    wire signal_9582 ;
    wire signal_9583 ;
    wire signal_9584 ;
    wire signal_9585 ;
    wire signal_9586 ;
    wire signal_9587 ;
    wire signal_9588 ;
    wire signal_9589 ;
    wire signal_9590 ;
    wire signal_9591 ;
    wire signal_9592 ;
    wire signal_9593 ;
    wire signal_9594 ;
    wire signal_9595 ;
    wire signal_9596 ;
    wire signal_9597 ;
    wire signal_9598 ;
    wire signal_9599 ;
    wire signal_9600 ;
    wire signal_9601 ;
    wire signal_9602 ;
    wire signal_9603 ;
    wire signal_9604 ;
    wire signal_9605 ;
    wire signal_9606 ;
    wire signal_9607 ;
    wire signal_9608 ;
    wire signal_9609 ;
    wire signal_9610 ;
    wire signal_9611 ;
    wire signal_9612 ;
    wire signal_9613 ;
    wire signal_9614 ;
    wire signal_9615 ;
    wire signal_9616 ;
    wire signal_9617 ;
    wire signal_9618 ;
    wire signal_9619 ;
    wire signal_9620 ;
    wire signal_9621 ;
    wire signal_9622 ;
    wire signal_9623 ;
    wire signal_9624 ;
    wire signal_9625 ;
    wire signal_9626 ;
    wire signal_9627 ;
    wire signal_9628 ;
    wire signal_9629 ;
    wire signal_9630 ;
    wire signal_9631 ;
    wire signal_9632 ;
    wire signal_9633 ;
    wire signal_9634 ;
    wire signal_9635 ;
    wire signal_9636 ;
    wire signal_9637 ;
    wire signal_9638 ;
    wire signal_9639 ;
    wire signal_9640 ;
    wire signal_9641 ;
    wire signal_9642 ;
    wire signal_9643 ;
    wire signal_9644 ;
    wire signal_9645 ;
    wire signal_9646 ;
    wire signal_9647 ;
    wire signal_9648 ;
    wire signal_9649 ;
    wire signal_9650 ;
    wire signal_9651 ;
    wire signal_9652 ;
    wire signal_9653 ;
    wire signal_9654 ;
    wire signal_9655 ;
    wire signal_9656 ;
    wire signal_9657 ;
    wire signal_9658 ;
    wire signal_9659 ;
    wire signal_9660 ;
    wire signal_9661 ;
    wire signal_9662 ;
    wire signal_9663 ;
    wire signal_9664 ;
    wire signal_9665 ;
    wire signal_9666 ;
    wire signal_9667 ;
    wire signal_9668 ;
    wire signal_9669 ;
    wire signal_9670 ;
    wire signal_9671 ;
    wire signal_9672 ;
    wire signal_9673 ;
    wire signal_9674 ;
    wire signal_9675 ;
    wire signal_9676 ;
    wire signal_9677 ;
    wire signal_9678 ;
    wire signal_9679 ;
    wire signal_9680 ;
    wire signal_9681 ;
    wire signal_9682 ;
    wire signal_9683 ;
    wire signal_9684 ;
    wire signal_9685 ;
    wire signal_9686 ;
    wire signal_9687 ;
    wire signal_9688 ;
    wire signal_9689 ;
    wire signal_9690 ;
    wire signal_9691 ;
    wire signal_9692 ;
    wire signal_9693 ;
    wire signal_9694 ;
    wire signal_9695 ;
    wire signal_9696 ;
    wire signal_9697 ;
    wire signal_9698 ;
    wire signal_9699 ;
    wire signal_9700 ;
    wire signal_9701 ;
    wire signal_9702 ;
    wire signal_9703 ;
    wire signal_9704 ;
    wire signal_9705 ;
    wire signal_9706 ;
    wire signal_9707 ;
    wire signal_9708 ;
    wire signal_9709 ;
    wire signal_9710 ;
    wire signal_9711 ;
    wire signal_9712 ;
    wire signal_9713 ;
    wire signal_9714 ;
    wire signal_9715 ;
    wire signal_9716 ;
    wire signal_9717 ;
    wire signal_9718 ;
    wire signal_9719 ;
    wire signal_9720 ;
    wire signal_9721 ;
    wire signal_9722 ;
    wire signal_9723 ;
    wire signal_9724 ;
    wire signal_9725 ;
    wire signal_9726 ;
    wire signal_9727 ;
    wire signal_9728 ;
    wire signal_9729 ;
    wire signal_9730 ;
    wire signal_9731 ;
    wire signal_9732 ;
    wire signal_9733 ;
    wire signal_9734 ;
    wire signal_9735 ;
    wire signal_9736 ;
    wire signal_9737 ;
    wire signal_9738 ;
    wire signal_9739 ;
    wire signal_9740 ;
    wire signal_9741 ;
    wire signal_9742 ;
    wire signal_9743 ;
    wire signal_9744 ;
    wire signal_9745 ;
    wire signal_9746 ;
    wire signal_9747 ;
    wire signal_9748 ;
    wire signal_9749 ;
    wire signal_9750 ;
    wire signal_9751 ;
    wire signal_9752 ;
    wire signal_9753 ;
    wire signal_9754 ;
    wire signal_9755 ;
    wire signal_9756 ;
    wire signal_9757 ;
    wire signal_9758 ;
    wire signal_9759 ;
    wire signal_9760 ;
    wire signal_9761 ;
    wire signal_9762 ;
    wire signal_9763 ;
    wire signal_9764 ;
    wire signal_9765 ;
    wire signal_9766 ;
    wire signal_9767 ;
    wire signal_9768 ;
    wire signal_9769 ;
    wire signal_9770 ;
    wire signal_9771 ;
    wire signal_9772 ;
    wire signal_9773 ;
    wire signal_9774 ;
    wire signal_9775 ;
    wire signal_9776 ;
    wire signal_9777 ;
    wire signal_9778 ;
    wire signal_9779 ;
    wire signal_9780 ;
    wire signal_9781 ;
    wire signal_9782 ;
    wire signal_9783 ;
    wire signal_9784 ;
    wire signal_9785 ;
    wire signal_9786 ;
    wire signal_9787 ;
    wire signal_9788 ;
    wire signal_9789 ;
    wire signal_9790 ;
    wire signal_9791 ;
    wire signal_9792 ;
    wire signal_9793 ;
    wire signal_9794 ;
    wire signal_9795 ;
    wire signal_9796 ;
    wire signal_9797 ;
    wire signal_9798 ;
    wire signal_9799 ;
    wire signal_9800 ;
    wire signal_9801 ;
    wire signal_9802 ;
    wire signal_9803 ;
    wire signal_9804 ;
    wire signal_9805 ;
    wire signal_9806 ;
    wire signal_9807 ;
    wire signal_9808 ;
    wire signal_9809 ;
    wire signal_9810 ;
    wire signal_9811 ;
    wire signal_9812 ;
    wire signal_9813 ;
    wire signal_9814 ;
    wire signal_9815 ;
    wire signal_9816 ;
    wire signal_9817 ;
    wire signal_9818 ;
    wire signal_9819 ;
    wire signal_9820 ;
    wire signal_9821 ;
    wire signal_9822 ;
    wire signal_9823 ;
    wire signal_9824 ;
    wire signal_9825 ;
    wire signal_9826 ;
    wire signal_9827 ;
    wire signal_9828 ;
    wire signal_9829 ;
    wire signal_9830 ;
    wire signal_9831 ;
    wire signal_9832 ;
    wire signal_9833 ;
    wire signal_9834 ;
    wire signal_9835 ;
    wire signal_9836 ;
    wire signal_9837 ;
    wire signal_9838 ;
    wire signal_9839 ;
    wire signal_9840 ;
    wire signal_9841 ;
    wire signal_9842 ;
    wire signal_9843 ;
    wire signal_9844 ;
    wire signal_9845 ;
    wire signal_9846 ;
    wire signal_9847 ;
    wire signal_9848 ;
    wire signal_9849 ;
    wire signal_9850 ;
    wire signal_9851 ;
    wire signal_9852 ;
    wire signal_9853 ;
    wire signal_9854 ;
    wire signal_9855 ;
    wire signal_9856 ;
    wire signal_9857 ;
    wire signal_9858 ;
    wire signal_9859 ;
    wire signal_9860 ;
    wire signal_9861 ;
    wire signal_9862 ;
    wire signal_9863 ;
    wire signal_9864 ;
    wire signal_9865 ;
    wire signal_9866 ;
    wire signal_9867 ;
    wire signal_9868 ;
    wire signal_9869 ;
    wire signal_9870 ;
    wire signal_9871 ;
    wire signal_9872 ;
    wire signal_9873 ;
    wire signal_9874 ;
    wire signal_9875 ;
    wire signal_9876 ;
    wire signal_9877 ;
    wire signal_9878 ;
    wire signal_9879 ;
    wire signal_9880 ;
    wire signal_9881 ;
    wire signal_9882 ;
    wire signal_9883 ;
    wire signal_9884 ;
    wire signal_9885 ;
    wire signal_9886 ;
    wire signal_9887 ;
    wire signal_9888 ;
    wire signal_9889 ;
    wire signal_9890 ;
    wire signal_9891 ;
    wire signal_9892 ;
    wire signal_9893 ;
    wire signal_9894 ;
    wire signal_9895 ;
    wire signal_9896 ;
    wire signal_9897 ;
    wire signal_9898 ;
    wire signal_9899 ;
    wire signal_9900 ;
    wire signal_9901 ;
    wire signal_9902 ;
    wire signal_9903 ;
    wire signal_9904 ;
    wire signal_9905 ;
    wire signal_9906 ;
    wire signal_9907 ;
    wire signal_9908 ;
    wire signal_9909 ;
    wire signal_9910 ;
    wire signal_9911 ;
    wire signal_9912 ;
    wire signal_9913 ;
    wire signal_9914 ;
    wire signal_9915 ;
    wire signal_9916 ;
    wire signal_9917 ;
    wire signal_9918 ;
    wire signal_9919 ;
    wire signal_9920 ;
    wire signal_9921 ;
    wire signal_9922 ;
    wire signal_9923 ;
    wire signal_9924 ;
    wire signal_9925 ;
    wire signal_9926 ;
    wire signal_9927 ;
    wire signal_9928 ;
    wire signal_9929 ;
    wire signal_9930 ;
    wire signal_9931 ;
    wire signal_9932 ;
    wire signal_9933 ;
    wire signal_9934 ;
    wire signal_9935 ;
    wire signal_9936 ;
    wire signal_9937 ;
    wire signal_9938 ;
    wire signal_9939 ;
    wire signal_9940 ;
    wire signal_9941 ;
    wire signal_9942 ;
    wire signal_9943 ;
    wire signal_9944 ;
    wire signal_9945 ;
    wire signal_9946 ;
    wire signal_9947 ;
    wire signal_9948 ;
    wire signal_9949 ;
    wire signal_9950 ;
    wire signal_9951 ;
    wire signal_9952 ;
    wire signal_9953 ;
    wire signal_9954 ;
    wire signal_9955 ;
    wire signal_9956 ;
    wire signal_9957 ;
    wire signal_9958 ;
    wire signal_9959 ;
    wire signal_9960 ;
    wire signal_9961 ;
    wire signal_9962 ;
    wire signal_9963 ;
    wire signal_9964 ;
    wire signal_9965 ;
    wire signal_9966 ;
    wire signal_9967 ;
    wire signal_9968 ;
    wire signal_9969 ;
    wire signal_9970 ;
    wire signal_9971 ;
    wire signal_9972 ;
    wire signal_9973 ;
    wire signal_9974 ;
    wire signal_9975 ;
    wire signal_9976 ;
    wire signal_9977 ;
    wire signal_9978 ;
    wire signal_9979 ;
    wire signal_9980 ;
    wire signal_9981 ;
    wire signal_9982 ;
    wire signal_9983 ;
    wire signal_9984 ;
    wire signal_9985 ;
    wire signal_9986 ;
    wire signal_9987 ;
    wire signal_9988 ;
    wire signal_9989 ;
    wire signal_9990 ;
    wire signal_9991 ;
    wire signal_9992 ;
    wire signal_9993 ;
    wire signal_9994 ;
    wire signal_9995 ;
    wire signal_9996 ;
    wire signal_9997 ;
    wire signal_9998 ;
    wire signal_9999 ;
    wire signal_10000 ;
    wire signal_10001 ;
    wire signal_10002 ;
    wire signal_10003 ;
    wire signal_10004 ;
    wire signal_10005 ;
    wire signal_10006 ;
    wire signal_10007 ;
    wire signal_10008 ;
    wire signal_10009 ;
    wire signal_10010 ;
    wire signal_10011 ;
    wire signal_10012 ;
    wire signal_10013 ;
    wire signal_10014 ;
    wire signal_10015 ;
    wire signal_10016 ;
    wire signal_10017 ;
    wire signal_10018 ;
    wire signal_10019 ;
    wire signal_10020 ;
    wire signal_10021 ;
    wire signal_10022 ;
    wire signal_10023 ;
    wire signal_10024 ;
    wire signal_10025 ;
    wire signal_10026 ;
    wire signal_10027 ;
    wire signal_10028 ;
    wire signal_10029 ;
    wire signal_10030 ;
    wire signal_10031 ;
    wire signal_10032 ;
    wire signal_10033 ;
    wire signal_10034 ;
    wire signal_10035 ;
    wire signal_10036 ;
    wire signal_10037 ;
    wire signal_10038 ;
    wire signal_10039 ;
    wire signal_10040 ;
    wire signal_10041 ;
    wire signal_10042 ;
    wire signal_10043 ;
    wire signal_10044 ;
    wire signal_10045 ;
    wire signal_10046 ;
    wire signal_10047 ;
    wire signal_10048 ;
    wire signal_10049 ;
    wire signal_10050 ;
    wire signal_10051 ;
    wire signal_10052 ;
    wire signal_10053 ;
    wire signal_10054 ;
    wire signal_10055 ;
    wire signal_10056 ;
    wire signal_10057 ;
    wire signal_10058 ;
    wire signal_10059 ;
    wire signal_10060 ;
    wire signal_10061 ;
    wire signal_10062 ;
    wire signal_10063 ;
    wire signal_10064 ;
    wire signal_10065 ;
    wire signal_10066 ;
    wire signal_10067 ;
    wire signal_10068 ;
    wire signal_10069 ;
    wire signal_10070 ;
    wire signal_10071 ;
    wire signal_10072 ;
    wire signal_10073 ;
    wire signal_10074 ;
    wire signal_10075 ;
    wire signal_10076 ;
    wire signal_10077 ;
    wire signal_10078 ;
    wire signal_10079 ;
    wire signal_10080 ;
    wire signal_10081 ;
    wire signal_10082 ;
    wire signal_10083 ;
    wire signal_10084 ;
    wire signal_10085 ;
    wire signal_10086 ;
    wire signal_10087 ;
    wire signal_10088 ;
    wire signal_10089 ;
    wire signal_10090 ;
    wire signal_10091 ;
    wire signal_10092 ;
    wire signal_10093 ;
    wire signal_10094 ;
    wire signal_10095 ;
    wire signal_10096 ;
    wire signal_10097 ;
    wire signal_10098 ;
    wire signal_10099 ;
    wire signal_10100 ;
    wire signal_10101 ;
    wire signal_10102 ;
    wire signal_10103 ;
    wire signal_10104 ;
    wire signal_10105 ;
    wire signal_10106 ;
    wire signal_10107 ;
    wire signal_10108 ;
    wire signal_10109 ;
    wire signal_10110 ;
    wire signal_10111 ;
    wire signal_10112 ;
    wire signal_10113 ;
    wire signal_10114 ;
    wire signal_10115 ;
    wire signal_10116 ;
    wire signal_10117 ;
    wire signal_10118 ;
    wire signal_10119 ;
    wire signal_10120 ;
    wire signal_10121 ;
    wire signal_10122 ;
    wire signal_10123 ;
    wire signal_10124 ;
    wire signal_10125 ;
    wire signal_10126 ;
    wire signal_10127 ;
    wire signal_10128 ;
    wire signal_10129 ;
    wire signal_10130 ;
    wire signal_10131 ;
    wire signal_10132 ;
    wire signal_10133 ;
    wire signal_10134 ;
    wire signal_10135 ;
    wire signal_10136 ;
    wire signal_10137 ;
    wire signal_10138 ;
    wire signal_10139 ;
    wire signal_10140 ;
    wire signal_10141 ;
    wire signal_10142 ;
    wire signal_10143 ;
    wire signal_10144 ;
    wire signal_10145 ;
    wire signal_10146 ;
    wire signal_10147 ;
    wire signal_10148 ;
    wire signal_10149 ;
    wire signal_10150 ;
    wire signal_10151 ;
    wire signal_10152 ;
    wire signal_10153 ;
    wire signal_10154 ;
    wire signal_10155 ;
    wire signal_10156 ;
    wire signal_10157 ;
    wire signal_10158 ;
    wire signal_10159 ;
    wire signal_10160 ;
    wire signal_10161 ;
    wire signal_10162 ;
    wire signal_10163 ;
    wire signal_10164 ;
    wire signal_10165 ;
    wire signal_10166 ;
    wire signal_10167 ;
    wire signal_10168 ;
    wire signal_10169 ;
    wire signal_10170 ;
    wire signal_10171 ;
    wire signal_10172 ;
    wire signal_10173 ;
    wire signal_10174 ;
    wire signal_10175 ;
    wire signal_10176 ;
    wire signal_10177 ;
    wire signal_10178 ;
    wire signal_10179 ;
    wire signal_10180 ;
    wire signal_10181 ;
    wire signal_10182 ;
    wire signal_10183 ;
    wire signal_10184 ;
    wire signal_10185 ;
    wire signal_10186 ;
    wire signal_10187 ;
    wire signal_10188 ;
    wire signal_10189 ;
    wire signal_10190 ;
    wire signal_10191 ;
    wire signal_10192 ;
    wire signal_10193 ;
    wire signal_10194 ;
    wire signal_10195 ;
    wire signal_10196 ;
    wire signal_10197 ;
    wire signal_10198 ;
    wire signal_10199 ;
    wire signal_10200 ;
    wire signal_10201 ;
    wire signal_10202 ;
    wire signal_10203 ;
    wire signal_10204 ;
    wire signal_10205 ;
    wire signal_10206 ;
    wire signal_10207 ;
    wire signal_10208 ;
    wire signal_10209 ;
    wire signal_10210 ;
    wire signal_10211 ;
    wire signal_10212 ;
    wire signal_10213 ;
    wire signal_10214 ;
    wire signal_10215 ;
    wire signal_10216 ;
    wire signal_10217 ;
    wire signal_10218 ;
    wire signal_10219 ;
    wire signal_10220 ;
    wire signal_10221 ;
    wire signal_10222 ;
    wire signal_10223 ;
    wire signal_10224 ;
    wire signal_10225 ;
    wire signal_10226 ;
    wire signal_10227 ;
    wire signal_10228 ;
    wire signal_10229 ;
    wire signal_10230 ;
    wire signal_10231 ;
    wire signal_10232 ;
    wire signal_10233 ;
    wire signal_10234 ;
    wire signal_10235 ;
    wire signal_10236 ;
    wire signal_10237 ;
    wire signal_10238 ;
    wire signal_10239 ;
    wire signal_10240 ;
    wire signal_10241 ;
    wire signal_10242 ;
    wire signal_10243 ;
    wire signal_10244 ;
    wire signal_10245 ;
    wire signal_10246 ;
    wire signal_10247 ;
    wire signal_10248 ;
    wire signal_10249 ;
    wire signal_10250 ;
    wire signal_10251 ;
    wire signal_10252 ;
    wire signal_10253 ;
    wire signal_10254 ;
    wire signal_10255 ;
    wire signal_10256 ;
    wire signal_10257 ;
    wire signal_10258 ;
    wire signal_10259 ;
    wire signal_10260 ;
    wire signal_10261 ;
    wire signal_10262 ;
    wire signal_10263 ;
    wire signal_10264 ;
    wire signal_10265 ;
    wire signal_10266 ;
    wire signal_10267 ;
    wire signal_10268 ;
    wire signal_10269 ;
    wire signal_10270 ;
    wire signal_10271 ;
    wire signal_10272 ;
    wire signal_10273 ;
    wire signal_10274 ;
    wire signal_10275 ;
    wire signal_10276 ;
    wire signal_10277 ;
    wire signal_10278 ;
    wire signal_10279 ;
    wire signal_10280 ;
    wire signal_10281 ;
    wire signal_10282 ;
    wire signal_10283 ;
    wire signal_10284 ;
    wire signal_10285 ;
    wire signal_10286 ;
    wire signal_10287 ;
    wire signal_10288 ;
    wire signal_10289 ;
    wire signal_10290 ;
    wire signal_10291 ;
    wire signal_10292 ;
    wire signal_10293 ;
    wire signal_10294 ;
    wire signal_10295 ;
    wire signal_10296 ;
    wire signal_10297 ;
    wire signal_10298 ;
    wire signal_10299 ;
    wire signal_10300 ;
    wire signal_10301 ;
    wire signal_10302 ;
    wire signal_10303 ;
    wire signal_10304 ;
    wire signal_10305 ;
    wire signal_10306 ;
    wire signal_10307 ;
    wire signal_10308 ;
    wire signal_10309 ;
    wire signal_10310 ;
    wire signal_10311 ;
    wire signal_10312 ;
    wire signal_10313 ;
    wire signal_10314 ;
    wire signal_10315 ;
    wire signal_10316 ;
    wire signal_10317 ;
    wire signal_10318 ;
    wire signal_10319 ;
    wire signal_10320 ;
    wire signal_10321 ;
    wire signal_10322 ;
    wire signal_10323 ;
    wire signal_10324 ;
    wire signal_10325 ;
    wire signal_10326 ;
    wire signal_10327 ;
    wire signal_10328 ;
    wire signal_10329 ;
    wire signal_10330 ;
    wire signal_10331 ;
    wire signal_10332 ;
    wire signal_10333 ;
    wire signal_10334 ;
    wire signal_10335 ;
    wire signal_10336 ;
    wire signal_10337 ;
    wire signal_10338 ;
    wire signal_10339 ;
    wire signal_10340 ;
    wire signal_10341 ;
    wire signal_10342 ;
    wire signal_10343 ;
    wire signal_10344 ;
    wire signal_10345 ;
    wire signal_10346 ;
    wire signal_10347 ;
    wire signal_10348 ;
    wire signal_10349 ;
    wire signal_10350 ;
    wire signal_10351 ;
    wire signal_10352 ;
    wire signal_10353 ;
    wire signal_10354 ;
    wire signal_10355 ;
    wire signal_10356 ;
    wire signal_10357 ;
    wire signal_10358 ;
    wire signal_10359 ;
    wire signal_10360 ;
    wire signal_10361 ;
    wire signal_10362 ;
    wire signal_10363 ;
    wire signal_10364 ;
    wire signal_10365 ;
    wire signal_10366 ;
    wire signal_10367 ;
    wire signal_10368 ;
    wire signal_10369 ;
    wire signal_10370 ;
    wire signal_10371 ;
    wire signal_10372 ;
    wire signal_10373 ;
    wire signal_10374 ;
    wire signal_10375 ;
    wire signal_10376 ;
    wire signal_10377 ;
    wire signal_10378 ;
    wire signal_10379 ;
    wire signal_10380 ;
    wire signal_10381 ;
    wire signal_10382 ;
    wire signal_10383 ;
    wire signal_10384 ;
    wire signal_10385 ;
    wire signal_10386 ;
    wire signal_10387 ;
    wire signal_10388 ;
    wire signal_10389 ;
    wire signal_10390 ;
    wire signal_10391 ;
    wire signal_10392 ;
    wire signal_10393 ;
    wire signal_10394 ;
    wire signal_10395 ;
    wire signal_10396 ;
    wire signal_10397 ;
    wire signal_10398 ;
    wire signal_10399 ;
    wire signal_10400 ;
    wire signal_10401 ;
    wire signal_10402 ;
    wire signal_10403 ;
    wire signal_10404 ;
    wire signal_10405 ;
    wire signal_10406 ;
    wire signal_10407 ;
    wire signal_10408 ;
    wire signal_10409 ;
    wire signal_10410 ;
    wire signal_10411 ;
    wire signal_10412 ;
    wire signal_10413 ;
    wire signal_10414 ;
    wire signal_10415 ;
    wire signal_10416 ;
    wire signal_10417 ;
    wire signal_10418 ;
    wire signal_10419 ;
    wire signal_10420 ;
    wire signal_10421 ;
    wire signal_10422 ;
    wire signal_10423 ;
    wire signal_10424 ;
    wire signal_10425 ;
    wire signal_10426 ;
    wire signal_10427 ;
    wire signal_10428 ;
    wire signal_10429 ;
    wire signal_10430 ;
    wire signal_10431 ;
    wire signal_10432 ;
    wire signal_10433 ;
    wire signal_10434 ;
    wire signal_10435 ;
    wire signal_10436 ;
    wire signal_10437 ;
    wire signal_10438 ;
    wire signal_10439 ;
    wire signal_10440 ;
    wire signal_10441 ;
    wire signal_10442 ;
    wire signal_10443 ;
    wire signal_10444 ;
    wire signal_10445 ;
    wire signal_10446 ;
    wire signal_10447 ;
    wire signal_10448 ;
    wire signal_10449 ;
    wire signal_10450 ;
    wire signal_10451 ;
    wire signal_10452 ;
    wire signal_10453 ;
    wire signal_10454 ;
    wire signal_10455 ;
    wire signal_10457 ;
    wire signal_10459 ;
    wire signal_10461 ;
    wire signal_10463 ;
    wire signal_10465 ;
    wire signal_10467 ;
    wire signal_10469 ;
    wire signal_10471 ;
    wire signal_10473 ;
    wire signal_10475 ;
    wire signal_10477 ;
    wire signal_10479 ;
    wire signal_10481 ;
    wire signal_10483 ;
    wire signal_10485 ;
    wire signal_10486 ;
    wire signal_10487 ;
    wire signal_10488 ;
    wire signal_10489 ;
    wire signal_10490 ;
    wire signal_10491 ;
    wire signal_10492 ;
    wire signal_10493 ;
    wire signal_10494 ;
    wire signal_10495 ;
    wire signal_10496 ;
    wire signal_10497 ;
    wire signal_10498 ;
    wire signal_10499 ;
    wire signal_10500 ;
    wire signal_10501 ;
    wire signal_10502 ;
    wire signal_10503 ;
    wire signal_10504 ;
    wire signal_10505 ;
    wire signal_10506 ;
    wire signal_10507 ;
    wire signal_10508 ;
    wire signal_10509 ;
    wire signal_10510 ;
    wire signal_10511 ;
    wire signal_10512 ;
    wire signal_10513 ;
    wire signal_10514 ;
    wire signal_10515 ;
    wire signal_10516 ;
    wire signal_10517 ;
    wire signal_10518 ;
    wire signal_10519 ;
    wire signal_10520 ;
    wire signal_10521 ;
    wire signal_10522 ;
    wire signal_10523 ;
    wire signal_10524 ;
    wire signal_10525 ;
    wire signal_10526 ;
    wire signal_10527 ;
    wire signal_10528 ;
    wire signal_10529 ;
    wire signal_10530 ;
    wire signal_10531 ;
    wire signal_10532 ;
    wire signal_10533 ;
    wire signal_10534 ;
    wire signal_10535 ;
    wire signal_10536 ;
    wire signal_10537 ;
    wire signal_10538 ;
    wire signal_10539 ;
    wire signal_10540 ;
    wire signal_10541 ;
    wire signal_10542 ;
    wire signal_10543 ;
    wire signal_10544 ;
    wire signal_10545 ;
    wire signal_10546 ;
    wire signal_10547 ;
    wire signal_10548 ;
    wire signal_10549 ;
    wire signal_10550 ;
    wire signal_10551 ;
    wire signal_10552 ;
    wire signal_10553 ;
    wire signal_10554 ;
    wire signal_10555 ;
    wire signal_10556 ;
    wire signal_10557 ;
    wire signal_10558 ;
    wire signal_10559 ;
    wire signal_10560 ;
    wire signal_10561 ;
    wire signal_10562 ;
    wire signal_10563 ;
    wire signal_10564 ;
    wire signal_10565 ;
    wire signal_10566 ;
    wire signal_10567 ;
    wire signal_10568 ;
    wire signal_10569 ;
    wire signal_10570 ;
    wire signal_10571 ;
    wire signal_10572 ;
    wire signal_10573 ;
    wire signal_10574 ;
    wire signal_10575 ;
    wire signal_10576 ;
    wire signal_10577 ;
    wire signal_10578 ;
    wire signal_10579 ;
    wire signal_10580 ;
    wire signal_10581 ;
    wire signal_10582 ;
    wire signal_10583 ;
    wire signal_10584 ;
    wire signal_10585 ;
    wire signal_10586 ;
    wire signal_10587 ;
    wire signal_10588 ;
    wire signal_10589 ;
    wire signal_10590 ;
    wire signal_10591 ;
    wire signal_10592 ;
    wire signal_10593 ;
    wire signal_10594 ;
    wire signal_10595 ;
    wire signal_10596 ;
    wire signal_10597 ;
    wire signal_10598 ;
    wire signal_10599 ;
    wire signal_10600 ;
    wire signal_10601 ;
    wire signal_10602 ;
    wire signal_10603 ;
    wire signal_10604 ;
    wire signal_10605 ;
    wire signal_10606 ;
    wire signal_10607 ;
    wire signal_10608 ;
    wire signal_10609 ;
    wire signal_10610 ;
    wire signal_10611 ;
    wire signal_10612 ;
    wire signal_10613 ;
    wire signal_10614 ;
    wire signal_10615 ;
    wire signal_10616 ;
    wire signal_10617 ;
    wire signal_10618 ;
    wire signal_10619 ;
    wire signal_10620 ;
    wire signal_10621 ;
    wire signal_10622 ;
    wire signal_10623 ;
    wire signal_10624 ;
    wire signal_10625 ;
    wire signal_10626 ;
    wire signal_10627 ;
    wire signal_10628 ;
    wire signal_10629 ;
    wire signal_10630 ;
    wire signal_10631 ;
    wire signal_10632 ;
    wire signal_10633 ;
    wire signal_10634 ;
    wire signal_10635 ;
    wire signal_10636 ;
    wire signal_10637 ;
    wire signal_10638 ;
    wire signal_10639 ;
    wire signal_10640 ;
    wire signal_10641 ;
    wire signal_10642 ;
    wire signal_10643 ;
    wire signal_10644 ;
    wire signal_10645 ;
    wire signal_10646 ;
    wire signal_10647 ;
    wire signal_10648 ;
    wire signal_10649 ;
    wire signal_10650 ;
    wire signal_10651 ;
    wire signal_10652 ;
    wire signal_10653 ;
    wire signal_10654 ;
    wire signal_10655 ;
    wire signal_10656 ;
    wire signal_10657 ;
    wire signal_10658 ;
    wire signal_10659 ;
    wire signal_10660 ;
    wire signal_10661 ;
    wire signal_10662 ;
    wire signal_10663 ;
    wire signal_10664 ;
    wire signal_10665 ;
    wire signal_10666 ;
    wire signal_10667 ;
    wire signal_10668 ;
    wire signal_10669 ;
    wire signal_10670 ;
    wire signal_10671 ;
    wire signal_10672 ;
    wire signal_10673 ;
    wire signal_10674 ;
    wire signal_10675 ;
    wire signal_10676 ;
    wire signal_10677 ;
    wire signal_10678 ;
    wire signal_10679 ;
    wire signal_10680 ;
    wire signal_10681 ;
    wire signal_10682 ;
    wire signal_10683 ;
    wire signal_10684 ;
    wire signal_10685 ;
    wire signal_10686 ;
    wire signal_10687 ;
    wire signal_10688 ;
    wire signal_10689 ;
    wire signal_10690 ;
    wire signal_10691 ;
    wire signal_10692 ;
    wire signal_10693 ;
    wire signal_10694 ;
    wire signal_10695 ;
    wire signal_10696 ;
    wire signal_10697 ;
    wire signal_10698 ;
    wire signal_10699 ;
    wire signal_10700 ;
    wire signal_10701 ;
    wire signal_10702 ;
    wire signal_10703 ;
    wire signal_10704 ;
    wire signal_10705 ;
    wire signal_10707 ;
    wire signal_10709 ;
    wire signal_10711 ;
    wire signal_10713 ;
    wire signal_10715 ;
    wire signal_10717 ;
    wire signal_10719 ;
    wire signal_10721 ;
    wire signal_10723 ;
    wire signal_10725 ;
    wire signal_10727 ;
    wire signal_10729 ;
    wire signal_10731 ;
    wire signal_10733 ;
    wire signal_10735 ;
    wire signal_10737 ;
    wire signal_10739 ;
    wire signal_10741 ;
    wire signal_10743 ;
    wire signal_10745 ;
    wire signal_10747 ;
    wire signal_10749 ;
    wire signal_10751 ;
    wire signal_10753 ;
    wire signal_10755 ;
    wire signal_10757 ;
    wire signal_10759 ;
    wire signal_10761 ;
    wire signal_10763 ;
    wire signal_10764 ;
    wire signal_10765 ;
    wire signal_10766 ;
    wire signal_10767 ;
    wire signal_10768 ;
    wire signal_10769 ;
    wire signal_10770 ;
    wire signal_10771 ;
    wire signal_10772 ;
    wire signal_10773 ;
    wire signal_10774 ;
    wire signal_10775 ;
    wire signal_10776 ;
    wire signal_10777 ;
    wire signal_10778 ;
    wire signal_10779 ;
    wire signal_10780 ;
    wire signal_10781 ;
    wire signal_10782 ;
    wire signal_10783 ;
    wire signal_10784 ;
    wire signal_10785 ;
    wire signal_10786 ;
    wire signal_10787 ;
    wire signal_10788 ;
    wire signal_10789 ;
    wire signal_10790 ;
    wire signal_10791 ;
    wire signal_10792 ;
    wire signal_10793 ;
    wire signal_10794 ;
    wire signal_10795 ;
    wire signal_10796 ;
    wire signal_10797 ;
    wire signal_10798 ;
    wire signal_10799 ;
    wire signal_10800 ;
    wire signal_10801 ;
    wire signal_10802 ;
    wire signal_10803 ;
    wire signal_10804 ;
    wire signal_10805 ;
    wire signal_10806 ;
    wire signal_10807 ;
    wire signal_10808 ;
    wire signal_10809 ;
    wire signal_10810 ;
    wire signal_10811 ;
    wire signal_10812 ;
    wire signal_10813 ;
    wire signal_10814 ;
    wire signal_10815 ;
    wire signal_10816 ;
    wire signal_10817 ;
    wire signal_10818 ;
    wire signal_10819 ;
    wire signal_10820 ;
    wire signal_10821 ;
    wire signal_10822 ;
    wire signal_10823 ;
    wire signal_10824 ;
    wire signal_10825 ;
    wire signal_10826 ;
    wire signal_10827 ;
    wire signal_10828 ;
    wire signal_10829 ;
    wire signal_10830 ;
    wire signal_10831 ;
    wire signal_10832 ;
    wire signal_10833 ;
    wire signal_10834 ;
    wire signal_10835 ;
    wire signal_10836 ;
    wire signal_10837 ;
    wire signal_10838 ;
    wire signal_10839 ;
    wire signal_10840 ;
    wire signal_10841 ;
    wire signal_10842 ;
    wire signal_10843 ;
    wire signal_10844 ;
    wire signal_10845 ;
    wire signal_10846 ;
    wire signal_10847 ;
    wire signal_10848 ;
    wire signal_10849 ;
    wire signal_10850 ;
    wire signal_10851 ;
    wire signal_10852 ;
    wire signal_10853 ;
    wire signal_10854 ;
    wire signal_10855 ;
    wire signal_10856 ;
    wire signal_10857 ;
    wire signal_10858 ;
    wire signal_10859 ;
    wire signal_10860 ;
    wire signal_10861 ;
    wire signal_10862 ;
    wire signal_10863 ;
    wire signal_10864 ;
    wire signal_10865 ;
    wire signal_10866 ;
    wire signal_10867 ;
    wire signal_10868 ;
    wire signal_10869 ;
    wire signal_10870 ;
    wire signal_10871 ;
    wire signal_10872 ;
    wire signal_10873 ;
    wire signal_10874 ;
    wire signal_10875 ;
    wire signal_10876 ;
    wire signal_10877 ;
    wire signal_10878 ;
    wire signal_10879 ;
    wire signal_10880 ;
    wire signal_10881 ;
    wire signal_10882 ;
    wire signal_10883 ;
    wire signal_10884 ;
    wire signal_10885 ;
    wire signal_10886 ;
    wire signal_10887 ;
    wire signal_10888 ;
    wire signal_10889 ;
    wire signal_10890 ;
    wire signal_10891 ;
    wire signal_10892 ;
    wire signal_10893 ;
    wire signal_10894 ;
    wire signal_10895 ;
    wire signal_10896 ;
    wire signal_10897 ;
    wire signal_10898 ;
    wire signal_10899 ;
    wire signal_10900 ;
    wire signal_10901 ;
    wire signal_10902 ;
    wire signal_10903 ;
    wire signal_10904 ;
    wire signal_10905 ;
    wire signal_10906 ;
    wire signal_10907 ;
    wire signal_10908 ;
    wire signal_10909 ;
    wire signal_10910 ;
    wire signal_10911 ;
    wire signal_10912 ;
    wire signal_10913 ;
    wire signal_10914 ;
    wire signal_10915 ;
    wire signal_10916 ;
    wire signal_10917 ;
    wire signal_10918 ;
    wire signal_10919 ;
    wire signal_10920 ;
    wire signal_10921 ;
    wire signal_10922 ;
    wire signal_10923 ;
    wire signal_10924 ;
    wire signal_10925 ;
    wire signal_10926 ;
    wire signal_10927 ;
    wire signal_10928 ;
    wire signal_10929 ;
    wire signal_10930 ;
    wire signal_10931 ;
    wire signal_10932 ;
    wire signal_10933 ;
    wire signal_10934 ;
    wire signal_10935 ;
    wire signal_10937 ;
    wire signal_10939 ;
    wire signal_10941 ;
    wire signal_10943 ;
    wire signal_10945 ;
    wire signal_10947 ;
    wire signal_10949 ;
    wire signal_10951 ;
    wire signal_10953 ;
    wire signal_10955 ;
    wire signal_10957 ;
    wire signal_10959 ;
    wire signal_10961 ;
    wire signal_10963 ;
    wire signal_10965 ;
    wire signal_10967 ;
    wire signal_10969 ;
    wire signal_10971 ;
    wire signal_10973 ;
    wire signal_10975 ;
    wire signal_10977 ;
    wire signal_10979 ;
    wire signal_10981 ;
    wire signal_10983 ;
    wire signal_10985 ;
    wire signal_10987 ;
    wire signal_10989 ;
    wire signal_10991 ;
    wire signal_10993 ;
    wire signal_10995 ;
    wire signal_10997 ;
    wire signal_10999 ;
    wire signal_11000 ;
    wire signal_11001 ;
    wire signal_11002 ;
    wire signal_11003 ;
    wire signal_11004 ;
    wire signal_11005 ;
    wire signal_11006 ;
    wire signal_11007 ;
    wire signal_11008 ;
    wire signal_11009 ;
    wire signal_11010 ;
    wire signal_11011 ;
    wire signal_11012 ;
    wire signal_11013 ;
    wire signal_11014 ;
    wire signal_11015 ;
    wire signal_11016 ;
    wire signal_11017 ;
    wire signal_11018 ;
    wire signal_11019 ;
    wire signal_11020 ;
    wire signal_11021 ;
    wire signal_11022 ;
    wire signal_11023 ;
    wire signal_11024 ;
    wire signal_11025 ;
    wire signal_11026 ;
    wire signal_11027 ;
    wire signal_11028 ;
    wire signal_11029 ;
    wire signal_11030 ;
    wire signal_11031 ;
    wire signal_11032 ;
    wire signal_11033 ;
    wire signal_11034 ;
    wire signal_11035 ;
    wire signal_11036 ;
    wire signal_11037 ;
    wire signal_11038 ;
    wire signal_11039 ;
    wire signal_11040 ;
    wire signal_11041 ;
    wire signal_11042 ;
    wire signal_11043 ;
    wire signal_11044 ;
    wire signal_11045 ;
    wire signal_11046 ;
    wire signal_11047 ;
    wire signal_11048 ;
    wire signal_11049 ;
    wire signal_11050 ;
    wire signal_11051 ;
    wire signal_11052 ;
    wire signal_11053 ;
    wire signal_11054 ;
    wire signal_11055 ;
    wire signal_11056 ;
    wire signal_11057 ;
    wire signal_11058 ;
    wire signal_11059 ;
    wire signal_11060 ;
    wire signal_11061 ;
    wire signal_11062 ;
    wire signal_11063 ;
    wire signal_11064 ;
    wire signal_11065 ;
    wire signal_11066 ;
    wire signal_11067 ;
    wire signal_11068 ;
    wire signal_11069 ;
    wire signal_11070 ;
    wire signal_11071 ;
    wire signal_11072 ;
    wire signal_11073 ;
    wire signal_11074 ;
    wire signal_11075 ;
    wire signal_11076 ;
    wire signal_11077 ;
    wire signal_11078 ;
    wire signal_11079 ;
    wire signal_11080 ;
    wire signal_11081 ;
    wire signal_11082 ;
    wire signal_11083 ;
    wire signal_11084 ;
    wire signal_11085 ;
    wire signal_11086 ;
    wire signal_11087 ;
    wire signal_11088 ;
    wire signal_11089 ;
    wire signal_11090 ;
    wire signal_11091 ;
    wire signal_11092 ;
    wire signal_11093 ;
    wire signal_11094 ;
    wire signal_11095 ;
    wire signal_11096 ;
    wire signal_11097 ;
    wire signal_11098 ;
    wire signal_11099 ;
    wire signal_11100 ;
    wire signal_11101 ;
    wire signal_11102 ;
    wire signal_11103 ;
    wire signal_11104 ;
    wire signal_11105 ;
    wire signal_11106 ;
    wire signal_11107 ;
    wire signal_11108 ;
    wire signal_11109 ;
    wire signal_11110 ;
    wire signal_11111 ;
    wire signal_11112 ;
    wire signal_11113 ;
    wire signal_11114 ;
    wire signal_11115 ;
    wire signal_11116 ;
    wire signal_11117 ;
    wire signal_11118 ;
    wire signal_11119 ;
    wire signal_11120 ;
    wire signal_11121 ;
    wire signal_11122 ;
    wire signal_11123 ;
    wire signal_11124 ;
    wire signal_11125 ;
    wire signal_11126 ;
    wire signal_11127 ;
    wire signal_11128 ;
    wire signal_11129 ;
    wire signal_11130 ;
    wire signal_11131 ;
    wire signal_11132 ;
    wire signal_11133 ;
    wire signal_11134 ;
    wire signal_11135 ;
    wire signal_11136 ;
    wire signal_11137 ;
    wire signal_11138 ;
    wire signal_11139 ;
    wire signal_11140 ;
    wire signal_11141 ;
    wire signal_11142 ;
    wire signal_11143 ;
    wire signal_11144 ;
    wire signal_11145 ;
    wire signal_11146 ;
    wire signal_11147 ;
    wire signal_11148 ;
    wire signal_11149 ;
    wire signal_11150 ;
    wire signal_11151 ;
    wire signal_11152 ;
    wire signal_11153 ;
    wire signal_11154 ;
    wire signal_11155 ;
    wire signal_11156 ;
    wire signal_11157 ;
    wire signal_11158 ;
    wire signal_11159 ;
    wire signal_11160 ;
    wire signal_11161 ;
    wire signal_11162 ;
    wire signal_11163 ;
    wire signal_11164 ;
    wire signal_11165 ;
    wire signal_11166 ;
    wire signal_11167 ;
    wire signal_11168 ;
    wire signal_11169 ;
    wire signal_11170 ;
    wire signal_11171 ;
    wire signal_11172 ;
    wire signal_11173 ;
    wire signal_11174 ;
    wire signal_11175 ;
    wire signal_11176 ;
    wire signal_11177 ;
    wire signal_11178 ;
    wire signal_11179 ;
    wire signal_11180 ;
    wire signal_11181 ;
    wire signal_11182 ;
    wire signal_11183 ;
    wire signal_11184 ;
    wire signal_11185 ;
    wire signal_11186 ;
    wire signal_11187 ;
    wire signal_11188 ;
    wire signal_11189 ;
    wire signal_11190 ;
    wire signal_11191 ;
    wire signal_11192 ;
    wire signal_11193 ;
    wire signal_11194 ;
    wire signal_11195 ;
    wire signal_11196 ;
    wire signal_11197 ;
    wire signal_11198 ;
    wire signal_11199 ;
    wire signal_11200 ;
    wire signal_11202 ;
    wire signal_11204 ;
    wire signal_11206 ;
    wire signal_11208 ;
    wire signal_11210 ;
    wire signal_11212 ;
    wire signal_11214 ;
    wire signal_11216 ;
    wire signal_11218 ;
    wire signal_11220 ;
    wire signal_11222 ;
    wire signal_11224 ;
    wire signal_11226 ;
    wire signal_11228 ;
    wire signal_11230 ;
    wire signal_11232 ;
    wire signal_11234 ;
    wire signal_11236 ;
    wire signal_11238 ;
    wire signal_11240 ;
    wire signal_11242 ;
    wire signal_11244 ;
    wire signal_11246 ;
    wire signal_11248 ;
    wire signal_11250 ;
    wire signal_11252 ;
    wire signal_11254 ;
    wire signal_11256 ;
    wire signal_11258 ;
    wire signal_11260 ;
    wire signal_11262 ;
    wire signal_11264 ;
    wire signal_11265 ;
    wire signal_11266 ;
    wire signal_11267 ;
    wire signal_11268 ;
    wire signal_11269 ;
    wire signal_11270 ;
    wire signal_11271 ;
    wire signal_11272 ;
    wire signal_11273 ;
    wire signal_11274 ;
    wire signal_11275 ;
    wire signal_11276 ;
    wire signal_11277 ;
    wire signal_11278 ;
    wire signal_11279 ;
    wire signal_11280 ;
    wire signal_11281 ;
    wire signal_11282 ;
    wire signal_11283 ;
    wire signal_11284 ;
    wire signal_11285 ;
    wire signal_11286 ;
    wire signal_11287 ;
    wire signal_11288 ;
    wire signal_11289 ;
    wire signal_11290 ;
    wire signal_11291 ;
    wire signal_11292 ;
    wire signal_11293 ;
    wire signal_11294 ;
    wire signal_11295 ;
    wire signal_11296 ;
    wire signal_11297 ;
    wire signal_11298 ;
    wire signal_11299 ;
    wire signal_11300 ;
    wire signal_11301 ;
    wire signal_11302 ;
    wire signal_11303 ;
    wire signal_11304 ;
    wire signal_11305 ;
    wire signal_11306 ;
    wire signal_11307 ;
    wire signal_11308 ;
    wire signal_11309 ;
    wire signal_11310 ;
    wire signal_11311 ;
    wire signal_11312 ;
    wire signal_11313 ;
    wire signal_11314 ;
    wire signal_11315 ;
    wire signal_11316 ;
    wire signal_11317 ;
    wire signal_11318 ;
    wire signal_11319 ;
    wire signal_11320 ;
    wire signal_11321 ;
    wire signal_11322 ;
    wire signal_11323 ;
    wire signal_11324 ;
    wire signal_11325 ;
    wire signal_11326 ;
    wire signal_11327 ;
    wire signal_11328 ;
    wire signal_11329 ;
    wire signal_11330 ;
    wire signal_11331 ;
    wire signal_11332 ;
    wire signal_11333 ;
    wire signal_11334 ;
    wire signal_11335 ;
    wire signal_11336 ;
    wire signal_11337 ;
    wire signal_11338 ;
    wire signal_11339 ;
    wire signal_11340 ;
    wire signal_11341 ;
    wire signal_11342 ;
    wire signal_11343 ;
    wire signal_11344 ;
    wire signal_11345 ;
    wire signal_11346 ;
    wire signal_11347 ;
    wire signal_11348 ;
    wire signal_11349 ;
    wire signal_11350 ;
    wire signal_11351 ;
    wire signal_11352 ;
    wire signal_11353 ;
    wire signal_11354 ;
    wire signal_11355 ;
    wire signal_11356 ;
    wire signal_11357 ;
    wire signal_11358 ;
    wire signal_11359 ;
    wire signal_11360 ;
    wire signal_11361 ;
    wire signal_11362 ;
    wire signal_11363 ;
    wire signal_11364 ;
    wire signal_11365 ;
    wire signal_11366 ;
    wire signal_11367 ;
    wire signal_11368 ;
    wire signal_11369 ;
    wire signal_11370 ;
    wire signal_11371 ;
    wire signal_11372 ;
    wire signal_11373 ;
    wire signal_11374 ;
    wire signal_11375 ;
    wire signal_11376 ;
    wire signal_11377 ;
    wire signal_11378 ;
    wire signal_11379 ;
    wire signal_11380 ;
    wire signal_11381 ;
    wire signal_11382 ;
    wire signal_11383 ;
    wire signal_11384 ;
    wire signal_11385 ;
    wire signal_11386 ;
    wire signal_11387 ;
    wire signal_11388 ;
    wire signal_11389 ;
    wire signal_11390 ;
    wire signal_11391 ;
    wire signal_11392 ;
    wire signal_11393 ;
    wire signal_11394 ;
    wire signal_11395 ;
    wire signal_11396 ;
    wire signal_11397 ;
    wire signal_11398 ;
    wire signal_11399 ;
    wire signal_11400 ;
    wire signal_11401 ;
    wire signal_11402 ;
    wire signal_11403 ;
    wire signal_11404 ;
    wire signal_11405 ;
    wire signal_11406 ;
    wire signal_11407 ;
    wire signal_11408 ;
    wire signal_11409 ;
    wire signal_11410 ;
    wire signal_11411 ;
    wire signal_11412 ;
    wire signal_11413 ;
    wire signal_11414 ;
    wire signal_11415 ;
    wire signal_11416 ;
    wire signal_11417 ;
    wire signal_11418 ;
    wire signal_11419 ;
    wire signal_11420 ;
    wire signal_11421 ;
    wire signal_11422 ;
    wire signal_11423 ;
    wire signal_11424 ;
    wire signal_11425 ;
    wire signal_11426 ;
    wire signal_11427 ;
    wire signal_11428 ;
    wire signal_11429 ;
    wire signal_11430 ;
    wire signal_11431 ;
    wire signal_11432 ;
    wire signal_11433 ;
    wire signal_11434 ;
    wire signal_11435 ;
    wire signal_11436 ;
    wire signal_11437 ;
    wire signal_11438 ;
    wire signal_11439 ;
    wire signal_11440 ;
    wire signal_11441 ;
    wire signal_11442 ;
    wire signal_11443 ;
    wire signal_11444 ;
    wire signal_11445 ;
    wire signal_11446 ;
    wire signal_11447 ;
    wire signal_11448 ;
    wire signal_11449 ;
    wire signal_11450 ;
    wire signal_11451 ;
    wire signal_11452 ;
    wire signal_11453 ;
    wire signal_11454 ;
    wire signal_11455 ;
    wire signal_11456 ;
    wire signal_11457 ;
    wire signal_11459 ;
    wire signal_11461 ;
    wire signal_11463 ;
    wire signal_11465 ;
    wire signal_11467 ;
    wire signal_11469 ;
    wire signal_11471 ;
    wire signal_11473 ;
    wire signal_11475 ;
    wire signal_11477 ;
    wire signal_11479 ;
    wire signal_11481 ;
    wire signal_11483 ;
    wire signal_11485 ;
    wire signal_11487 ;
    wire signal_11489 ;
    wire signal_11491 ;
    wire signal_11493 ;
    wire signal_11495 ;
    wire signal_11497 ;
    wire signal_11499 ;
    wire signal_11501 ;
    wire signal_11503 ;
    wire signal_11505 ;
    wire signal_11507 ;
    wire signal_11509 ;
    wire signal_11511 ;
    wire signal_11513 ;
    wire signal_11515 ;
    wire signal_11517 ;
    wire signal_11519 ;
    wire signal_11521 ;
    wire signal_11523 ;
    wire signal_11525 ;
    wire signal_11527 ;
    wire signal_11529 ;
    wire signal_11531 ;
    wire signal_11533 ;
    wire signal_11535 ;
    wire signal_11537 ;
    wire signal_11539 ;
    wire signal_11541 ;
    wire signal_11543 ;
    wire signal_11545 ;
    wire signal_11547 ;
    wire signal_11549 ;
    wire signal_11551 ;
    wire signal_11553 ;
    wire signal_11555 ;
    wire signal_11556 ;
    wire signal_11557 ;
    wire signal_11558 ;
    wire signal_11559 ;
    wire signal_11560 ;
    wire signal_11561 ;
    wire signal_11562 ;
    wire signal_11563 ;
    wire signal_11564 ;
    wire signal_11565 ;
    wire signal_11566 ;
    wire signal_11567 ;
    wire signal_11568 ;
    wire signal_11569 ;
    wire signal_11570 ;
    wire signal_11571 ;
    wire signal_11572 ;
    wire signal_11573 ;
    wire signal_11574 ;
    wire signal_11575 ;
    wire signal_11576 ;
    wire signal_11577 ;
    wire signal_11578 ;
    wire signal_11579 ;
    wire signal_11580 ;
    wire signal_11581 ;
    wire signal_11582 ;
    wire signal_11583 ;
    wire signal_11584 ;
    wire signal_11585 ;
    wire signal_11586 ;
    wire signal_11587 ;
    wire signal_11588 ;
    wire signal_11589 ;
    wire signal_11590 ;
    wire signal_11592 ;
    wire signal_11594 ;
    wire signal_11596 ;
    wire signal_11598 ;
    wire signal_11600 ;
    wire signal_11602 ;
    wire signal_11604 ;
    wire signal_11606 ;
    wire signal_11608 ;
    wire signal_11610 ;
    wire signal_11612 ;
    wire signal_11614 ;
    wire signal_11616 ;
    wire signal_11618 ;
    wire signal_11620 ;
    wire signal_11622 ;
    wire signal_11624 ;
    wire signal_11626 ;
    wire signal_11628 ;
    wire signal_11630 ;
    wire signal_11632 ;
    wire signal_11634 ;
    wire signal_11636 ;
    wire signal_11638 ;
    wire signal_11640 ;
    wire signal_11642 ;
    wire signal_11644 ;
    wire signal_11646 ;
    wire signal_11648 ;
    wire signal_11650 ;
    wire signal_11652 ;
    wire signal_11654 ;
    wire signal_11656 ;
    wire signal_11658 ;
    wire signal_11660 ;
    wire signal_11662 ;
    wire signal_11664 ;
    wire signal_11666 ;
    wire signal_11668 ;
    wire signal_11670 ;
    wire signal_11672 ;
    wire signal_11674 ;
    wire signal_11676 ;
    wire signal_11678 ;
    wire signal_11680 ;
    wire signal_11682 ;
    wire signal_11684 ;
    wire signal_11686 ;
    wire signal_11688 ;
    wire signal_11690 ;
    wire signal_11692 ;
    wire signal_11694 ;
    wire signal_11696 ;
    wire signal_11698 ;
    wire signal_11700 ;
    wire signal_11702 ;
    wire signal_11704 ;
    wire signal_11706 ;
    wire signal_11708 ;
    wire signal_11710 ;
    wire signal_11712 ;
    wire signal_11714 ;
    wire signal_11716 ;
    wire signal_11718 ;
    wire signal_11720 ;
    wire signal_11722 ;
    wire signal_11724 ;
    wire signal_11726 ;
    wire signal_11728 ;
    wire signal_11730 ;
    wire signal_11732 ;
    wire signal_11734 ;
    wire signal_11736 ;
    wire signal_11738 ;
    wire signal_11740 ;
    wire signal_11742 ;
    wire signal_11744 ;
    wire signal_11746 ;
    wire signal_11748 ;
    wire signal_11750 ;
    wire signal_11752 ;
    wire signal_11754 ;
    wire signal_11756 ;
    wire signal_11758 ;
    wire signal_11760 ;
    wire signal_11762 ;
    wire signal_11764 ;
    wire signal_11766 ;
    wire signal_11768 ;
    wire signal_11770 ;
    wire signal_11772 ;
    wire signal_11774 ;
    wire signal_11776 ;
    wire signal_11778 ;
    wire signal_11780 ;
    wire signal_11782 ;
    wire signal_11784 ;
    wire signal_11786 ;
    wire signal_11788 ;
    wire signal_12469 ;
    wire signal_12470 ;
    wire signal_12471 ;
    wire signal_12472 ;
    wire signal_12473 ;
    wire signal_12474 ;
    wire signal_12475 ;
    wire signal_12476 ;
    wire signal_12477 ;
    wire signal_12478 ;
    wire signal_12479 ;
    wire signal_12480 ;
    wire signal_12481 ;
    wire signal_12482 ;
    wire signal_12483 ;
    wire signal_12484 ;
    wire signal_12485 ;
    wire signal_12486 ;
    wire signal_12487 ;
    wire signal_12488 ;
    wire signal_12489 ;
    wire signal_12490 ;
    wire signal_12491 ;
    wire signal_12492 ;
    wire signal_12493 ;
    wire signal_12494 ;
    wire signal_12495 ;
    wire signal_12496 ;
    wire signal_12497 ;
    wire signal_12498 ;
    wire signal_12499 ;
    wire signal_12500 ;
    wire signal_12501 ;
    wire signal_12502 ;
    wire signal_12503 ;
    wire signal_12504 ;
    wire signal_12505 ;
    wire signal_12506 ;
    wire signal_12507 ;
    wire signal_12508 ;
    wire signal_12509 ;
    wire signal_12510 ;
    wire signal_12511 ;
    wire signal_12512 ;
    wire signal_12513 ;
    wire signal_12514 ;
    wire signal_12515 ;
    wire signal_12516 ;
    wire signal_12517 ;
    wire signal_12518 ;
    wire signal_12519 ;
    wire signal_12520 ;
    wire signal_12521 ;
    wire signal_12522 ;
    wire signal_12523 ;
    wire signal_12524 ;
    wire signal_12525 ;
    wire signal_12526 ;
    wire signal_12527 ;
    wire signal_12528 ;
    wire signal_12529 ;
    wire signal_12530 ;
    wire signal_12531 ;
    wire signal_12532 ;
    wire signal_12533 ;
    wire signal_12534 ;
    wire signal_12535 ;
    wire signal_12536 ;
    wire signal_12537 ;
    wire signal_12538 ;
    wire signal_12539 ;
    wire signal_12540 ;
    wire signal_12541 ;
    wire signal_12542 ;
    wire signal_12543 ;
    wire signal_12544 ;
    wire signal_12545 ;
    wire signal_12546 ;
    wire signal_12547 ;
    wire signal_12548 ;
    wire signal_12549 ;
    wire signal_12550 ;
    wire signal_12551 ;
    wire signal_12552 ;
    wire signal_12553 ;
    wire signal_12554 ;
    wire signal_12555 ;
    wire signal_12556 ;
    wire signal_12557 ;
    wire signal_12558 ;
    wire signal_12559 ;
    wire signal_12560 ;
    wire signal_12561 ;
    wire signal_12562 ;
    wire signal_12563 ;
    wire signal_12564 ;
    wire signal_12565 ;
    wire signal_12566 ;
    wire signal_12567 ;
    wire signal_12568 ;
    wire signal_12569 ;
    wire signal_12570 ;
    wire signal_12571 ;
    wire signal_12572 ;
    wire signal_12573 ;
    wire signal_12574 ;
    wire signal_12575 ;
    wire signal_12576 ;
    wire signal_12577 ;
    wire signal_12578 ;
    wire signal_12579 ;
    wire signal_12580 ;
    wire signal_12581 ;
    wire signal_12582 ;
    wire signal_12583 ;
    wire signal_12584 ;
    wire signal_12585 ;
    wire signal_12586 ;
    wire signal_12587 ;
    wire signal_12588 ;
    wire signal_12589 ;
    wire signal_12590 ;
    wire signal_12591 ;
    wire signal_12592 ;
    wire signal_12593 ;
    wire signal_12594 ;
    wire signal_12595 ;
    wire signal_12596 ;
    wire signal_12597 ;
    wire signal_12598 ;
    wire signal_12599 ;
    wire signal_12600 ;
    wire signal_12601 ;
    wire signal_12602 ;
    wire signal_12603 ;
    wire signal_12604 ;
    wire signal_12605 ;
    wire signal_12606 ;
    wire signal_12607 ;
    wire signal_12608 ;
    wire signal_12609 ;
    wire signal_12610 ;
    wire signal_12611 ;
    wire signal_12612 ;
    wire signal_12613 ;
    wire signal_12614 ;
    wire signal_12615 ;
    wire signal_12616 ;
    wire signal_12617 ;
    wire signal_12618 ;
    wire signal_12619 ;
    wire signal_12620 ;
    wire signal_12621 ;
    wire signal_12622 ;
    wire signal_12623 ;
    wire signal_12624 ;
    wire signal_12625 ;
    wire signal_12626 ;
    wire signal_12627 ;
    wire signal_12628 ;
    wire signal_12629 ;
    wire signal_12630 ;
    wire signal_12631 ;
    wire signal_12632 ;
    wire signal_12633 ;
    wire signal_12634 ;
    wire signal_12635 ;
    wire signal_12636 ;
    wire signal_12637 ;
    wire signal_12638 ;
    wire signal_12639 ;
    wire signal_12640 ;
    wire signal_12641 ;
    wire signal_12642 ;
    wire signal_12643 ;
    wire signal_12644 ;
    wire signal_12645 ;
    wire signal_12646 ;
    wire signal_12647 ;
    wire signal_12648 ;
    wire signal_12649 ;
    wire signal_12650 ;
    wire signal_12651 ;
    wire signal_12652 ;
    wire signal_12653 ;
    wire signal_12654 ;
    wire signal_12655 ;
    wire signal_12656 ;
    wire signal_12657 ;
    wire signal_12658 ;
    wire signal_12659 ;
    wire signal_12660 ;
    wire signal_12661 ;
    wire signal_12662 ;
    wire signal_12663 ;
    wire signal_12664 ;
    wire signal_12665 ;
    wire signal_12666 ;
    wire signal_12667 ;
    wire signal_12668 ;
    wire signal_12669 ;
    wire signal_12670 ;
    wire signal_12671 ;
    wire signal_12672 ;
    wire signal_12673 ;
    wire signal_12674 ;
    wire signal_12675 ;
    wire signal_12676 ;
    wire signal_12677 ;
    wire signal_12678 ;
    wire signal_12679 ;
    wire signal_12680 ;
    wire signal_12681 ;
    wire signal_12682 ;
    wire signal_12683 ;
    wire signal_12684 ;
    wire signal_12685 ;
    wire signal_12686 ;
    wire signal_12687 ;
    wire signal_12688 ;
    wire signal_12689 ;
    wire signal_12690 ;
    wire signal_12691 ;
    wire signal_12692 ;
    wire signal_12693 ;
    wire signal_12694 ;
    wire signal_12695 ;
    wire signal_12696 ;
    wire signal_12697 ;
    wire signal_12698 ;
    wire signal_12699 ;
    wire signal_12700 ;
    wire signal_12701 ;
    wire signal_12702 ;
    wire signal_12703 ;
    wire signal_12704 ;
    wire signal_12705 ;
    wire signal_12706 ;
    wire signal_12707 ;
    wire signal_12708 ;
    wire signal_12709 ;
    wire signal_12710 ;
    wire signal_12711 ;
    wire signal_12712 ;
    wire signal_12713 ;
    wire signal_12714 ;
    wire signal_12715 ;
    wire signal_12716 ;
    wire signal_12717 ;
    wire signal_12718 ;
    wire signal_12719 ;
    wire signal_12720 ;
    wire signal_12721 ;
    wire signal_12722 ;
    wire signal_12723 ;
    wire signal_12724 ;
    wire signal_12725 ;
    wire signal_12726 ;
    wire signal_12727 ;
    wire signal_12728 ;
    wire signal_12729 ;
    wire signal_12730 ;
    wire signal_12731 ;
    wire signal_12732 ;
    wire signal_12733 ;
    wire signal_12734 ;
    wire signal_12735 ;
    wire signal_12736 ;
    wire signal_12737 ;
    wire signal_12738 ;
    wire signal_12739 ;
    wire signal_12740 ;
    wire signal_12741 ;
    wire signal_12742 ;
    wire signal_12743 ;
    wire signal_12744 ;
    wire signal_12745 ;
    wire signal_12746 ;
    wire signal_12747 ;
    wire signal_12748 ;
    wire signal_12749 ;
    wire signal_12750 ;
    wire signal_12751 ;
    wire signal_12752 ;
    wire signal_12753 ;
    wire signal_12754 ;
    wire signal_12755 ;
    wire signal_12756 ;
    wire signal_12757 ;
    wire signal_12758 ;
    wire signal_12759 ;
    wire signal_12760 ;
    wire signal_12761 ;
    wire signal_12762 ;
    wire signal_12763 ;
    wire signal_12764 ;
    wire signal_12765 ;
    wire signal_12766 ;
    wire signal_12767 ;
    wire signal_12768 ;
    wire signal_12769 ;
    wire signal_12770 ;
    wire signal_12771 ;
    wire signal_12772 ;
    wire signal_12773 ;
    wire signal_12774 ;
    wire signal_12775 ;
    wire signal_12776 ;
    wire signal_12777 ;
    wire signal_12778 ;
    wire signal_12779 ;
    wire signal_12780 ;
    wire signal_12781 ;
    wire signal_12782 ;
    wire signal_12783 ;
    wire signal_12784 ;
    wire signal_12785 ;
    wire signal_12786 ;
    wire signal_12787 ;
    wire signal_12788 ;
    wire signal_12789 ;
    wire signal_12790 ;
    wire signal_12791 ;
    wire signal_12792 ;
    wire signal_12793 ;
    wire signal_12794 ;
    wire signal_12795 ;
    wire signal_12796 ;
    wire signal_12797 ;
    wire signal_12798 ;
    wire signal_12799 ;
    wire signal_12800 ;
    wire signal_12801 ;
    wire signal_12802 ;
    wire signal_12803 ;
    wire signal_12804 ;
    wire signal_12805 ;
    wire signal_12806 ;
    wire signal_12807 ;
    wire signal_12808 ;
    wire signal_12809 ;
    wire signal_12810 ;
    wire signal_12811 ;
    wire signal_12812 ;
    wire signal_12813 ;
    wire signal_12814 ;
    wire signal_12815 ;
    wire signal_12816 ;
    wire signal_12817 ;
    wire signal_12818 ;
    wire signal_12819 ;
    wire signal_12820 ;
    wire signal_12821 ;
    wire signal_12822 ;
    wire signal_12823 ;
    wire signal_12824 ;
    wire signal_12825 ;
    wire signal_12826 ;
    wire signal_12827 ;
    wire signal_12828 ;
    wire signal_12829 ;
    wire signal_12830 ;
    wire signal_12831 ;
    wire signal_12832 ;
    wire signal_12833 ;
    wire signal_12834 ;
    wire signal_12835 ;
    wire signal_12836 ;
    wire signal_12837 ;
    wire signal_12838 ;
    wire signal_12839 ;
    wire signal_12840 ;
    wire signal_12841 ;
    wire signal_12842 ;
    wire signal_12843 ;
    wire signal_12844 ;
    wire signal_12845 ;
    wire signal_12846 ;
    wire signal_12847 ;
    wire signal_12848 ;
    wire signal_12849 ;
    wire signal_12850 ;
    wire signal_12851 ;
    wire signal_12852 ;
    wire signal_12853 ;
    wire signal_12854 ;
    wire signal_12855 ;
    wire signal_12856 ;
    wire signal_12857 ;
    wire signal_12858 ;
    wire signal_12859 ;
    wire signal_12860 ;
    wire signal_12861 ;
    wire signal_12862 ;
    wire signal_12863 ;
    wire signal_12864 ;
    wire signal_12865 ;
    wire signal_12866 ;
    wire signal_12867 ;
    wire signal_12868 ;
    wire signal_12869 ;
    wire signal_12870 ;
    wire signal_12871 ;
    wire signal_12872 ;
    wire signal_12873 ;
    wire signal_12874 ;
    wire signal_12875 ;
    wire signal_12876 ;
    wire signal_12877 ;
    wire signal_12878 ;
    wire signal_12879 ;
    wire signal_12880 ;
    wire signal_12881 ;
    wire signal_12882 ;
    wire signal_12883 ;
    wire signal_12884 ;
    wire signal_12885 ;
    wire signal_12886 ;
    wire signal_12887 ;
    wire signal_12888 ;
    wire signal_12889 ;
    wire signal_12890 ;
    wire signal_12891 ;
    wire signal_12892 ;
    wire signal_12893 ;
    wire signal_12894 ;
    wire signal_12895 ;
    wire signal_12896 ;
    wire signal_12897 ;
    wire signal_12898 ;
    wire signal_12899 ;
    wire signal_12900 ;
    wire signal_12901 ;
    wire signal_12902 ;
    wire signal_12903 ;
    wire signal_12904 ;
    wire signal_12905 ;
    wire signal_12906 ;
    wire signal_12907 ;
    wire signal_12908 ;
    wire signal_12909 ;
    wire signal_12910 ;
    wire signal_12911 ;
    wire signal_12912 ;
    wire signal_12913 ;
    wire signal_12914 ;
    wire signal_12915 ;
    wire signal_12916 ;
    wire signal_12917 ;
    wire signal_12918 ;
    wire signal_12919 ;
    wire signal_12920 ;
    wire signal_12921 ;
    wire signal_12922 ;
    wire signal_12923 ;
    wire signal_12924 ;
    wire signal_12925 ;
    wire signal_12926 ;
    wire signal_12927 ;
    wire signal_12928 ;
    wire signal_12929 ;
    wire signal_12930 ;
    wire signal_12931 ;
    wire signal_12932 ;
    wire signal_12933 ;
    wire signal_12934 ;
    wire signal_12935 ;
    wire signal_12936 ;
    wire signal_12937 ;
    wire signal_12938 ;
    wire signal_12939 ;
    wire signal_12940 ;
    wire signal_12941 ;
    wire signal_12942 ;
    wire signal_12943 ;
    wire signal_12944 ;
    wire signal_12945 ;
    wire signal_12946 ;
    wire signal_12947 ;
    wire signal_12948 ;
    wire signal_12949 ;
    wire signal_12950 ;
    wire signal_12951 ;
    wire signal_12952 ;
    wire signal_12953 ;
    wire signal_12954 ;
    wire signal_12955 ;
    wire signal_12956 ;
    wire signal_12957 ;
    wire signal_12958 ;
    wire signal_12959 ;
    wire signal_12960 ;
    wire signal_12961 ;
    wire signal_12962 ;
    wire signal_12963 ;
    wire signal_12964 ;
    wire signal_12965 ;
    wire signal_12966 ;
    wire signal_12967 ;
    wire signal_12968 ;
    wire signal_12969 ;
    wire signal_12970 ;
    wire signal_12971 ;
    wire signal_12972 ;
    wire signal_12973 ;
    wire signal_12974 ;
    wire signal_12975 ;
    wire signal_12976 ;
    wire signal_12977 ;
    wire signal_12978 ;
    wire signal_12979 ;
    wire signal_12980 ;
    wire signal_12981 ;
    wire signal_12982 ;
    wire signal_12983 ;
    wire signal_12984 ;
    wire signal_12985 ;
    wire signal_12986 ;
    wire signal_12987 ;
    wire signal_12988 ;
    wire signal_12989 ;
    wire signal_12990 ;
    wire signal_12991 ;
    wire signal_12992 ;
    wire signal_12993 ;
    wire signal_12994 ;
    wire signal_12995 ;
    wire signal_12996 ;
    wire signal_12997 ;
    wire signal_12998 ;
    wire signal_12999 ;
    wire signal_13000 ;
    wire signal_13001 ;
    wire signal_13002 ;
    wire signal_13003 ;
    wire signal_13004 ;
    wire signal_13005 ;
    wire signal_13006 ;
    wire signal_13007 ;
    wire signal_13008 ;
    wire signal_13009 ;
    wire signal_13010 ;
    wire signal_13011 ;
    wire signal_13012 ;
    wire signal_13013 ;
    wire signal_13014 ;
    wire signal_13015 ;
    wire signal_13016 ;
    wire signal_13017 ;
    wire signal_13018 ;
    wire signal_13019 ;
    wire signal_13020 ;
    wire signal_13021 ;
    wire signal_13022 ;
    wire signal_13023 ;
    wire signal_13024 ;
    wire signal_13025 ;
    wire signal_13026 ;
    wire signal_13027 ;
    wire signal_13028 ;
    wire signal_13029 ;
    wire signal_13030 ;
    wire signal_13031 ;
    wire signal_13032 ;
    wire signal_13033 ;
    wire signal_13034 ;
    wire signal_13035 ;
    wire signal_13036 ;
    wire signal_13037 ;
    wire signal_13038 ;
    wire signal_13039 ;
    wire signal_13040 ;
    wire signal_13041 ;
    wire signal_13042 ;
    wire signal_13043 ;
    wire signal_13044 ;
    wire signal_13045 ;
    wire signal_13046 ;
    wire signal_13047 ;
    wire signal_13048 ;
    wire signal_13049 ;
    wire signal_13050 ;
    wire signal_13051 ;
    wire signal_13052 ;
    wire signal_13053 ;
    wire signal_13054 ;
    wire signal_13055 ;
    wire signal_13056 ;
    wire signal_13057 ;
    wire signal_13058 ;
    wire signal_13059 ;
    wire signal_13060 ;
    wire signal_13061 ;
    wire signal_13062 ;
    wire signal_13063 ;
    wire signal_13064 ;
    wire signal_13065 ;
    wire signal_13066 ;
    wire signal_13067 ;
    wire signal_13068 ;
    wire signal_13069 ;
    wire signal_13070 ;
    wire signal_13071 ;
    wire signal_13072 ;
    wire signal_13073 ;
    wire signal_13074 ;
    wire signal_13075 ;
    wire signal_13076 ;
    wire signal_13077 ;
    wire signal_13078 ;
    wire signal_13079 ;
    wire signal_13080 ;
    wire signal_13081 ;
    wire signal_13082 ;
    wire signal_13083 ;
    wire signal_13084 ;
    wire signal_13085 ;
    wire signal_13086 ;
    wire signal_13087 ;
    wire signal_13088 ;
    wire signal_13089 ;
    wire signal_13090 ;
    wire signal_13091 ;
    wire signal_13092 ;
    wire signal_13093 ;
    wire signal_13094 ;
    wire signal_13095 ;
    wire signal_13096 ;
    wire signal_13097 ;
    wire signal_13098 ;
    wire signal_13099 ;
    wire signal_13100 ;
    wire signal_13101 ;
    wire signal_13102 ;
    wire signal_13103 ;
    wire signal_13104 ;
    wire signal_13105 ;
    wire signal_13106 ;
    wire signal_13107 ;
    wire signal_13108 ;
    wire signal_13109 ;
    wire signal_13110 ;
    wire signal_13111 ;
    wire signal_13112 ;
    wire signal_13113 ;
    wire signal_13114 ;
    wire signal_13115 ;
    wire signal_13116 ;
    wire signal_13117 ;
    wire signal_13118 ;
    wire signal_13119 ;
    wire signal_13120 ;
    wire signal_13121 ;
    wire signal_13122 ;
    wire signal_13123 ;
    wire signal_13124 ;
    wire signal_13125 ;
    wire signal_13126 ;
    wire signal_13127 ;
    wire signal_13128 ;
    wire signal_13129 ;
    wire signal_13130 ;
    wire signal_13131 ;
    wire signal_13132 ;
    wire signal_13133 ;
    wire signal_13134 ;
    wire signal_13135 ;
    wire signal_13136 ;
    wire signal_13137 ;
    wire signal_13138 ;
    wire signal_13139 ;
    wire signal_13140 ;
    wire signal_13141 ;
    wire signal_13142 ;
    wire signal_13143 ;
    wire signal_13144 ;
    wire signal_13145 ;
    wire signal_13146 ;
    wire signal_13147 ;
    wire signal_13148 ;
    wire signal_13149 ;
    wire signal_13150 ;
    wire signal_13151 ;
    wire signal_13152 ;
    wire signal_13153 ;
    wire signal_13154 ;
    wire signal_13155 ;
    wire signal_13156 ;
    wire signal_13157 ;
    wire signal_13158 ;
    wire signal_13159 ;
    wire signal_13160 ;
    wire signal_13161 ;
    wire signal_13162 ;
    wire signal_13163 ;
    wire signal_13164 ;
    wire signal_13165 ;
    wire signal_13166 ;
    wire signal_13167 ;
    wire signal_13168 ;
    wire signal_13169 ;
    wire signal_13170 ;
    wire signal_13171 ;
    wire signal_13172 ;
    wire signal_13173 ;
    wire signal_13174 ;
    wire signal_13175 ;
    wire signal_13176 ;
    wire signal_13177 ;
    wire signal_13178 ;
    wire signal_13179 ;
    wire signal_13180 ;
    wire signal_13181 ;
    wire signal_13182 ;
    wire signal_13183 ;
    wire signal_13184 ;
    wire signal_13185 ;
    wire signal_13186 ;
    wire signal_13187 ;
    wire signal_13188 ;
    wire signal_13189 ;
    wire signal_13190 ;
    wire signal_13191 ;
    wire signal_13192 ;
    wire signal_13193 ;
    wire signal_13194 ;
    wire signal_13195 ;
    wire signal_13196 ;
    wire signal_13197 ;
    wire signal_13198 ;
    wire signal_13199 ;
    wire signal_13200 ;
    wire signal_13201 ;
    wire signal_13202 ;
    wire signal_13203 ;
    wire signal_13204 ;
    wire signal_13205 ;
    wire signal_13206 ;
    wire signal_13207 ;
    wire signal_13208 ;
    wire signal_13209 ;
    wire signal_13210 ;
    wire signal_13211 ;
    wire signal_13212 ;
    wire signal_13213 ;
    wire signal_13214 ;
    wire signal_13215 ;
    wire signal_13216 ;
    wire signal_13217 ;
    wire signal_13218 ;
    wire signal_13219 ;
    wire signal_13220 ;
    wire signal_13221 ;
    wire signal_13222 ;
    wire signal_13223 ;
    wire signal_13224 ;
    wire signal_13225 ;
    wire signal_13226 ;
    wire signal_13227 ;
    wire signal_13228 ;
    wire signal_13229 ;
    wire signal_13230 ;
    wire signal_13231 ;
    wire signal_13232 ;
    wire signal_13233 ;
    wire signal_13234 ;
    wire signal_13235 ;
    wire signal_13236 ;
    wire signal_13237 ;
    wire signal_13238 ;
    wire signal_13239 ;
    wire signal_13240 ;
    wire signal_13241 ;
    wire signal_13242 ;
    wire signal_13243 ;
    wire signal_13244 ;
    wire signal_13245 ;
    wire signal_13246 ;
    wire signal_13247 ;
    wire signal_13248 ;
    wire signal_13249 ;
    wire signal_13250 ;
    wire signal_13251 ;
    wire signal_13252 ;
    wire signal_13253 ;
    wire signal_13254 ;
    wire signal_13255 ;
    wire signal_13256 ;
    wire signal_13257 ;
    wire signal_13258 ;
    wire signal_13259 ;
    wire signal_13260 ;
    wire signal_13261 ;
    wire signal_13262 ;
    wire signal_13263 ;
    wire signal_13264 ;
    wire signal_13265 ;
    wire signal_13266 ;
    wire signal_13267 ;
    wire signal_13268 ;
    wire signal_13269 ;
    wire signal_13270 ;
    wire signal_13271 ;
    wire signal_13272 ;
    wire signal_13273 ;
    wire signal_13274 ;
    wire signal_13275 ;
    wire signal_13276 ;
    wire signal_13277 ;
    wire signal_13278 ;
    wire signal_13279 ;
    wire signal_13280 ;
    wire signal_13281 ;
    wire signal_13282 ;
    wire signal_13283 ;
    wire signal_13284 ;
    wire signal_13285 ;
    wire signal_13286 ;
    wire signal_13287 ;
    wire signal_13288 ;
    wire signal_13289 ;
    wire signal_13290 ;
    wire signal_13291 ;
    wire signal_13292 ;
    wire signal_13293 ;
    wire signal_13294 ;
    wire signal_13295 ;
    wire signal_13296 ;
    wire signal_13297 ;
    wire signal_13298 ;
    wire signal_13299 ;
    wire signal_13300 ;
    wire signal_13301 ;
    wire signal_13302 ;
    wire signal_13303 ;
    wire signal_13304 ;
    wire signal_13305 ;
    wire signal_13306 ;
    wire signal_13307 ;
    wire signal_13308 ;
    wire signal_13309 ;
    wire signal_13310 ;
    wire signal_13311 ;
    wire signal_13312 ;
    wire signal_13313 ;
    wire signal_13314 ;
    wire signal_13315 ;
    wire signal_13316 ;
    wire signal_13317 ;
    wire signal_13318 ;
    wire signal_13319 ;
    wire signal_13320 ;
    wire signal_13321 ;
    wire signal_13322 ;
    wire signal_13323 ;
    wire signal_13324 ;
    wire signal_13325 ;
    wire signal_13326 ;
    wire signal_13327 ;
    wire signal_13328 ;
    wire signal_13329 ;
    wire signal_13330 ;
    wire signal_13331 ;
    wire signal_13332 ;
    wire signal_13333 ;
    wire signal_13334 ;
    wire signal_13335 ;
    wire signal_13336 ;
    wire signal_13337 ;
    wire signal_13338 ;
    wire signal_13339 ;
    wire signal_13340 ;
    wire signal_13341 ;
    wire signal_13342 ;
    wire signal_13343 ;
    wire signal_13344 ;
    wire signal_13345 ;
    wire signal_13346 ;
    wire signal_13347 ;
    wire signal_13348 ;
    wire signal_13349 ;
    wire signal_13350 ;
    wire signal_13351 ;
    wire signal_13352 ;
    wire signal_13353 ;
    wire signal_13354 ;
    wire signal_13355 ;
    wire signal_13356 ;
    wire signal_13357 ;
    wire signal_13358 ;
    wire signal_13359 ;
    wire signal_13360 ;
    wire signal_13361 ;
    wire signal_13362 ;
    wire signal_13363 ;
    wire signal_13364 ;
    wire signal_13365 ;
    wire signal_13366 ;
    wire signal_13367 ;
    wire signal_13368 ;
    wire signal_13369 ;
    wire signal_13370 ;
    wire signal_13371 ;
    wire signal_13372 ;
    wire signal_13373 ;
    wire signal_13374 ;
    wire signal_13375 ;
    wire signal_13376 ;
    wire signal_13377 ;
    wire signal_13378 ;
    wire signal_13379 ;
    wire signal_13380 ;
    wire signal_13381 ;
    wire signal_13382 ;
    wire signal_13383 ;
    wire signal_13384 ;
    wire signal_13385 ;
    wire signal_13386 ;
    wire signal_13387 ;
    wire signal_13388 ;
    wire signal_13389 ;
    wire signal_13390 ;
    wire signal_13391 ;
    wire signal_13392 ;
    wire signal_13393 ;
    wire signal_13394 ;
    wire signal_13395 ;
    wire signal_13396 ;
    wire signal_13397 ;
    wire signal_13398 ;
    wire signal_13399 ;
    wire signal_13400 ;
    wire signal_13401 ;
    wire signal_13402 ;
    wire signal_13403 ;
    wire signal_13404 ;
    wire signal_13405 ;
    wire signal_13406 ;
    wire signal_13407 ;
    wire signal_13408 ;
    wire signal_13409 ;
    wire signal_13410 ;
    wire signal_13411 ;
    wire signal_13412 ;
    wire signal_13413 ;
    wire signal_13414 ;
    wire signal_13415 ;
    wire signal_13416 ;
    wire signal_13417 ;
    wire signal_13418 ;
    wire signal_13419 ;
    wire signal_13420 ;
    wire signal_13421 ;
    wire signal_13422 ;
    wire signal_13423 ;
    wire signal_13424 ;
    wire signal_13425 ;
    wire signal_13426 ;
    wire signal_13427 ;
    wire signal_13428 ;
    wire signal_13429 ;
    wire signal_13430 ;
    wire signal_13431 ;
    wire signal_13432 ;
    wire signal_13433 ;
    wire signal_13434 ;
    wire signal_13435 ;
    wire signal_13436 ;
    wire signal_13437 ;
    wire signal_13438 ;
    wire signal_13439 ;
    wire signal_13440 ;
    wire signal_13441 ;
    wire signal_13442 ;
    wire signal_13443 ;
    wire signal_13444 ;
    wire signal_13445 ;
    wire signal_13446 ;
    wire signal_13447 ;
    wire signal_13448 ;
    wire signal_13449 ;
    wire signal_13450 ;
    wire signal_13451 ;
    wire signal_13452 ;
    wire signal_13453 ;
    wire signal_13454 ;
    wire signal_13455 ;
    wire signal_13456 ;
    wire signal_13457 ;
    wire signal_13458 ;
    wire signal_13459 ;
    wire signal_13460 ;
    wire signal_13461 ;
    wire signal_13462 ;
    wire signal_13463 ;
    wire signal_13464 ;
    wire signal_13465 ;
    wire signal_13466 ;
    wire signal_13467 ;
    wire signal_13468 ;
    wire signal_13469 ;
    wire signal_13470 ;
    wire signal_13471 ;
    wire signal_13472 ;
    wire signal_13473 ;
    wire signal_13474 ;
    wire signal_13475 ;
    wire signal_13476 ;
    wire signal_13477 ;
    wire signal_13478 ;
    wire signal_13479 ;
    wire signal_13480 ;
    wire signal_13481 ;
    wire signal_13482 ;
    wire signal_13483 ;
    wire signal_13484 ;
    wire signal_13485 ;
    wire signal_13486 ;
    wire signal_13487 ;
    wire signal_13488 ;
    wire signal_13489 ;
    wire signal_13490 ;
    wire signal_13491 ;
    wire signal_13492 ;
    wire signal_13493 ;
    wire signal_13494 ;
    wire signal_13495 ;
    wire signal_13496 ;
    wire signal_13497 ;
    wire signal_13498 ;
    wire signal_13499 ;
    wire signal_13500 ;
    wire signal_13501 ;
    wire signal_13502 ;
    wire signal_13503 ;
    wire signal_13504 ;
    wire signal_13505 ;
    wire signal_13506 ;
    wire signal_13507 ;
    wire signal_13508 ;
    wire signal_13509 ;
    wire signal_13510 ;
    wire signal_13511 ;
    wire signal_13512 ;
    wire signal_13513 ;
    wire signal_13514 ;
    wire signal_13515 ;
    wire signal_13516 ;
    wire signal_13517 ;
    wire signal_13518 ;
    wire signal_13519 ;
    wire signal_13520 ;
    wire signal_13521 ;
    wire signal_13522 ;
    wire signal_13523 ;
    wire signal_13524 ;
    wire signal_13525 ;
    wire signal_13526 ;
    wire signal_13527 ;
    wire signal_13528 ;
    wire signal_13529 ;
    wire signal_13530 ;
    wire signal_13531 ;
    wire signal_13532 ;
    wire signal_13533 ;
    wire signal_13534 ;
    wire signal_13535 ;
    wire signal_13536 ;
    wire signal_13537 ;
    wire signal_13538 ;
    wire signal_13539 ;
    wire signal_13540 ;
    wire signal_13541 ;
    wire signal_13542 ;
    wire signal_13543 ;
    wire signal_13544 ;
    wire signal_13545 ;
    wire signal_13546 ;
    wire signal_13547 ;
    wire signal_13548 ;
    wire signal_13549 ;
    wire signal_13550 ;
    wire signal_13551 ;
    wire signal_13552 ;
    wire signal_13553 ;
    wire signal_13554 ;
    wire signal_13555 ;
    wire signal_13556 ;
    wire signal_13557 ;
    wire signal_13558 ;
    wire signal_13559 ;
    wire signal_13560 ;
    wire signal_13561 ;
    wire signal_13562 ;
    wire signal_13563 ;
    wire signal_13564 ;
    wire signal_13565 ;
    wire signal_13566 ;
    wire signal_13567 ;
    wire signal_13568 ;
    wire signal_13569 ;
    wire signal_13570 ;
    wire signal_13571 ;
    wire signal_13572 ;
    wire signal_13573 ;
    wire signal_13574 ;
    wire signal_13575 ;
    wire signal_13576 ;
    wire signal_13577 ;
    wire signal_13578 ;
    wire signal_13579 ;
    wire signal_13580 ;
    wire signal_13581 ;
    wire signal_13582 ;
    wire signal_13583 ;
    wire signal_13584 ;
    wire signal_13585 ;
    wire signal_13586 ;
    wire signal_13587 ;
    wire signal_13588 ;
    wire signal_13589 ;
    wire signal_13590 ;
    wire signal_13591 ;
    wire signal_13592 ;
    wire signal_13593 ;
    wire signal_13594 ;
    wire signal_13595 ;
    wire signal_13596 ;
    wire signal_13597 ;
    wire signal_13598 ;
    wire signal_13599 ;
    wire signal_13600 ;
    wire signal_13601 ;
    wire signal_13602 ;
    wire signal_13603 ;
    wire signal_13604 ;
    wire signal_13605 ;
    wire signal_13606 ;
    wire signal_13607 ;
    wire signal_13608 ;
    wire signal_13609 ;
    wire signal_13610 ;
    wire signal_13611 ;
    wire signal_13612 ;
    wire signal_13613 ;
    wire signal_13614 ;
    wire signal_13615 ;
    wire signal_13616 ;
    wire signal_13617 ;
    wire signal_13618 ;
    wire signal_13619 ;
    wire signal_13620 ;
    wire signal_13621 ;
    wire signal_13622 ;
    wire signal_13623 ;
    wire signal_13624 ;
    wire signal_13625 ;
    wire signal_13626 ;
    wire signal_13627 ;
    wire signal_13628 ;
    wire signal_13629 ;
    wire signal_13630 ;
    wire signal_13631 ;
    wire signal_13632 ;
    wire signal_13633 ;
    wire signal_13634 ;
    wire signal_13635 ;
    wire signal_13636 ;
    wire signal_13637 ;
    wire signal_13638 ;
    wire signal_13639 ;
    wire signal_13640 ;
    wire signal_13641 ;
    wire signal_13642 ;
    wire signal_13643 ;
    wire signal_13644 ;
    wire signal_13645 ;
    wire signal_13646 ;
    wire signal_13647 ;
    wire signal_13648 ;
    wire signal_13649 ;
    wire signal_13650 ;
    wire signal_13651 ;
    wire signal_13652 ;
    wire signal_13653 ;
    wire signal_13654 ;
    wire signal_13655 ;
    wire signal_13656 ;
    wire signal_13657 ;
    wire signal_13658 ;
    wire signal_13659 ;
    wire signal_13660 ;
    wire signal_13661 ;
    wire signal_13662 ;
    wire signal_13663 ;
    wire signal_13664 ;
    wire signal_13665 ;
    wire signal_13666 ;
    wire signal_13667 ;
    wire signal_13668 ;
    wire signal_13669 ;
    wire signal_13670 ;
    wire signal_13671 ;
    wire signal_13672 ;
    wire signal_13673 ;
    wire signal_13674 ;
    wire signal_13675 ;
    wire signal_13676 ;
    wire signal_13677 ;
    wire signal_13678 ;
    wire signal_13679 ;
    wire signal_13680 ;
    wire signal_13681 ;
    wire signal_13682 ;
    wire signal_13683 ;
    wire signal_13684 ;
    wire signal_13685 ;
    wire signal_13686 ;
    wire signal_13687 ;
    wire signal_13688 ;
    wire signal_13689 ;
    wire signal_13690 ;
    wire signal_13691 ;
    wire signal_13692 ;
    wire signal_13693 ;
    wire signal_13694 ;
    wire signal_13695 ;
    wire signal_13696 ;
    wire signal_13697 ;
    wire signal_13698 ;
    wire signal_13699 ;
    wire signal_13700 ;
    wire signal_13701 ;
    wire signal_13702 ;
    wire signal_13703 ;
    wire signal_13704 ;
    wire signal_13705 ;
    wire signal_13706 ;
    wire signal_13707 ;
    wire signal_13708 ;
    wire signal_13709 ;
    wire signal_13710 ;
    wire signal_13711 ;
    wire signal_13712 ;
    wire signal_13713 ;
    wire signal_13714 ;
    wire signal_13715 ;
    wire signal_13716 ;
    wire signal_13717 ;
    wire signal_13718 ;
    wire signal_13719 ;
    wire signal_13720 ;
    wire signal_13721 ;
    wire signal_13722 ;
    wire signal_13723 ;
    wire signal_13724 ;
    wire signal_13725 ;
    wire signal_13726 ;
    wire signal_13727 ;
    wire signal_13728 ;
    wire signal_13729 ;
    wire signal_13730 ;
    wire signal_13731 ;
    wire signal_13732 ;
    wire signal_13733 ;
    wire signal_13734 ;
    wire signal_13735 ;
    wire signal_13736 ;
    wire signal_13737 ;
    wire signal_13738 ;
    wire signal_13739 ;
    wire signal_13740 ;
    wire signal_13741 ;
    wire signal_13742 ;
    wire signal_13743 ;
    wire signal_13744 ;
    wire signal_13745 ;
    wire signal_13746 ;
    wire signal_13747 ;
    wire signal_13748 ;
    wire signal_13749 ;
    wire signal_13750 ;
    wire signal_13751 ;
    wire signal_13752 ;
    wire signal_13753 ;
    wire signal_13754 ;
    wire signal_13755 ;
    wire signal_13756 ;
    wire signal_13757 ;
    wire signal_13758 ;
    wire signal_13759 ;
    wire signal_13760 ;
    wire signal_13761 ;
    wire signal_13762 ;
    wire signal_13763 ;
    wire signal_13764 ;
    wire signal_13765 ;
    wire signal_13766 ;
    wire signal_13767 ;
    wire signal_13768 ;
    wire signal_13769 ;
    wire signal_13770 ;
    wire signal_13771 ;
    wire signal_13772 ;
    wire signal_13773 ;
    wire signal_13774 ;
    wire signal_13775 ;
    wire signal_13776 ;
    wire signal_13777 ;
    wire signal_13778 ;
    wire signal_13779 ;
    wire signal_13780 ;
    wire signal_13781 ;
    wire signal_13782 ;
    wire signal_13783 ;
    wire signal_13784 ;
    wire signal_13785 ;
    wire signal_13786 ;
    wire signal_13787 ;
    wire signal_13788 ;
    wire signal_13789 ;
    wire signal_13790 ;
    wire signal_13791 ;
    wire signal_13792 ;
    wire signal_13793 ;
    wire signal_13794 ;
    wire signal_13795 ;
    wire signal_13796 ;
    wire signal_13797 ;
    wire signal_13798 ;
    wire signal_13799 ;
    wire signal_13800 ;
    wire signal_13801 ;
    wire signal_13802 ;
    wire signal_13803 ;
    wire signal_13804 ;
    wire signal_13805 ;
    wire signal_13806 ;
    wire signal_13807 ;
    wire signal_13808 ;
    wire signal_13809 ;
    wire signal_13810 ;
    wire signal_13811 ;
    wire signal_13812 ;
    wire signal_13813 ;
    wire signal_13814 ;
    wire signal_13815 ;
    wire signal_13816 ;
    wire signal_13817 ;
    wire signal_13818 ;
    wire signal_13819 ;
    wire signal_13820 ;
    wire signal_13821 ;
    wire signal_13822 ;
    wire signal_13823 ;
    wire signal_13824 ;
    wire signal_13825 ;
    wire signal_13826 ;
    wire signal_13827 ;
    wire signal_13828 ;
    wire signal_13829 ;
    wire signal_13830 ;
    wire signal_13831 ;
    wire signal_13832 ;
    wire signal_13833 ;
    wire signal_13834 ;
    wire signal_13835 ;
    wire signal_13836 ;
    wire signal_13837 ;
    wire signal_13838 ;
    wire signal_13839 ;
    wire signal_13840 ;
    wire signal_13841 ;
    wire signal_13842 ;
    wire signal_13843 ;
    wire signal_13844 ;
    wire signal_13845 ;
    wire signal_13846 ;
    wire signal_13847 ;
    wire signal_13848 ;
    wire signal_13849 ;
    wire signal_13850 ;
    wire signal_13851 ;
    wire signal_13852 ;
    wire signal_13853 ;
    wire signal_13854 ;
    wire signal_13855 ;
    wire signal_13856 ;
    wire signal_13857 ;
    wire signal_13858 ;
    wire signal_13859 ;
    wire signal_13860 ;
    wire signal_13861 ;
    wire signal_13862 ;
    wire signal_13863 ;
    wire signal_13864 ;
    wire signal_13865 ;
    wire signal_13866 ;
    wire signal_13867 ;
    wire signal_13868 ;
    wire signal_13869 ;
    wire signal_13870 ;
    wire signal_13871 ;
    wire signal_13872 ;
    wire signal_13873 ;
    wire signal_13874 ;
    wire signal_13875 ;
    wire signal_13876 ;
    wire signal_13877 ;
    wire signal_13878 ;
    wire signal_13879 ;
    wire signal_13880 ;
    wire signal_13881 ;
    wire signal_13882 ;
    wire signal_13883 ;
    wire signal_13884 ;
    wire signal_13885 ;
    wire signal_13886 ;
    wire signal_13887 ;
    wire signal_13888 ;
    wire signal_13889 ;
    wire signal_13890 ;
    wire signal_13891 ;
    wire signal_13892 ;
    wire signal_13893 ;
    wire signal_13894 ;
    wire signal_13895 ;
    wire signal_13896 ;
    wire signal_13897 ;
    wire signal_13898 ;
    wire signal_13899 ;
    wire signal_13900 ;
    wire signal_13901 ;
    wire signal_13902 ;
    wire signal_13903 ;
    wire signal_13904 ;
    wire signal_13905 ;
    wire signal_13906 ;
    wire signal_13907 ;
    wire signal_13908 ;
    wire signal_13909 ;
    wire signal_13910 ;
    wire signal_13911 ;
    wire signal_13912 ;
    wire signal_13913 ;
    wire signal_13914 ;
    wire signal_13915 ;
    wire signal_13916 ;
    wire signal_13917 ;
    wire signal_13918 ;
    wire signal_13919 ;
    wire signal_13920 ;
    wire signal_13921 ;
    wire signal_13922 ;
    wire signal_13923 ;
    wire signal_13924 ;
    wire signal_13925 ;
    wire signal_13926 ;
    wire signal_13927 ;
    wire signal_13928 ;
    wire signal_13929 ;
    wire signal_13930 ;
    wire signal_13931 ;
    wire signal_13932 ;
    wire signal_13933 ;
    wire signal_13934 ;
    wire signal_13935 ;
    wire signal_13936 ;
    wire signal_13937 ;
    wire signal_13938 ;
    wire signal_13939 ;
    wire signal_13940 ;
    wire signal_13941 ;
    wire signal_13942 ;
    wire signal_13943 ;
    wire signal_13944 ;
    wire signal_13945 ;
    wire signal_13946 ;
    wire signal_13947 ;
    wire signal_13948 ;
    wire signal_13949 ;
    wire signal_13950 ;
    wire signal_13951 ;
    wire signal_13952 ;
    wire signal_13953 ;
    wire signal_13954 ;
    wire signal_13955 ;
    wire signal_13956 ;
    wire signal_13957 ;
    wire signal_13958 ;
    wire signal_13959 ;
    wire signal_13960 ;
    wire signal_13961 ;
    wire signal_13962 ;
    wire signal_13963 ;
    wire signal_13964 ;
    wire signal_13965 ;
    wire signal_13966 ;
    wire signal_13967 ;
    wire signal_13968 ;
    wire signal_13969 ;
    wire signal_13970 ;
    wire signal_13971 ;
    wire signal_13972 ;
    wire signal_13973 ;
    wire signal_13974 ;
    wire signal_13975 ;
    wire signal_13976 ;
    wire signal_13977 ;
    wire signal_13978 ;
    wire signal_13979 ;
    wire signal_13980 ;
    wire signal_13981 ;
    wire signal_13982 ;
    wire signal_13983 ;
    wire signal_13984 ;
    wire signal_13985 ;
    wire signal_13986 ;
    wire signal_13987 ;
    wire signal_13988 ;
    wire signal_13989 ;
    wire signal_13990 ;
    wire signal_13991 ;
    wire signal_13992 ;
    wire signal_13993 ;
    wire signal_13994 ;
    wire signal_13995 ;
    wire signal_13996 ;
    wire signal_13997 ;
    wire signal_13998 ;
    wire signal_13999 ;
    wire signal_14000 ;
    wire signal_14001 ;
    wire signal_14002 ;
    wire signal_14003 ;
    wire signal_14004 ;
    wire signal_14005 ;
    wire signal_14006 ;
    wire signal_14007 ;
    wire signal_14008 ;
    wire signal_14009 ;
    wire signal_14010 ;
    wire signal_14011 ;
    wire signal_14012 ;
    wire signal_14013 ;
    wire signal_14014 ;
    wire signal_14015 ;
    wire signal_14016 ;
    wire signal_14017 ;
    wire signal_14018 ;
    wire signal_14019 ;
    wire signal_14020 ;
    wire signal_14021 ;
    wire signal_14022 ;
    wire signal_14023 ;
    wire signal_14024 ;
    wire signal_14025 ;
    wire signal_14026 ;
    wire signal_14027 ;
    wire signal_14028 ;
    wire signal_14029 ;
    wire signal_14030 ;
    wire signal_14031 ;
    wire signal_14032 ;
    wire signal_14033 ;
    wire signal_14034 ;
    wire signal_14035 ;
    wire signal_14036 ;
    wire signal_14037 ;
    wire signal_14038 ;
    wire signal_14039 ;
    wire signal_14040 ;
    wire signal_14041 ;
    wire signal_14042 ;
    wire signal_14043 ;
    wire signal_14044 ;
    wire signal_14045 ;
    wire signal_14046 ;
    wire signal_14047 ;
    wire signal_14048 ;
    wire signal_14049 ;
    wire signal_14050 ;
    wire signal_14051 ;
    wire signal_14052 ;
    wire signal_14053 ;
    wire signal_14054 ;
    wire signal_14055 ;
    wire signal_14056 ;
    wire signal_14057 ;
    wire signal_14058 ;
    wire signal_14059 ;
    wire signal_14060 ;
    wire signal_14061 ;
    wire signal_14062 ;
    wire signal_14063 ;
    wire signal_14064 ;
    wire signal_14065 ;
    wire signal_14066 ;
    wire signal_14067 ;
    wire signal_14068 ;
    wire signal_14069 ;
    wire signal_14070 ;
    wire signal_14071 ;
    wire signal_14072 ;
    wire signal_14073 ;
    wire signal_14074 ;
    wire signal_14075 ;
    wire signal_14076 ;
    wire signal_14077 ;
    wire signal_14078 ;
    wire signal_14079 ;
    wire signal_14080 ;
    wire signal_14081 ;
    wire signal_14082 ;
    wire signal_14083 ;
    wire signal_14084 ;
    wire signal_14085 ;
    wire signal_14086 ;
    wire signal_14087 ;
    wire signal_14088 ;
    wire signal_14089 ;
    wire signal_14090 ;
    wire signal_14091 ;
    wire signal_14092 ;
    wire signal_14093 ;
    wire signal_14094 ;
    wire signal_14095 ;
    wire signal_14096 ;
    wire signal_14097 ;
    wire signal_14098 ;
    wire signal_14099 ;
    wire signal_14100 ;
    wire signal_14101 ;
    wire signal_14102 ;
    wire signal_14103 ;
    wire signal_14104 ;
    wire signal_14105 ;
    wire signal_14106 ;
    wire signal_14107 ;
    wire signal_14108 ;
    wire signal_14109 ;
    wire signal_14110 ;
    wire signal_14111 ;
    wire signal_14112 ;
    wire signal_14113 ;
    wire signal_14114 ;
    wire signal_14115 ;
    wire signal_14116 ;
    wire signal_14117 ;
    wire signal_14118 ;
    wire signal_14119 ;
    wire signal_14120 ;
    wire signal_14121 ;
    wire signal_14122 ;
    wire signal_14123 ;
    wire signal_14124 ;
    wire signal_14125 ;
    wire signal_14126 ;
    wire signal_14127 ;
    wire signal_14128 ;
    wire signal_14129 ;
    wire signal_14130 ;
    wire signal_14131 ;
    wire signal_14132 ;
    wire signal_14133 ;
    wire signal_14134 ;
    wire signal_14135 ;
    wire signal_14136 ;
    wire signal_14137 ;
    wire signal_14138 ;
    wire signal_14139 ;
    wire signal_14140 ;
    wire signal_14141 ;
    wire signal_14142 ;
    wire signal_14143 ;
    wire signal_14144 ;
    wire signal_14145 ;
    wire signal_14146 ;
    wire signal_14147 ;
    wire signal_14148 ;
    wire signal_14149 ;
    wire signal_14150 ;
    wire signal_14151 ;
    wire signal_14152 ;
    wire signal_14153 ;
    wire signal_14154 ;
    wire signal_14155 ;
    wire signal_14156 ;
    wire signal_14157 ;
    wire signal_14158 ;
    wire signal_14159 ;
    wire signal_14160 ;
    wire signal_14161 ;
    wire signal_14162 ;
    wire signal_14163 ;
    wire signal_14164 ;
    wire signal_14165 ;
    wire signal_14166 ;
    wire signal_14167 ;
    wire signal_14168 ;
    wire signal_14169 ;
    wire signal_14170 ;
    wire signal_14171 ;
    wire signal_14172 ;
    wire signal_14173 ;
    wire signal_14174 ;
    wire signal_14175 ;
    wire signal_14176 ;
    wire signal_14177 ;
    wire signal_14178 ;
    wire signal_14179 ;
    wire signal_14180 ;
    wire signal_14181 ;
    wire signal_14182 ;
    wire signal_14183 ;
    wire signal_14184 ;
    wire signal_14185 ;
    wire signal_14186 ;
    wire signal_14187 ;
    wire signal_14188 ;
    wire signal_14189 ;
    wire signal_14190 ;
    wire signal_14191 ;
    wire signal_14192 ;
    wire signal_14193 ;
    wire signal_14194 ;
    wire signal_14195 ;
    wire signal_14196 ;
    wire signal_14197 ;
    wire signal_14198 ;
    wire signal_14199 ;
    wire signal_14200 ;
    wire signal_14201 ;
    wire signal_14202 ;
    wire signal_14203 ;
    wire signal_14204 ;
    wire signal_14205 ;
    wire signal_14206 ;
    wire signal_14207 ;
    wire signal_14208 ;
    wire signal_14209 ;
    wire signal_14210 ;
    wire signal_14211 ;
    wire signal_14212 ;
    wire signal_14213 ;
    wire signal_14214 ;
    wire signal_14215 ;
    wire signal_14216 ;
    wire signal_14217 ;
    wire signal_14218 ;
    wire signal_14219 ;
    wire signal_14220 ;
    wire signal_14221 ;
    wire signal_14222 ;
    wire signal_14223 ;
    wire signal_14224 ;
    wire signal_14225 ;
    wire signal_14226 ;
    wire signal_14227 ;
    wire signal_14228 ;
    wire signal_14229 ;
    wire signal_14230 ;
    wire signal_14231 ;
    wire signal_14232 ;
    wire signal_14233 ;
    wire signal_14234 ;
    wire signal_14235 ;
    wire signal_14236 ;
    wire signal_14237 ;
    wire signal_14238 ;
    wire signal_14239 ;
    wire signal_14240 ;
    wire signal_14241 ;
    wire signal_14242 ;
    wire signal_14243 ;
    wire signal_14244 ;
    wire signal_14245 ;
    wire signal_14246 ;
    wire signal_14247 ;
    wire signal_14248 ;
    wire signal_14249 ;
    wire signal_14250 ;
    wire signal_14251 ;
    wire signal_14252 ;
    wire signal_14253 ;
    wire signal_14254 ;
    wire signal_14255 ;
    wire signal_14256 ;
    wire signal_14257 ;
    wire signal_14258 ;
    wire signal_14259 ;
    wire signal_14260 ;
    wire signal_14261 ;
    wire signal_14262 ;
    wire signal_14263 ;
    wire signal_14264 ;
    wire signal_14265 ;
    wire signal_14266 ;
    wire signal_14267 ;
    wire signal_14268 ;
    wire signal_14269 ;
    wire signal_14270 ;
    wire signal_14271 ;
    wire signal_14272 ;
    wire signal_14273 ;
    wire signal_14274 ;
    wire signal_14275 ;
    wire signal_14276 ;
    wire signal_14277 ;
    wire signal_14278 ;
    wire signal_14279 ;
    wire signal_14280 ;
    wire signal_14281 ;
    wire signal_14282 ;
    wire signal_14283 ;
    wire signal_14284 ;
    wire signal_14285 ;
    wire signal_14286 ;
    wire signal_14287 ;
    wire signal_14288 ;
    wire signal_14289 ;
    wire signal_14290 ;
    wire signal_14291 ;
    wire signal_14292 ;
    wire signal_14293 ;
    wire signal_14294 ;
    wire signal_14295 ;
    wire signal_14296 ;
    wire signal_14297 ;
    wire signal_14298 ;
    wire signal_14299 ;
    wire signal_14300 ;
    wire signal_14301 ;
    wire signal_14302 ;
    wire signal_14303 ;
    wire signal_14304 ;
    wire signal_14305 ;
    wire signal_14306 ;
    wire signal_14307 ;
    wire signal_14308 ;
    wire signal_14309 ;
    wire signal_14310 ;
    wire signal_14311 ;
    wire signal_14312 ;
    wire signal_14313 ;
    wire signal_14314 ;
    wire signal_14315 ;
    wire signal_14316 ;
    wire signal_14317 ;
    wire signal_14318 ;
    wire signal_14319 ;
    wire signal_14320 ;
    wire signal_14321 ;
    wire signal_14322 ;
    wire signal_14323 ;
    wire signal_14324 ;
    wire signal_14325 ;
    wire signal_14326 ;
    wire signal_14327 ;
    wire signal_14328 ;
    wire signal_14329 ;
    wire signal_14330 ;
    wire signal_14331 ;
    wire signal_14332 ;
    wire signal_14333 ;
    wire signal_14334 ;
    wire signal_14335 ;
    wire signal_14336 ;
    wire signal_14337 ;
    wire signal_14338 ;
    wire signal_14339 ;
    wire signal_14340 ;
    wire signal_14341 ;
    wire signal_14342 ;
    wire signal_14343 ;
    wire signal_14344 ;
    wire signal_14345 ;
    wire signal_14346 ;
    wire signal_14347 ;
    wire signal_14348 ;
    wire signal_14349 ;
    wire signal_14350 ;
    wire signal_14351 ;
    wire signal_14352 ;
    wire signal_14353 ;
    wire signal_14354 ;
    wire signal_14355 ;
    wire signal_14356 ;
    wire signal_14357 ;
    wire signal_14358 ;
    wire signal_14359 ;
    wire signal_14360 ;
    wire signal_14361 ;
    wire signal_14362 ;
    wire signal_14363 ;
    wire signal_14364 ;
    wire signal_14365 ;
    wire signal_14366 ;
    wire signal_14367 ;
    wire signal_14368 ;
    wire signal_14369 ;
    wire signal_14370 ;
    wire signal_14371 ;
    wire signal_14372 ;
    wire signal_14373 ;
    wire signal_14374 ;
    wire signal_14375 ;
    wire signal_14376 ;
    wire signal_14377 ;
    wire signal_14378 ;
    wire signal_14379 ;
    wire signal_14380 ;
    wire signal_14381 ;
    wire signal_14382 ;
    wire signal_14383 ;
    wire signal_14384 ;
    wire signal_14385 ;
    wire signal_14386 ;
    wire signal_14387 ;
    wire signal_14388 ;
    wire signal_14389 ;
    wire signal_14390 ;
    wire signal_14391 ;
    wire signal_14392 ;
    wire signal_14393 ;
    wire signal_14394 ;
    wire signal_14395 ;
    wire signal_14396 ;
    wire signal_14397 ;
    wire signal_14398 ;
    wire signal_14399 ;
    wire signal_14400 ;
    wire signal_14401 ;
    wire signal_14402 ;
    wire signal_14403 ;
    wire signal_14404 ;
    wire signal_14405 ;
    wire signal_14406 ;
    wire signal_14407 ;
    wire signal_14408 ;
    wire signal_14409 ;
    wire signal_14410 ;
    wire signal_14411 ;
    wire signal_14412 ;
    wire signal_14413 ;
    wire signal_14414 ;
    wire signal_14415 ;
    wire signal_14416 ;
    wire signal_14417 ;
    wire signal_14418 ;
    wire signal_14419 ;
    wire signal_14420 ;
    wire signal_14421 ;
    wire signal_14422 ;
    wire signal_14423 ;
    wire signal_14424 ;
    wire signal_14425 ;
    wire signal_14426 ;
    wire signal_14427 ;
    wire signal_14428 ;
    wire signal_14429 ;
    wire signal_14430 ;
    wire signal_14431 ;
    wire signal_14432 ;
    wire signal_14433 ;
    wire signal_14434 ;
    wire signal_14435 ;
    wire signal_14436 ;
    wire signal_14437 ;
    wire signal_14438 ;
    wire signal_14439 ;
    wire signal_14440 ;
    wire signal_14441 ;
    wire signal_14442 ;
    wire signal_14443 ;
    wire signal_14444 ;
    wire signal_14445 ;
    wire signal_14446 ;
    wire signal_14447 ;
    wire signal_14448 ;
    wire signal_14449 ;
    wire signal_14450 ;
    wire signal_14451 ;
    wire signal_14452 ;
    wire signal_14453 ;
    wire signal_14454 ;
    wire signal_14455 ;
    wire signal_14456 ;
    wire signal_14457 ;
    wire signal_14458 ;
    wire signal_14459 ;
    wire signal_14460 ;
    wire signal_14461 ;
    wire signal_14462 ;
    wire signal_14463 ;
    wire signal_14464 ;
    wire signal_14465 ;
    wire signal_14466 ;
    wire signal_14467 ;
    wire signal_14468 ;
    wire signal_14469 ;
    wire signal_14470 ;
    wire signal_14471 ;
    wire signal_14472 ;
    wire signal_14473 ;
    wire signal_14474 ;
    wire signal_14475 ;
    wire signal_14476 ;
    wire signal_14477 ;
    wire signal_14478 ;
    wire signal_14479 ;
    wire signal_14480 ;
    wire signal_14481 ;
    wire signal_14482 ;
    wire signal_14483 ;
    wire signal_14484 ;
    wire signal_14485 ;
    wire signal_14486 ;
    wire signal_14487 ;
    wire signal_14488 ;
    wire signal_14489 ;
    wire signal_14490 ;
    wire signal_14491 ;
    wire signal_14492 ;
    wire signal_14493 ;
    wire signal_14494 ;
    wire signal_14495 ;
    wire signal_14496 ;
    wire signal_14497 ;
    wire signal_14498 ;
    wire signal_14499 ;
    wire signal_14500 ;
    wire signal_14501 ;
    wire signal_14502 ;
    wire signal_14503 ;
    wire signal_14504 ;
    wire signal_14505 ;
    wire signal_14506 ;
    wire signal_14507 ;
    wire signal_14508 ;
    wire signal_14509 ;
    wire signal_14510 ;
    wire signal_14511 ;
    wire signal_14512 ;
    wire signal_14513 ;
    wire signal_14514 ;
    wire signal_14515 ;
    wire signal_14516 ;
    wire signal_14517 ;
    wire signal_14518 ;
    wire signal_14519 ;
    wire signal_14520 ;
    wire signal_14521 ;
    wire signal_14522 ;
    wire signal_14523 ;
    wire signal_14524 ;
    wire signal_14525 ;
    wire signal_14526 ;
    wire signal_14527 ;
    wire signal_14528 ;
    wire signal_14529 ;
    wire signal_14530 ;
    wire signal_14531 ;
    wire signal_14532 ;
    wire signal_14533 ;
    wire signal_14534 ;
    wire signal_14535 ;
    wire signal_14536 ;
    wire signal_14537 ;
    wire signal_14538 ;
    wire signal_14539 ;
    wire signal_14540 ;
    wire signal_14541 ;
    wire signal_14542 ;
    wire signal_14543 ;
    wire signal_14544 ;
    wire signal_14545 ;
    wire signal_14546 ;
    wire signal_14547 ;
    wire signal_14548 ;
    wire signal_14549 ;
    wire signal_14550 ;
    wire signal_14551 ;
    wire signal_14552 ;
    wire signal_14553 ;
    wire signal_14554 ;
    wire signal_14555 ;
    wire signal_14556 ;
    wire signal_14557 ;
    wire signal_14558 ;
    wire signal_14559 ;
    wire signal_14560 ;
    wire signal_14561 ;
    wire signal_14562 ;
    wire signal_14563 ;
    wire signal_14564 ;
    wire signal_14565 ;
    wire signal_14566 ;
    wire signal_14567 ;
    wire signal_14568 ;
    wire signal_14569 ;
    wire signal_14570 ;
    wire signal_14571 ;
    wire signal_14572 ;
    wire signal_14573 ;
    wire signal_14574 ;
    wire signal_14575 ;
    wire signal_14576 ;
    wire signal_14577 ;
    wire signal_14578 ;
    wire signal_14579 ;
    wire signal_14580 ;
    wire signal_14581 ;
    wire signal_14582 ;
    wire signal_14583 ;
    wire signal_14584 ;
    wire signal_14585 ;
    wire signal_14586 ;
    wire signal_14587 ;
    wire signal_14588 ;
    wire signal_14589 ;
    wire signal_14590 ;
    wire signal_14591 ;
    wire signal_14592 ;
    wire signal_14593 ;
    wire signal_14594 ;
    wire signal_14595 ;
    wire signal_14596 ;
    wire signal_14597 ;
    wire signal_14598 ;
    wire signal_14599 ;
    wire signal_14600 ;
    wire signal_14601 ;
    wire signal_14602 ;
    wire signal_14603 ;
    wire signal_14604 ;
    wire signal_14605 ;
    wire signal_14606 ;
    wire signal_14607 ;
    wire signal_14608 ;
    wire signal_14609 ;
    wire signal_14610 ;
    wire signal_14611 ;
    wire signal_14612 ;
    wire signal_14613 ;
    wire signal_14614 ;
    wire signal_14615 ;
    wire signal_14616 ;
    wire signal_14617 ;
    wire signal_14618 ;
    wire signal_14619 ;
    wire signal_14620 ;
    wire signal_14621 ;
    wire signal_14622 ;
    wire signal_14623 ;
    wire signal_14624 ;
    wire signal_14625 ;
    wire signal_14626 ;
    wire signal_14627 ;
    wire signal_14628 ;
    wire signal_14629 ;
    wire signal_14630 ;
    wire signal_14631 ;
    wire signal_14632 ;
    wire signal_14633 ;
    wire signal_14634 ;
    wire signal_14635 ;
    wire signal_14636 ;
    wire signal_14637 ;
    wire signal_14638 ;
    wire signal_14639 ;
    wire signal_14640 ;
    wire signal_14641 ;
    wire signal_14642 ;
    wire signal_14643 ;
    wire signal_14644 ;
    wire signal_14645 ;
    wire signal_14646 ;
    wire signal_14647 ;
    wire signal_14648 ;
    wire signal_14649 ;
    wire signal_14650 ;
    wire signal_14651 ;
    wire signal_14652 ;
    wire signal_14653 ;
    wire signal_14654 ;
    wire signal_14655 ;
    wire signal_14656 ;
    wire signal_14657 ;
    wire signal_14658 ;
    wire signal_14659 ;
    wire signal_14660 ;
    wire signal_14661 ;
    wire signal_14662 ;
    wire signal_14663 ;
    wire signal_14664 ;
    wire signal_14665 ;
    wire signal_14666 ;
    wire signal_14667 ;
    wire signal_14668 ;
    wire signal_14669 ;
    wire signal_14670 ;
    wire signal_14671 ;
    wire signal_14672 ;
    wire signal_14673 ;
    wire signal_14674 ;
    wire signal_14675 ;
    wire signal_14676 ;
    wire signal_14677 ;
    wire signal_14678 ;
    wire signal_14679 ;
    wire signal_14680 ;
    wire signal_14681 ;
    wire signal_14682 ;
    wire signal_14683 ;
    wire signal_14684 ;
    wire signal_14685 ;
    wire signal_14686 ;
    wire signal_14687 ;
    wire signal_14688 ;
    wire signal_14689 ;
    wire signal_14690 ;
    wire signal_14691 ;
    wire signal_14692 ;
    wire signal_14693 ;
    wire signal_14694 ;
    wire signal_14695 ;
    wire signal_14696 ;
    wire signal_14697 ;
    wire signal_14698 ;
    wire signal_14699 ;
    wire signal_14700 ;
    wire signal_14701 ;
    wire signal_14702 ;
    wire signal_14703 ;
    wire signal_14704 ;
    wire signal_14705 ;
    wire signal_14706 ;
    wire signal_14707 ;
    wire signal_14708 ;
    wire signal_14709 ;
    wire signal_14710 ;
    wire signal_14711 ;
    wire signal_14712 ;
    wire signal_14713 ;
    wire signal_14714 ;
    wire signal_14715 ;
    wire signal_14716 ;
    wire signal_14717 ;
    wire signal_14718 ;
    wire signal_14719 ;
    wire signal_14720 ;
    wire signal_14721 ;
    wire signal_14722 ;
    wire signal_14723 ;
    wire signal_14724 ;
    wire signal_14725 ;
    wire signal_14726 ;
    wire signal_14727 ;
    wire signal_14728 ;
    wire signal_14729 ;
    wire signal_14730 ;
    wire signal_14731 ;
    wire signal_14732 ;
    wire signal_14733 ;
    wire signal_14734 ;
    wire signal_14735 ;
    wire signal_14736 ;
    wire signal_14737 ;
    wire signal_14738 ;
    wire signal_14739 ;
    wire signal_14740 ;
    wire signal_14741 ;
    wire signal_14742 ;
    wire signal_14743 ;
    wire signal_14744 ;
    wire signal_14745 ;
    wire signal_14746 ;
    wire signal_14747 ;
    wire signal_14748 ;
    wire signal_14749 ;
    wire signal_14750 ;
    wire signal_14751 ;
    wire signal_14752 ;
    wire signal_14753 ;
    wire signal_14754 ;
    wire signal_14755 ;
    wire signal_14756 ;
    wire signal_14757 ;
    wire signal_14758 ;
    wire signal_14759 ;
    wire signal_14760 ;
    wire signal_14761 ;
    wire signal_14762 ;
    wire signal_14763 ;
    wire signal_14764 ;
    wire signal_14765 ;
    wire signal_14766 ;
    wire signal_14767 ;
    wire signal_14768 ;
    wire signal_14769 ;
    wire signal_14770 ;
    wire signal_14771 ;
    wire signal_14772 ;
    wire signal_14773 ;
    wire signal_14774 ;
    wire signal_14775 ;
    wire signal_14776 ;
    wire signal_14777 ;
    wire signal_14778 ;
    wire signal_14779 ;
    wire signal_14780 ;
    wire signal_14781 ;
    wire signal_14782 ;
    wire signal_14783 ;
    wire signal_14784 ;
    wire signal_14785 ;
    wire signal_14786 ;
    wire signal_14787 ;
    wire signal_14788 ;
    wire signal_14789 ;
    wire signal_14790 ;
    wire signal_14791 ;
    wire signal_14792 ;
    wire signal_14793 ;
    wire signal_14794 ;
    wire signal_14795 ;
    wire signal_14796 ;
    wire signal_14797 ;
    wire signal_14798 ;
    wire signal_14799 ;
    wire signal_14800 ;
    wire signal_14801 ;
    wire signal_14802 ;
    wire signal_14803 ;
    wire signal_14804 ;
    wire signal_14805 ;
    wire signal_14806 ;
    wire signal_14807 ;
    wire signal_14808 ;
    wire signal_14809 ;
    wire signal_14810 ;
    wire signal_14811 ;
    wire signal_14812 ;
    wire signal_14813 ;
    wire signal_14814 ;
    wire signal_14815 ;
    wire signal_14816 ;
    wire signal_14817 ;
    wire signal_14818 ;
    wire signal_14819 ;
    wire signal_14820 ;
    wire signal_14821 ;
    wire signal_14822 ;
    wire signal_14823 ;
    wire signal_14824 ;
    wire signal_14825 ;
    wire signal_14826 ;
    wire signal_14827 ;
    wire signal_14828 ;
    wire signal_14829 ;
    wire signal_14830 ;
    wire signal_14831 ;
    wire signal_14832 ;
    wire signal_14833 ;
    wire signal_14834 ;
    wire signal_14835 ;
    wire signal_14836 ;
    wire signal_14837 ;
    wire signal_14838 ;
    wire signal_14839 ;
    wire signal_14840 ;
    wire signal_14841 ;
    wire signal_14842 ;
    wire signal_14843 ;
    wire signal_14844 ;
    wire signal_14845 ;
    wire signal_14846 ;
    wire signal_14847 ;
    wire signal_14848 ;
    wire signal_14849 ;
    wire signal_14850 ;
    wire signal_14851 ;
    wire signal_14852 ;
    wire signal_14853 ;
    wire signal_14854 ;
    wire signal_14855 ;
    wire signal_14856 ;
    wire signal_14857 ;
    wire signal_14858 ;
    wire signal_14859 ;
    wire signal_14860 ;
    wire signal_14861 ;
    wire signal_14862 ;
    wire signal_14863 ;
    wire signal_14864 ;
    wire signal_14865 ;
    wire signal_14866 ;
    wire signal_14867 ;
    wire signal_14868 ;
    wire signal_14869 ;
    wire signal_14870 ;
    wire signal_14871 ;
    wire signal_14872 ;
    wire signal_14873 ;
    wire signal_14874 ;
    wire signal_14875 ;
    wire signal_14876 ;
    wire signal_14877 ;
    wire signal_14878 ;
    wire signal_14879 ;
    wire signal_14880 ;
    wire signal_14881 ;
    wire signal_14882 ;
    wire signal_14883 ;
    wire signal_14884 ;
    wire signal_14885 ;
    wire signal_14886 ;
    wire signal_14887 ;
    wire signal_14888 ;
    wire signal_14889 ;
    wire signal_14890 ;
    wire signal_14891 ;
    wire signal_14892 ;
    wire signal_14893 ;
    wire signal_14894 ;
    wire signal_14895 ;
    wire signal_14896 ;
    wire signal_14897 ;
    wire signal_14898 ;
    wire signal_14899 ;
    wire signal_14900 ;
    wire signal_14901 ;
    wire signal_14902 ;
    wire signal_14903 ;
    wire signal_14904 ;
    wire signal_14905 ;
    wire signal_14906 ;
    wire signal_14907 ;
    wire signal_14908 ;
    wire signal_14909 ;
    wire signal_14910 ;
    wire signal_14911 ;
    wire signal_14912 ;
    wire signal_14913 ;
    wire signal_14914 ;
    wire signal_14915 ;
    wire signal_14916 ;
    wire signal_14917 ;
    wire signal_14918 ;
    wire signal_14919 ;
    wire signal_14920 ;
    wire signal_14921 ;
    wire signal_14922 ;
    wire signal_14923 ;
    wire signal_14924 ;
    wire signal_14925 ;
    wire signal_14926 ;
    wire signal_14927 ;
    wire signal_14928 ;
    wire signal_14929 ;
    wire signal_14930 ;
    wire signal_14931 ;
    wire signal_14932 ;
    wire signal_14933 ;
    wire signal_14934 ;
    wire signal_14935 ;
    wire signal_14936 ;
    wire signal_14937 ;
    wire signal_14938 ;
    wire signal_14939 ;
    wire signal_14940 ;
    wire signal_14941 ;
    wire signal_14942 ;
    wire signal_14943 ;
    wire signal_14944 ;
    wire signal_14945 ;
    wire signal_14946 ;
    wire signal_14947 ;
    wire signal_14948 ;
    wire signal_14949 ;
    wire signal_14950 ;
    wire signal_14951 ;
    wire signal_14952 ;
    wire signal_14953 ;
    wire signal_14954 ;
    wire signal_14955 ;
    wire signal_14956 ;
    wire signal_14957 ;
    wire signal_14958 ;
    wire signal_14959 ;
    wire signal_14960 ;
    wire signal_14961 ;
    wire signal_14962 ;
    wire signal_14963 ;
    wire signal_14964 ;
    wire signal_14965 ;
    wire signal_14966 ;
    wire signal_14967 ;
    wire signal_14968 ;
    wire signal_14969 ;
    wire signal_14970 ;
    wire signal_14971 ;
    wire signal_14972 ;
    wire signal_14973 ;
    wire signal_14974 ;
    wire signal_14975 ;
    wire signal_14976 ;
    wire signal_14977 ;
    wire signal_14978 ;
    wire signal_14979 ;
    wire signal_14980 ;
    wire signal_14981 ;
    wire signal_14982 ;
    wire signal_14983 ;
    wire signal_14984 ;
    wire signal_14985 ;
    wire signal_14986 ;
    wire signal_14987 ;
    wire signal_14988 ;
    wire signal_14989 ;
    wire signal_14990 ;
    wire signal_14991 ;
    wire signal_14992 ;
    wire signal_14993 ;
    wire signal_14994 ;
    wire signal_14995 ;
    wire signal_14996 ;
    wire signal_14997 ;
    wire signal_14998 ;
    wire signal_14999 ;
    wire signal_15000 ;
    wire signal_15001 ;
    wire signal_15002 ;
    wire signal_15003 ;
    wire signal_15004 ;
    wire signal_15005 ;
    wire signal_15006 ;
    wire signal_15007 ;
    wire signal_15008 ;
    wire signal_15009 ;
    wire signal_15010 ;
    wire signal_15011 ;
    wire signal_15012 ;
    wire signal_15013 ;
    wire signal_15014 ;
    wire signal_15015 ;
    wire signal_15016 ;
    wire signal_15017 ;
    wire signal_15018 ;
    wire signal_15019 ;
    wire signal_15020 ;
    wire signal_15021 ;
    wire signal_15022 ;
    wire signal_15023 ;
    wire signal_15024 ;
    wire signal_15025 ;
    wire signal_15026 ;
    wire signal_15027 ;
    wire signal_15028 ;
    wire signal_15029 ;
    wire signal_15030 ;
    wire signal_15031 ;
    wire signal_15032 ;
    wire signal_15033 ;
    wire signal_15034 ;
    wire signal_15035 ;
    wire signal_15036 ;
    wire signal_15037 ;
    wire signal_15038 ;
    wire signal_15039 ;
    wire signal_15040 ;
    wire signal_15041 ;
    wire signal_15042 ;
    wire signal_15043 ;
    wire signal_15044 ;
    wire signal_15045 ;
    wire signal_15046 ;
    wire signal_15047 ;
    wire signal_15048 ;
    wire signal_15049 ;
    wire signal_15050 ;
    wire signal_15051 ;
    wire signal_15052 ;
    wire signal_15053 ;
    wire signal_15054 ;
    wire signal_15055 ;
    wire signal_15056 ;
    wire signal_15057 ;
    wire signal_15058 ;
    wire signal_15059 ;
    wire signal_15060 ;
    wire signal_15061 ;
    wire signal_15062 ;
    wire signal_15063 ;
    wire signal_15064 ;
    wire signal_15065 ;
    wire signal_15066 ;
    wire signal_15067 ;
    wire signal_15068 ;
    wire signal_15069 ;
    wire signal_15070 ;
    wire signal_15071 ;
    wire signal_15072 ;
    wire signal_15073 ;
    wire signal_15074 ;
    wire signal_15075 ;
    wire signal_15076 ;
    wire signal_15077 ;
    wire signal_15078 ;
    wire signal_15079 ;
    wire signal_15080 ;
    wire signal_15081 ;
    wire signal_15082 ;
    wire signal_15083 ;
    wire signal_15084 ;
    wire signal_15085 ;
    wire signal_15086 ;
    wire signal_15087 ;
    wire signal_15088 ;
    wire signal_15089 ;
    wire signal_15090 ;
    wire signal_15091 ;
    wire signal_15092 ;
    wire signal_15093 ;
    wire signal_15094 ;
    wire signal_15095 ;
    wire signal_15096 ;
    wire signal_15097 ;
    wire signal_15098 ;
    wire signal_15099 ;
    wire signal_15100 ;
    wire signal_15101 ;
    wire signal_15102 ;
    wire signal_15103 ;
    wire signal_15104 ;
    wire signal_15105 ;
    wire signal_15106 ;
    wire signal_15107 ;
    wire signal_15108 ;
    wire signal_15109 ;
    wire signal_15110 ;
    wire signal_15111 ;
    wire signal_15112 ;
    wire signal_15113 ;
    wire signal_15114 ;
    wire signal_15115 ;
    wire signal_15116 ;
    wire signal_15117 ;
    wire signal_15118 ;
    wire signal_15119 ;
    wire signal_15120 ;
    wire signal_15121 ;
    wire signal_15122 ;
    wire signal_15123 ;
    wire signal_15124 ;
    wire signal_15125 ;
    wire signal_15126 ;
    wire signal_15127 ;
    wire signal_15128 ;
    wire signal_15129 ;
    wire signal_15130 ;
    wire signal_15131 ;
    wire signal_15132 ;
    wire signal_15133 ;
    wire signal_15134 ;
    wire signal_15135 ;
    wire signal_15136 ;
    wire signal_15137 ;
    wire signal_15138 ;
    wire signal_15139 ;
    wire signal_15140 ;
    wire signal_15141 ;
    wire signal_15142 ;
    wire signal_15143 ;
    wire signal_15144 ;
    wire signal_15145 ;
    wire signal_15146 ;
    wire signal_15147 ;
    wire signal_15148 ;
    wire signal_15149 ;
    wire signal_15150 ;
    wire signal_15151 ;
    wire signal_15152 ;
    wire signal_15153 ;
    wire signal_15154 ;
    wire signal_15155 ;
    wire signal_15156 ;
    wire signal_15157 ;
    wire signal_15158 ;
    wire signal_15159 ;
    wire signal_15160 ;
    wire signal_15161 ;
    wire signal_15162 ;
    wire signal_15163 ;
    wire signal_15164 ;
    wire signal_15165 ;
    wire signal_15166 ;
    wire signal_15167 ;
    wire signal_15168 ;
    wire signal_15169 ;
    wire signal_15170 ;
    wire signal_15171 ;
    wire signal_15172 ;
    wire signal_15173 ;
    wire signal_15174 ;
    wire signal_15175 ;
    wire signal_15176 ;
    wire signal_15177 ;
    wire signal_15178 ;
    wire signal_15179 ;
    wire signal_15180 ;
    wire signal_15181 ;
    wire signal_15182 ;
    wire signal_15183 ;
    wire signal_15184 ;
    wire signal_15185 ;
    wire signal_15186 ;
    wire signal_15187 ;
    wire signal_15188 ;
    wire signal_15189 ;
    wire signal_15190 ;
    wire signal_15191 ;
    wire signal_15192 ;
    wire signal_15193 ;
    wire signal_15194 ;
    wire signal_15195 ;
    wire signal_15196 ;
    wire signal_15197 ;
    wire signal_15198 ;
    wire signal_15199 ;
    wire signal_15200 ;
    wire signal_15201 ;
    wire signal_15202 ;
    wire signal_15203 ;
    wire signal_15204 ;
    wire signal_15205 ;
    wire signal_15206 ;
    wire signal_15207 ;
    wire signal_15208 ;
    wire signal_15209 ;
    wire signal_15210 ;
    wire signal_15211 ;
    wire signal_15212 ;
    wire signal_15213 ;
    wire signal_15214 ;
    wire signal_15215 ;
    wire signal_15216 ;
    wire signal_15217 ;
    wire signal_15218 ;
    wire signal_15219 ;
    wire signal_15220 ;
    wire signal_15221 ;
    wire signal_15222 ;
    wire signal_15223 ;
    wire signal_15224 ;
    wire signal_15225 ;
    wire signal_15226 ;
    wire signal_15227 ;
    wire signal_15228 ;
    wire signal_15229 ;
    wire signal_15230 ;
    wire signal_15231 ;
    wire signal_15232 ;
    wire signal_15233 ;
    wire signal_15234 ;
    wire signal_15235 ;
    wire signal_15236 ;
    wire signal_15237 ;
    wire signal_15238 ;
    wire signal_15239 ;
    wire signal_15240 ;
    wire signal_15241 ;
    wire signal_15242 ;
    wire signal_15243 ;
    wire signal_15244 ;
    wire signal_15245 ;
    wire signal_15246 ;
    wire signal_15247 ;
    wire signal_15248 ;
    wire signal_15249 ;
    wire signal_15250 ;
    wire signal_15251 ;
    wire signal_15252 ;
    wire signal_15253 ;
    wire signal_15254 ;
    wire signal_15255 ;
    wire signal_15256 ;
    wire signal_15257 ;
    wire signal_15258 ;
    wire signal_15259 ;
    wire signal_15260 ;
    wire signal_15261 ;
    wire signal_15262 ;
    wire signal_15263 ;
    wire signal_15264 ;
    wire signal_15265 ;
    wire signal_15266 ;
    wire signal_15267 ;
    wire signal_15268 ;
    wire signal_15269 ;
    wire signal_15270 ;
    wire signal_15271 ;
    wire signal_15272 ;
    wire signal_15273 ;
    wire signal_15274 ;
    wire signal_15275 ;
    wire signal_15276 ;
    wire signal_15277 ;
    wire signal_15278 ;
    wire signal_15279 ;
    wire signal_15280 ;
    wire signal_15281 ;
    wire signal_15282 ;
    wire signal_15283 ;
    wire signal_15284 ;
    wire signal_15285 ;
    wire signal_15286 ;
    wire signal_15287 ;
    wire signal_15288 ;
    wire signal_15289 ;
    wire signal_15290 ;
    wire signal_15291 ;
    wire signal_15292 ;
    wire signal_15293 ;
    wire signal_15294 ;
    wire signal_15295 ;
    wire signal_15296 ;
    wire signal_15297 ;
    wire signal_15298 ;
    wire signal_15299 ;
    wire signal_15300 ;
    wire signal_15301 ;
    wire signal_15302 ;
    wire signal_15303 ;
    wire signal_15304 ;
    wire signal_15305 ;
    wire signal_15306 ;
    wire signal_15307 ;
    wire signal_15308 ;
    wire signal_15309 ;
    wire signal_15310 ;
    wire signal_15311 ;
    wire signal_15312 ;
    wire signal_15313 ;
    wire signal_15314 ;
    wire signal_15315 ;
    wire signal_15316 ;
    wire signal_15317 ;
    wire signal_15318 ;
    wire signal_15319 ;
    wire signal_15320 ;
    wire signal_15321 ;
    wire signal_15322 ;
    wire signal_15323 ;
    wire signal_15324 ;
    wire signal_15325 ;
    wire signal_15326 ;
    wire signal_15327 ;
    wire signal_15328 ;
    wire signal_15329 ;
    wire signal_15330 ;
    wire signal_15331 ;
    wire signal_15332 ;
    wire signal_15333 ;
    wire signal_15334 ;
    wire signal_15335 ;
    wire signal_15336 ;
    wire signal_15337 ;
    wire signal_15338 ;
    wire signal_15339 ;
    wire signal_15340 ;
    wire signal_15341 ;
    wire signal_15342 ;
    wire signal_15343 ;
    wire signal_15344 ;
    wire signal_15345 ;
    wire signal_15346 ;
    wire signal_15347 ;
    wire signal_15348 ;
    wire signal_15349 ;
    wire signal_15350 ;
    wire signal_15351 ;
    wire signal_15352 ;
    wire signal_15353 ;
    wire signal_15354 ;
    wire signal_15355 ;
    wire signal_15356 ;
    wire signal_15357 ;
    wire signal_15358 ;
    wire signal_15359 ;
    wire signal_15360 ;
    wire signal_15361 ;
    wire signal_15362 ;
    wire signal_15363 ;
    wire signal_15364 ;
    wire signal_15365 ;
    wire signal_15366 ;
    wire signal_15367 ;
    wire signal_15368 ;
    wire signal_15369 ;
    wire signal_15370 ;
    wire signal_15371 ;
    wire signal_15372 ;
    wire signal_15373 ;
    wire signal_15374 ;
    wire signal_15375 ;
    wire signal_15376 ;
    wire signal_15377 ;
    wire signal_15378 ;
    wire signal_15379 ;
    wire signal_15380 ;
    wire signal_15381 ;
    wire signal_15382 ;
    wire signal_15383 ;
    wire signal_15384 ;
    wire signal_15385 ;
    wire signal_15386 ;
    wire signal_15387 ;
    wire signal_15388 ;
    wire signal_15389 ;
    wire signal_15390 ;
    wire signal_15391 ;
    wire signal_15392 ;
    wire signal_15393 ;
    wire signal_15394 ;
    wire signal_15395 ;
    wire signal_15396 ;
    wire signal_15397 ;
    wire signal_15398 ;
    wire signal_15399 ;
    wire signal_15400 ;
    wire signal_15401 ;
    wire signal_15402 ;
    wire signal_15403 ;
    wire signal_15404 ;
    wire signal_15405 ;
    wire signal_15406 ;
    wire signal_15407 ;
    wire signal_15408 ;
    wire signal_15409 ;
    wire signal_15410 ;
    wire signal_15411 ;
    wire signal_15412 ;
    wire signal_15413 ;
    wire signal_15414 ;
    wire signal_15415 ;
    wire signal_15416 ;
    wire signal_15417 ;
    wire signal_15418 ;
    wire signal_15419 ;
    wire signal_15420 ;
    wire signal_15421 ;
    wire signal_15422 ;
    wire signal_15423 ;
    wire signal_15424 ;
    wire signal_15425 ;
    wire signal_15426 ;
    wire signal_15427 ;
    wire signal_15428 ;
    wire signal_15429 ;
    wire signal_15430 ;
    wire signal_15431 ;
    wire signal_15432 ;
    wire signal_15433 ;
    wire signal_15434 ;
    wire signal_15435 ;
    wire signal_15436 ;
    wire signal_15437 ;
    wire signal_15438 ;
    wire signal_15439 ;
    wire signal_15440 ;
    wire signal_15441 ;
    wire signal_15442 ;
    wire signal_15443 ;
    wire signal_15444 ;
    wire signal_15445 ;
    wire signal_15446 ;
    wire signal_15447 ;
    wire signal_15448 ;
    wire signal_15449 ;
    wire signal_15450 ;
    wire signal_15451 ;
    wire signal_15452 ;
    wire signal_15453 ;
    wire signal_15454 ;
    wire signal_15455 ;
    wire signal_15456 ;
    wire signal_15457 ;
    wire signal_15458 ;
    wire signal_15459 ;
    wire signal_15460 ;
    wire signal_15461 ;
    wire signal_15462 ;
    wire signal_15463 ;
    wire signal_15464 ;
    wire signal_15465 ;
    wire signal_15466 ;
    wire signal_15467 ;
    wire signal_15468 ;
    wire signal_15469 ;
    wire signal_15470 ;
    wire signal_15471 ;
    wire signal_15472 ;
    wire signal_15473 ;
    wire signal_15474 ;
    wire signal_15475 ;
    wire signal_15476 ;
    wire signal_15477 ;
    wire signal_15478 ;
    wire signal_15479 ;
    wire signal_15480 ;
    wire signal_15481 ;
    wire signal_15482 ;
    wire signal_15483 ;
    wire signal_15484 ;
    wire signal_15485 ;
    wire signal_15486 ;
    wire signal_15487 ;
    wire signal_15488 ;
    wire signal_15489 ;
    wire signal_15490 ;
    wire signal_15491 ;
    wire signal_15492 ;
    wire signal_15493 ;
    wire signal_15494 ;
    wire signal_15495 ;
    wire signal_15496 ;
    wire signal_15497 ;
    wire signal_15498 ;
    wire signal_15499 ;
    wire signal_15500 ;
    wire signal_15501 ;
    wire signal_15502 ;
    wire signal_15503 ;
    wire signal_15504 ;
    wire signal_15505 ;
    wire signal_15506 ;
    wire signal_15507 ;
    wire signal_15508 ;
    wire signal_15509 ;
    wire signal_15510 ;
    wire signal_15511 ;
    wire signal_15512 ;
    wire signal_15513 ;
    wire signal_15514 ;
    wire signal_15515 ;
    wire signal_15516 ;
    wire signal_15517 ;
    wire signal_15518 ;
    wire signal_15519 ;
    wire signal_15520 ;
    wire signal_15521 ;
    wire signal_15522 ;
    wire signal_15523 ;
    wire signal_15524 ;
    wire signal_15525 ;
    wire signal_15526 ;
    wire signal_15527 ;
    wire signal_15528 ;
    wire signal_15529 ;
    wire signal_15530 ;
    wire signal_15531 ;
    wire signal_15532 ;
    wire signal_15533 ;
    wire signal_15534 ;
    wire signal_15535 ;
    wire signal_15536 ;
    wire signal_15537 ;
    wire signal_15538 ;
    wire signal_15539 ;
    wire signal_15540 ;
    wire signal_15541 ;
    wire signal_15542 ;
    wire signal_15543 ;
    wire signal_15544 ;
    wire signal_15545 ;
    wire signal_15546 ;
    wire signal_15547 ;
    wire signal_15548 ;
    wire signal_15549 ;
    wire signal_15550 ;
    wire signal_15551 ;
    wire signal_15552 ;
    wire signal_15553 ;
    wire signal_15554 ;
    wire signal_15555 ;
    wire signal_15556 ;
    wire signal_15557 ;
    wire signal_15558 ;
    wire signal_15559 ;
    wire signal_15560 ;
    wire signal_15561 ;
    wire signal_15562 ;
    wire signal_15563 ;
    wire signal_15564 ;
    wire signal_15565 ;
    wire signal_15566 ;
    wire signal_15567 ;
    wire signal_15568 ;
    wire signal_15569 ;
    wire signal_15570 ;
    wire signal_15571 ;
    wire signal_15572 ;
    wire signal_15573 ;
    wire signal_15574 ;
    wire signal_15575 ;
    wire signal_15576 ;
    wire signal_15577 ;
    wire signal_15578 ;
    wire signal_15579 ;
    wire signal_15580 ;
    wire signal_15581 ;
    wire signal_15582 ;
    wire signal_15583 ;
    wire signal_15584 ;
    wire signal_15585 ;
    wire signal_15586 ;
    wire signal_15587 ;
    wire signal_15588 ;
    wire signal_15589 ;
    wire signal_15590 ;
    wire signal_15591 ;
    wire signal_15592 ;
    wire signal_15593 ;
    wire signal_15594 ;
    wire signal_15595 ;
    wire signal_15596 ;
    wire signal_15597 ;
    wire signal_15598 ;
    wire signal_15599 ;
    wire signal_15600 ;
    wire signal_15601 ;
    wire signal_15602 ;
    wire signal_15603 ;
    wire signal_15604 ;
    wire signal_15605 ;
    wire signal_15606 ;
    wire signal_15607 ;
    wire signal_15608 ;
    wire signal_15609 ;
    wire signal_15610 ;
    wire signal_15611 ;
    wire signal_15612 ;
    wire signal_15613 ;
    wire signal_15614 ;
    wire signal_15615 ;
    wire signal_15616 ;
    wire signal_15617 ;
    wire signal_15618 ;
    wire signal_15619 ;
    wire signal_15620 ;
    wire signal_15621 ;
    wire signal_15622 ;
    wire signal_15623 ;
    wire signal_15624 ;
    wire signal_15625 ;
    wire signal_15626 ;
    wire signal_15627 ;
    wire signal_15628 ;
    wire signal_15629 ;
    wire signal_15630 ;
    wire signal_15631 ;
    wire signal_15632 ;
    wire signal_15633 ;
    wire signal_15634 ;
    wire signal_15635 ;
    wire signal_15636 ;
    wire signal_15637 ;
    wire signal_15638 ;
    wire signal_15639 ;
    wire signal_15640 ;
    wire signal_15641 ;
    wire signal_15642 ;
    wire signal_15643 ;
    wire signal_15644 ;
    wire signal_15645 ;
    wire signal_15646 ;
    wire signal_15647 ;
    wire signal_15648 ;
    wire signal_15649 ;
    wire signal_15650 ;
    wire signal_15651 ;
    wire signal_15652 ;
    wire signal_15653 ;
    wire signal_15654 ;
    wire signal_15655 ;
    wire signal_15656 ;
    wire signal_15657 ;
    wire signal_15658 ;
    wire signal_15659 ;
    wire signal_15660 ;
    wire signal_15661 ;
    wire signal_15662 ;
    wire signal_15663 ;
    wire signal_15664 ;
    wire signal_15665 ;
    wire signal_15666 ;
    wire signal_15667 ;
    wire signal_15668 ;
    wire signal_15669 ;
    wire signal_15670 ;
    wire signal_15671 ;
    wire signal_15672 ;
    wire signal_15673 ;
    wire signal_15674 ;
    wire signal_15675 ;
    wire signal_15676 ;
    wire signal_15677 ;
    wire signal_15678 ;
    wire signal_15679 ;
    wire signal_15680 ;
    wire signal_15681 ;
    wire signal_15682 ;
    wire signal_15683 ;
    wire signal_15684 ;
    wire signal_15685 ;
    wire signal_15686 ;
    wire signal_15687 ;
    wire signal_15688 ;
    wire signal_15689 ;
    wire signal_15690 ;
    wire signal_15691 ;
    wire signal_15692 ;
    wire signal_15693 ;
    wire signal_15694 ;
    wire signal_15695 ;
    wire signal_15696 ;
    wire signal_15697 ;
    wire signal_15698 ;
    wire signal_15699 ;
    wire signal_15700 ;
    wire signal_15701 ;
    wire signal_15702 ;
    wire signal_15703 ;
    wire signal_15704 ;
    wire signal_15705 ;
    wire signal_15706 ;
    wire signal_15707 ;
    wire signal_15708 ;
    wire signal_15709 ;
    wire signal_15710 ;
    wire signal_15711 ;
    wire signal_15712 ;
    wire signal_15713 ;
    wire signal_15714 ;
    wire signal_15715 ;
    wire signal_15716 ;
    wire signal_15717 ;
    wire signal_15718 ;
    wire signal_15719 ;
    wire signal_15720 ;
    wire signal_15721 ;
    wire signal_15722 ;
    wire signal_15723 ;
    wire signal_15724 ;
    wire signal_15725 ;
    wire signal_15726 ;
    wire signal_15727 ;
    wire signal_15728 ;
    wire signal_15729 ;
    wire signal_15730 ;
    wire signal_15731 ;
    wire signal_15732 ;
    wire signal_15733 ;
    wire signal_15734 ;
    wire signal_15735 ;
    wire signal_15736 ;
    wire signal_15737 ;
    wire signal_15738 ;
    wire signal_15739 ;
    wire signal_15740 ;
    wire signal_15741 ;
    wire signal_15742 ;
    wire signal_15743 ;
    wire signal_15744 ;
    wire signal_15745 ;
    wire signal_15746 ;
    wire signal_15747 ;
    wire signal_15748 ;
    wire signal_15749 ;
    wire signal_15750 ;
    wire signal_15751 ;
    wire signal_15752 ;
    wire signal_15753 ;
    wire signal_15754 ;
    wire signal_15755 ;
    wire signal_15756 ;
    wire signal_15757 ;
    wire signal_15758 ;
    wire signal_15759 ;
    wire signal_15760 ;
    wire signal_15761 ;
    wire signal_15762 ;
    wire signal_15763 ;
    wire signal_15764 ;
    wire signal_15765 ;
    wire signal_15766 ;
    wire signal_15767 ;
    wire signal_15768 ;
    wire signal_15769 ;
    wire signal_15770 ;
    wire signal_15771 ;
    wire signal_15772 ;
    wire signal_15773 ;
    wire signal_15774 ;
    wire signal_15775 ;
    wire signal_15776 ;
    wire signal_15777 ;
    wire signal_15778 ;
    wire signal_15779 ;
    wire signal_15780 ;
    wire signal_15781 ;
    wire signal_15782 ;
    wire signal_15783 ;
    wire signal_15784 ;
    wire signal_15785 ;
    wire signal_15786 ;
    wire signal_15787 ;
    wire signal_15788 ;
    wire signal_15789 ;
    wire signal_15790 ;
    wire signal_15791 ;
    wire signal_15792 ;
    wire signal_15793 ;
    wire signal_15794 ;
    wire signal_15795 ;
    wire signal_15796 ;
    wire signal_15797 ;
    wire signal_15798 ;
    wire signal_15799 ;
    wire signal_15800 ;
    wire signal_15801 ;
    wire signal_15802 ;
    wire signal_15803 ;
    wire signal_15804 ;
    wire signal_15805 ;
    wire signal_15806 ;
    wire signal_15807 ;
    wire signal_15808 ;
    wire signal_15809 ;
    wire signal_15810 ;
    wire signal_15811 ;
    wire signal_15812 ;
    wire signal_15813 ;
    wire signal_15814 ;
    wire signal_15815 ;
    wire signal_15816 ;
    wire signal_15817 ;
    wire signal_15818 ;
    wire signal_15819 ;
    wire signal_15820 ;
    wire signal_15821 ;
    wire signal_15822 ;
    wire signal_15823 ;
    wire signal_15824 ;
    wire signal_15825 ;
    wire signal_15826 ;
    wire signal_15827 ;
    wire signal_15828 ;
    wire signal_15829 ;
    wire signal_15830 ;
    wire signal_15831 ;
    wire signal_15832 ;
    wire signal_15833 ;
    wire signal_15834 ;
    wire signal_15835 ;
    wire signal_15836 ;
    wire signal_15837 ;
    wire signal_15838 ;
    wire signal_15839 ;
    wire signal_15840 ;
    wire signal_15841 ;
    wire signal_15842 ;
    wire signal_15843 ;
    wire signal_15844 ;
    wire signal_15845 ;
    wire signal_15846 ;
    wire signal_15847 ;
    wire signal_15848 ;
    wire signal_15849 ;
    wire signal_15850 ;
    wire signal_15851 ;
    wire signal_15852 ;
    wire signal_15853 ;
    wire signal_15854 ;
    wire signal_15855 ;
    wire signal_15856 ;
    wire signal_15857 ;
    wire signal_15858 ;
    wire signal_15859 ;
    wire signal_15860 ;
    wire signal_15861 ;
    wire signal_15862 ;
    wire signal_15863 ;
    wire signal_15864 ;
    wire signal_15865 ;
    wire signal_15866 ;
    wire signal_15867 ;
    wire signal_15868 ;
    wire signal_15869 ;
    wire signal_15870 ;
    wire signal_15871 ;
    wire signal_15872 ;
    wire signal_15873 ;
    wire signal_15874 ;
    wire signal_15875 ;
    wire signal_15876 ;
    wire signal_15877 ;
    wire signal_15878 ;
    wire signal_15879 ;
    wire signal_15880 ;
    wire signal_15881 ;
    wire signal_15882 ;
    wire signal_15883 ;
    wire signal_15884 ;
    wire signal_15885 ;
    wire signal_15886 ;
    wire signal_15887 ;
    wire signal_15888 ;
    wire signal_15889 ;
    wire signal_15890 ;
    wire signal_15891 ;
    wire signal_15892 ;
    wire signal_15893 ;
    wire signal_15894 ;
    wire signal_15895 ;
    wire signal_15896 ;
    wire signal_15897 ;
    wire signal_15898 ;
    wire signal_15899 ;
    wire signal_15900 ;
    wire signal_15901 ;
    wire signal_15902 ;
    wire signal_15903 ;
    wire signal_15904 ;
    wire signal_15905 ;
    wire signal_15906 ;
    wire signal_15907 ;
    wire signal_15908 ;
    wire signal_15909 ;
    wire signal_15910 ;
    wire signal_15911 ;
    wire signal_15912 ;
    wire signal_15913 ;
    wire signal_15914 ;
    wire signal_15915 ;
    wire signal_15916 ;
    wire signal_15917 ;
    wire signal_15918 ;
    wire signal_15919 ;
    wire signal_15920 ;
    wire signal_15921 ;
    wire signal_15922 ;
    wire signal_15923 ;
    wire signal_15924 ;
    wire signal_15925 ;
    wire signal_15926 ;
    wire signal_15927 ;
    wire signal_15928 ;
    wire signal_15929 ;
    wire signal_15930 ;
    wire signal_15931 ;
    wire signal_15932 ;
    wire signal_15933 ;
    wire signal_15934 ;
    wire signal_15935 ;
    wire signal_15936 ;
    wire signal_15937 ;
    wire signal_15938 ;
    wire signal_15939 ;
    wire signal_15940 ;
    wire signal_15941 ;
    wire signal_15942 ;
    wire signal_15943 ;
    wire signal_15944 ;
    wire signal_15945 ;
    wire signal_15946 ;
    wire signal_15947 ;
    wire signal_15948 ;
    wire signal_15949 ;
    wire signal_15950 ;
    wire signal_15951 ;
    wire signal_15952 ;
    wire signal_15953 ;
    wire signal_15954 ;
    wire signal_15955 ;
    wire signal_15956 ;
    wire signal_15957 ;
    wire signal_15958 ;
    wire signal_15959 ;
    wire signal_15960 ;
    wire signal_15961 ;
    wire signal_15962 ;
    wire signal_15963 ;
    wire signal_15964 ;
    wire signal_15965 ;
    wire signal_15966 ;
    wire signal_15967 ;
    wire signal_15968 ;
    wire signal_15969 ;
    wire signal_15970 ;
    wire signal_15971 ;
    wire signal_15972 ;
    wire signal_15973 ;
    wire signal_15974 ;
    wire signal_15975 ;
    wire signal_15976 ;
    wire signal_15977 ;
    wire signal_15978 ;
    wire signal_15979 ;
    wire signal_15980 ;
    wire signal_15981 ;
    wire signal_15982 ;
    wire signal_15983 ;
    wire signal_15984 ;
    wire signal_15985 ;
    wire signal_15986 ;
    wire signal_15987 ;
    wire signal_15988 ;
    wire signal_15989 ;
    wire signal_15990 ;
    wire signal_15991 ;
    wire signal_15992 ;
    wire signal_15993 ;
    wire signal_15994 ;
    wire signal_15995 ;
    wire signal_15996 ;
    wire signal_15997 ;
    wire signal_15998 ;
    wire signal_15999 ;
    wire signal_16000 ;
    wire signal_16001 ;
    wire signal_16002 ;
    wire signal_16003 ;
    wire signal_16004 ;
    wire signal_16005 ;
    wire signal_16006 ;
    wire signal_16007 ;
    wire signal_16008 ;
    wire signal_16009 ;
    wire signal_16010 ;
    wire signal_16011 ;
    wire signal_16012 ;
    wire signal_16013 ;
    wire signal_16014 ;
    wire signal_16015 ;
    wire signal_16016 ;
    wire signal_16017 ;
    wire signal_16018 ;
    wire signal_16019 ;
    wire signal_16020 ;
    wire signal_16021 ;
    wire signal_16022 ;
    wire signal_16023 ;
    wire signal_16024 ;
    wire signal_16025 ;
    wire signal_16026 ;
    wire signal_16027 ;
    wire signal_16028 ;
    wire signal_16029 ;
    wire signal_16030 ;
    wire signal_16031 ;
    wire signal_16032 ;
    wire signal_16033 ;
    wire signal_16034 ;
    wire signal_16035 ;
    wire signal_16036 ;
    wire signal_16037 ;
    wire signal_16038 ;
    wire signal_16039 ;
    wire signal_16040 ;
    wire signal_16041 ;
    wire signal_16042 ;
    wire signal_16043 ;
    wire signal_16044 ;
    wire signal_16045 ;
    wire signal_16046 ;
    wire signal_16047 ;
    wire signal_16048 ;
    wire signal_16049 ;
    wire signal_16050 ;
    wire signal_16051 ;
    wire signal_16052 ;
    wire signal_16053 ;
    wire signal_16054 ;
    wire signal_16055 ;
    wire signal_16056 ;
    wire signal_16057 ;
    wire signal_16058 ;
    wire signal_16059 ;
    wire signal_16060 ;
    wire signal_16061 ;
    wire signal_16062 ;
    wire signal_16063 ;
    wire signal_16064 ;
    wire signal_16065 ;
    wire signal_16066 ;
    wire signal_16067 ;
    wire signal_16068 ;
    wire signal_16069 ;
    wire signal_16070 ;
    wire signal_16071 ;
    wire signal_16072 ;
    wire signal_16073 ;
    wire signal_16074 ;
    wire signal_16075 ;
    wire signal_16076 ;
    wire signal_16077 ;
    wire signal_16078 ;
    wire signal_16079 ;
    wire signal_16080 ;
    wire signal_16081 ;
    wire signal_16082 ;
    wire signal_16083 ;
    wire signal_16084 ;
    wire signal_16085 ;
    wire signal_16086 ;
    wire signal_16087 ;
    wire signal_16088 ;
    wire signal_16089 ;
    wire signal_16090 ;
    wire signal_16091 ;
    wire signal_16092 ;
    wire signal_16093 ;
    wire signal_16094 ;
    wire signal_16095 ;
    wire signal_16096 ;
    wire signal_16097 ;
    wire signal_16098 ;
    wire signal_16099 ;
    wire signal_16100 ;
    wire signal_16101 ;
    wire signal_16102 ;
    wire signal_16103 ;
    wire signal_16104 ;
    wire signal_16105 ;
    wire signal_16106 ;
    wire signal_16107 ;
    wire signal_16108 ;
    wire signal_16109 ;
    wire signal_16110 ;
    wire signal_16111 ;
    wire signal_16112 ;
    wire signal_16113 ;
    wire signal_16114 ;
    wire signal_16115 ;
    wire signal_16116 ;
    wire signal_16117 ;
    wire signal_16118 ;
    wire signal_16119 ;
    wire signal_16120 ;
    wire signal_16121 ;
    wire signal_16122 ;
    wire signal_16123 ;
    wire signal_16124 ;
    wire signal_16125 ;
    wire signal_16126 ;
    wire signal_16127 ;
    wire signal_16128 ;
    wire signal_16129 ;
    wire signal_16130 ;
    wire signal_16131 ;
    wire signal_16132 ;
    wire signal_16133 ;
    wire signal_16134 ;
    wire signal_16135 ;
    wire signal_16136 ;
    wire signal_16137 ;
    wire signal_16138 ;
    wire signal_16139 ;
    wire signal_16140 ;
    wire signal_16141 ;
    wire signal_16142 ;
    wire signal_16143 ;
    wire signal_16144 ;
    wire signal_16145 ;
    wire signal_16146 ;
    wire signal_16147 ;
    wire signal_16148 ;
    wire signal_16149 ;
    wire signal_16150 ;
    wire signal_16151 ;
    wire signal_16152 ;
    wire signal_16153 ;
    wire signal_16154 ;
    wire signal_16155 ;
    wire signal_16156 ;
    wire signal_16157 ;
    wire signal_16158 ;
    wire signal_16159 ;
    wire signal_16160 ;
    wire signal_16161 ;
    wire signal_16162 ;
    wire signal_16163 ;
    wire signal_16164 ;
    wire signal_16165 ;
    wire signal_16166 ;
    wire signal_16167 ;
    wire signal_16168 ;
    wire signal_16169 ;
    wire signal_16170 ;
    wire signal_16171 ;
    wire signal_16172 ;
    wire signal_16173 ;
    wire signal_16174 ;
    wire signal_16175 ;
    wire signal_16176 ;
    wire signal_16177 ;
    wire signal_16178 ;
    wire signal_16179 ;
    wire signal_16180 ;
    wire signal_16181 ;
    wire signal_16182 ;
    wire signal_16183 ;
    wire signal_16184 ;
    wire signal_16185 ;
    wire signal_16186 ;
    wire signal_16187 ;
    wire signal_16188 ;
    wire signal_16189 ;
    wire signal_16190 ;
    wire signal_16191 ;
    wire signal_16192 ;
    wire signal_16193 ;
    wire signal_16194 ;
    wire signal_16195 ;
    wire signal_16196 ;
    wire signal_16197 ;
    wire signal_16198 ;
    wire signal_16199 ;
    wire signal_16200 ;
    wire signal_16201 ;
    wire signal_16202 ;
    wire signal_16203 ;
    wire signal_16204 ;
    wire signal_16205 ;
    wire signal_16206 ;
    wire signal_16207 ;
    wire signal_16208 ;
    wire signal_16209 ;
    wire signal_16210 ;
    wire signal_16211 ;
    wire signal_16212 ;
    wire signal_16213 ;
    wire signal_16214 ;
    wire signal_16215 ;
    wire signal_16216 ;
    wire signal_16217 ;
    wire signal_16218 ;
    wire signal_16219 ;
    wire signal_16220 ;
    wire signal_16221 ;
    wire signal_16222 ;
    wire signal_16223 ;
    wire signal_16224 ;
    wire signal_16225 ;
    wire signal_16226 ;
    wire signal_16227 ;
    wire signal_16228 ;
    wire signal_16229 ;
    wire signal_16230 ;
    wire signal_16231 ;
    wire signal_16232 ;
    wire signal_16233 ;
    wire signal_16234 ;
    wire signal_16235 ;
    wire signal_16236 ;
    wire signal_16237 ;
    wire signal_16238 ;
    wire signal_16239 ;
    wire signal_16240 ;
    wire signal_16241 ;
    wire signal_16242 ;
    wire signal_16243 ;
    wire signal_16244 ;
    wire signal_16245 ;
    wire signal_16246 ;
    wire signal_16247 ;
    wire signal_16248 ;
    wire signal_16249 ;
    wire signal_16250 ;
    wire signal_16251 ;
    wire signal_16252 ;
    wire signal_16253 ;
    wire signal_16254 ;
    wire signal_16255 ;
    wire signal_16256 ;
    wire signal_16257 ;
    wire signal_16258 ;
    wire signal_16259 ;
    wire signal_16260 ;
    wire signal_16261 ;
    wire signal_16262 ;
    wire signal_16263 ;
    wire signal_16264 ;
    wire signal_16265 ;
    wire signal_16266 ;
    wire signal_16267 ;
    wire signal_16268 ;
    wire signal_16269 ;
    wire signal_16270 ;
    wire signal_16271 ;
    wire signal_16272 ;
    wire signal_16273 ;
    wire signal_16274 ;
    wire signal_16275 ;
    wire signal_16276 ;
    wire signal_16277 ;
    wire signal_16278 ;
    wire signal_16279 ;
    wire signal_16280 ;
    wire signal_16281 ;
    wire signal_16282 ;
    wire signal_16283 ;
    wire signal_16284 ;
    wire signal_16285 ;
    wire signal_16286 ;
    wire signal_16287 ;
    wire signal_16288 ;
    wire signal_16289 ;
    wire signal_16290 ;
    wire signal_16291 ;
    wire signal_16292 ;
    wire signal_16293 ;
    wire signal_16294 ;
    wire signal_16295 ;
    wire signal_16296 ;
    wire signal_16297 ;
    wire signal_16298 ;
    wire signal_16299 ;
    wire signal_16300 ;
    wire signal_16301 ;
    wire signal_16302 ;
    wire signal_16303 ;
    wire signal_16304 ;
    wire signal_16305 ;
    wire signal_16306 ;
    wire signal_16307 ;
    wire signal_16308 ;
    wire signal_16309 ;
    wire signal_16310 ;
    wire signal_16311 ;
    wire signal_16312 ;
    wire signal_16313 ;
    wire signal_16314 ;
    wire signal_16315 ;
    wire signal_16316 ;
    wire signal_16317 ;
    wire signal_16318 ;
    wire signal_16319 ;
    wire signal_16320 ;
    wire signal_16321 ;
    wire signal_16322 ;
    wire signal_16323 ;
    wire signal_16324 ;
    wire signal_16325 ;
    wire signal_16326 ;
    wire signal_16327 ;
    wire signal_16328 ;
    wire signal_16329 ;
    wire signal_16330 ;
    wire signal_16331 ;
    wire signal_16332 ;
    wire signal_16333 ;
    wire signal_16334 ;
    wire signal_16335 ;
    wire signal_16336 ;
    wire signal_16337 ;
    wire signal_16338 ;
    wire signal_16339 ;
    wire signal_16340 ;
    wire signal_16341 ;
    wire signal_16342 ;
    wire signal_16343 ;
    wire signal_16344 ;
    wire signal_16345 ;
    wire signal_16346 ;
    wire signal_16347 ;
    wire signal_16348 ;
    wire signal_16349 ;
    wire signal_16350 ;
    wire signal_16351 ;
    wire signal_16352 ;
    wire signal_16353 ;
    wire signal_16354 ;
    wire signal_16355 ;
    wire signal_16356 ;
    wire signal_16357 ;
    wire signal_16358 ;
    wire signal_16359 ;
    wire signal_16360 ;
    wire signal_16361 ;
    wire signal_16362 ;
    wire signal_16363 ;
    wire signal_16364 ;
    wire signal_16365 ;
    wire signal_16366 ;
    wire signal_16367 ;
    wire signal_16368 ;
    wire signal_16369 ;
    wire signal_16370 ;
    wire signal_16371 ;
    wire signal_16372 ;
    wire signal_16373 ;
    wire signal_16374 ;
    wire signal_16375 ;
    wire signal_16376 ;
    wire signal_16377 ;
    wire signal_16378 ;
    wire signal_16379 ;
    wire signal_16380 ;
    wire signal_16381 ;
    wire signal_16382 ;
    wire signal_16383 ;
    wire signal_16384 ;
    wire signal_16385 ;
    wire signal_16386 ;
    wire signal_16387 ;
    wire signal_16388 ;
    wire signal_16389 ;
    wire signal_16390 ;
    wire signal_16391 ;
    wire signal_16392 ;
    wire signal_16393 ;
    wire signal_16394 ;
    wire signal_16395 ;
    wire signal_16396 ;
    wire signal_16397 ;
    wire signal_16398 ;
    wire signal_16399 ;
    wire signal_16400 ;
    wire signal_16401 ;
    wire signal_16402 ;
    wire signal_16403 ;
    wire signal_16404 ;
    wire signal_16405 ;
    wire signal_16406 ;
    wire signal_16407 ;
    wire signal_16408 ;
    wire signal_16409 ;
    wire signal_16410 ;
    wire signal_16411 ;
    wire signal_16412 ;
    wire signal_16413 ;
    wire signal_16414 ;
    wire signal_16415 ;
    wire signal_16416 ;
    wire signal_16417 ;
    wire signal_16418 ;
    wire signal_16419 ;
    wire signal_16420 ;
    wire signal_16421 ;
    wire signal_16422 ;
    wire signal_16423 ;
    wire signal_16424 ;
    wire signal_16425 ;
    wire signal_16426 ;
    wire signal_16427 ;
    wire signal_16428 ;
    wire signal_16429 ;
    wire signal_16430 ;
    wire signal_16431 ;
    wire signal_16432 ;
    wire signal_16433 ;
    wire signal_16434 ;
    wire signal_16435 ;
    wire signal_16436 ;
    wire signal_16437 ;
    wire signal_16438 ;
    wire signal_16439 ;
    wire signal_16440 ;
    wire signal_16441 ;
    wire signal_16442 ;
    wire signal_16443 ;
    wire signal_16444 ;
    wire signal_16445 ;
    wire signal_16446 ;
    wire signal_16447 ;
    wire signal_16448 ;
    wire signal_16449 ;
    wire signal_16450 ;
    wire signal_16451 ;
    wire signal_16452 ;
    wire signal_16453 ;
    wire signal_16454 ;
    wire signal_16455 ;
    wire signal_16456 ;
    wire signal_16457 ;
    wire signal_16458 ;
    wire signal_16459 ;
    wire signal_16460 ;
    wire signal_16461 ;
    wire signal_16462 ;
    wire signal_16463 ;
    wire signal_16464 ;
    wire signal_16465 ;
    wire signal_16466 ;
    wire signal_16467 ;
    wire signal_16468 ;
    wire signal_16469 ;
    wire signal_16470 ;
    wire signal_16471 ;
    wire signal_16472 ;
    wire signal_16473 ;
    wire signal_16474 ;
    wire signal_16475 ;
    wire signal_16476 ;
    wire signal_16477 ;
    wire signal_16478 ;
    wire signal_16479 ;
    wire signal_16480 ;
    wire signal_16481 ;
    wire signal_16482 ;
    wire signal_16483 ;
    wire signal_16484 ;
    wire signal_16485 ;
    wire signal_16486 ;
    wire signal_16487 ;
    wire signal_16488 ;
    wire signal_16489 ;
    wire signal_16490 ;
    wire signal_16491 ;
    wire signal_16492 ;
    wire signal_16493 ;
    wire signal_16494 ;
    wire signal_16495 ;
    wire signal_16496 ;
    wire signal_16497 ;
    wire signal_16498 ;
    wire signal_16499 ;
    wire signal_16500 ;
    wire signal_16501 ;
    wire signal_16502 ;
    wire signal_16503 ;
    wire signal_16504 ;
    wire signal_16505 ;
    wire signal_16506 ;
    wire signal_16507 ;
    wire signal_16508 ;
    wire signal_16509 ;
    wire signal_16510 ;
    wire signal_16511 ;
    wire signal_16512 ;
    wire signal_16513 ;
    wire signal_16514 ;
    wire signal_16515 ;
    wire signal_16516 ;
    wire signal_16517 ;
    wire signal_16518 ;
    wire signal_16519 ;
    wire signal_16520 ;
    wire signal_16521 ;
    wire signal_16522 ;
    wire signal_16523 ;
    wire signal_16524 ;
    wire signal_16525 ;
    wire signal_16526 ;
    wire signal_16527 ;
    wire signal_16528 ;
    wire signal_16529 ;
    wire signal_16530 ;
    wire signal_16531 ;
    wire signal_16532 ;
    wire signal_16533 ;
    wire signal_16534 ;
    wire signal_16535 ;
    wire signal_16536 ;
    wire signal_16537 ;
    wire signal_16538 ;
    wire signal_16539 ;
    wire signal_16540 ;
    wire signal_16541 ;
    wire signal_16542 ;
    wire signal_16543 ;
    wire signal_16544 ;
    wire signal_16545 ;
    wire signal_16546 ;
    wire signal_16547 ;
    wire signal_16548 ;
    wire signal_16549 ;
    wire signal_16550 ;
    wire signal_16551 ;
    wire signal_16552 ;
    wire signal_16553 ;
    wire signal_16554 ;
    wire signal_16555 ;
    wire signal_16556 ;
    wire signal_16557 ;
    wire signal_16558 ;
    wire signal_16559 ;
    wire signal_16560 ;
    wire signal_16561 ;
    wire signal_16562 ;
    wire signal_16563 ;
    wire signal_16564 ;
    wire signal_16565 ;
    wire signal_16566 ;
    wire signal_16567 ;
    wire signal_16568 ;
    wire signal_16569 ;
    wire signal_16570 ;
    wire signal_16571 ;
    wire signal_16572 ;
    wire signal_16573 ;
    wire signal_16574 ;
    wire signal_16575 ;
    wire signal_16576 ;
    wire signal_16577 ;
    wire signal_16578 ;
    wire signal_16579 ;
    wire signal_16580 ;
    wire signal_16581 ;
    wire signal_16582 ;
    wire signal_16583 ;
    wire signal_16584 ;
    wire signal_16585 ;
    wire signal_16586 ;
    wire signal_16587 ;
    wire signal_16588 ;
    wire signal_16589 ;
    wire signal_16590 ;
    wire signal_16591 ;
    wire signal_16592 ;
    wire signal_16593 ;
    wire signal_16594 ;
    wire signal_16595 ;
    wire signal_16596 ;
    wire signal_16597 ;
    wire signal_16598 ;
    wire signal_16599 ;
    wire signal_16600 ;
    wire signal_16601 ;
    wire signal_16602 ;
    wire signal_16603 ;
    wire signal_16604 ;
    wire signal_16605 ;
    wire signal_16606 ;
    wire signal_16607 ;
    wire signal_16608 ;
    wire signal_16609 ;
    wire signal_16610 ;
    wire signal_16611 ;
    wire signal_16612 ;
    wire signal_16613 ;
    wire signal_16614 ;
    wire signal_16615 ;
    wire signal_16616 ;
    wire signal_16617 ;
    wire signal_16618 ;
    wire signal_16619 ;
    wire signal_16620 ;
    wire signal_16621 ;
    wire signal_16622 ;
    wire signal_16623 ;
    wire signal_16624 ;
    wire signal_16625 ;
    wire signal_16626 ;
    wire signal_16627 ;
    wire signal_16628 ;
    wire signal_16629 ;
    wire signal_16630 ;
    wire signal_16631 ;
    wire signal_16632 ;
    wire signal_16633 ;
    wire signal_16634 ;
    wire signal_16635 ;
    wire signal_16636 ;
    wire signal_16637 ;
    wire signal_16638 ;
    wire signal_16639 ;
    wire signal_16640 ;
    wire signal_16641 ;
    wire signal_16642 ;
    wire signal_16643 ;
    wire signal_16644 ;
    wire signal_16645 ;
    wire signal_16646 ;
    wire signal_16647 ;
    wire signal_16648 ;
    wire signal_16649 ;
    wire signal_16650 ;
    wire signal_16651 ;
    wire signal_16652 ;
    wire signal_16653 ;
    wire signal_16654 ;
    wire signal_16655 ;
    wire signal_16656 ;
    wire signal_16657 ;
    wire signal_16658 ;
    wire signal_16659 ;
    wire signal_16660 ;
    wire signal_16661 ;
    wire signal_16662 ;
    wire signal_16663 ;
    wire signal_16664 ;
    wire signal_16665 ;
    wire signal_16666 ;
    wire signal_16667 ;
    wire signal_16668 ;
    wire signal_16669 ;
    wire signal_16670 ;
    wire signal_16671 ;
    wire signal_16672 ;
    wire signal_16673 ;
    wire signal_16674 ;
    wire signal_16675 ;
    wire signal_16676 ;
    wire signal_16677 ;
    wire signal_16678 ;
    wire signal_16679 ;
    wire signal_16680 ;
    wire signal_16681 ;
    wire signal_16682 ;
    wire signal_16683 ;
    wire signal_16684 ;
    wire signal_16685 ;
    wire signal_16686 ;
    wire signal_16687 ;
    wire signal_16688 ;
    wire signal_16689 ;
    wire signal_16690 ;
    wire signal_16691 ;
    wire signal_16692 ;
    wire signal_16693 ;
    wire signal_16694 ;
    wire signal_16695 ;
    wire signal_16696 ;
    wire signal_16697 ;
    wire signal_16698 ;
    wire signal_16699 ;
    wire signal_16700 ;
    wire signal_16701 ;
    wire signal_16702 ;
    wire signal_16703 ;
    wire signal_16704 ;
    wire signal_16705 ;
    wire signal_16706 ;
    wire signal_16707 ;
    wire signal_16708 ;
    wire signal_16709 ;
    wire signal_16710 ;
    wire signal_16711 ;
    wire signal_16712 ;
    wire signal_16713 ;
    wire signal_16714 ;
    wire signal_16715 ;
    wire signal_16716 ;
    wire signal_16717 ;
    wire signal_16718 ;
    wire signal_16719 ;
    wire signal_16720 ;
    wire signal_16721 ;
    wire signal_16722 ;
    wire signal_16723 ;
    wire signal_16724 ;
    wire signal_16725 ;
    wire signal_16726 ;
    wire signal_16727 ;
    wire signal_16728 ;
    wire signal_16729 ;
    wire signal_16730 ;
    wire signal_16731 ;
    wire signal_16732 ;
    wire signal_16733 ;
    wire signal_16734 ;
    wire signal_16735 ;
    wire signal_16736 ;
    wire signal_16737 ;
    wire signal_16738 ;
    wire signal_16739 ;
    wire signal_16740 ;
    wire signal_16741 ;
    wire signal_16742 ;
    wire signal_16743 ;
    wire signal_16744 ;
    wire signal_16745 ;
    wire signal_16746 ;
    wire signal_16747 ;
    wire signal_16748 ;
    wire signal_16749 ;
    wire signal_16750 ;
    wire signal_16751 ;
    wire signal_16752 ;
    wire signal_16753 ;
    wire signal_16754 ;
    wire signal_16755 ;
    wire signal_16756 ;
    wire signal_16757 ;
    wire signal_16758 ;
    wire signal_16759 ;
    wire signal_16760 ;
    wire signal_16761 ;
    wire signal_16762 ;
    wire signal_16763 ;
    wire signal_16764 ;
    wire signal_16765 ;
    wire signal_16766 ;
    wire signal_16767 ;
    wire signal_16768 ;
    wire signal_16769 ;
    wire signal_16770 ;
    wire signal_16771 ;
    wire signal_16772 ;
    wire signal_16773 ;
    wire signal_16774 ;
    wire signal_16775 ;
    wire signal_16776 ;
    wire signal_16777 ;
    wire signal_16778 ;
    wire signal_16779 ;
    wire signal_16780 ;
    wire signal_16781 ;
    wire signal_16782 ;
    wire signal_16783 ;
    wire signal_16784 ;
    wire signal_16785 ;
    wire signal_16786 ;
    wire signal_16787 ;
    wire signal_16788 ;
    wire signal_16789 ;
    wire signal_16790 ;
    wire signal_16791 ;
    wire signal_16792 ;
    wire signal_16793 ;
    wire signal_16794 ;
    wire signal_16795 ;
    wire signal_16796 ;
    wire signal_16797 ;
    wire signal_16798 ;
    wire signal_16799 ;
    wire signal_16800 ;
    wire signal_16801 ;
    wire signal_16802 ;
    wire signal_16803 ;
    wire signal_16804 ;
    wire signal_16805 ;
    wire signal_16806 ;
    wire signal_16807 ;
    wire signal_16808 ;
    wire signal_16809 ;
    wire signal_16810 ;
    wire signal_16811 ;
    wire signal_16812 ;
    wire signal_16813 ;
    wire signal_16814 ;
    wire signal_16815 ;
    wire signal_16816 ;
    wire signal_16817 ;
    wire signal_16818 ;
    wire signal_16819 ;
    wire signal_16820 ;
    wire signal_16821 ;
    wire signal_16822 ;
    wire signal_16823 ;
    wire signal_16824 ;
    wire signal_16825 ;
    wire signal_16826 ;
    wire signal_16827 ;
    wire signal_16828 ;
    wire signal_16829 ;
    wire signal_16830 ;
    wire signal_16831 ;
    wire signal_16832 ;
    wire signal_16833 ;
    wire signal_16834 ;
    wire signal_16835 ;
    wire signal_16836 ;
    wire signal_16837 ;
    wire signal_16838 ;
    wire signal_16839 ;
    wire signal_16840 ;
    wire signal_16841 ;
    wire signal_16842 ;
    wire signal_16843 ;
    wire signal_16844 ;
    wire signal_16845 ;
    wire signal_16846 ;
    wire signal_16847 ;
    wire signal_16848 ;
    wire signal_16849 ;
    wire signal_16850 ;
    wire signal_16851 ;
    wire signal_16852 ;
    wire signal_16853 ;
    wire signal_16854 ;
    wire signal_16855 ;
    wire signal_16856 ;
    wire signal_16857 ;
    wire signal_16858 ;
    wire signal_16859 ;
    wire signal_16860 ;
    wire signal_16861 ;
    wire signal_16862 ;
    wire signal_16863 ;
    wire signal_16864 ;
    wire signal_16865 ;
    wire signal_16866 ;
    wire signal_16867 ;
    wire signal_16868 ;
    wire signal_16869 ;
    wire signal_16870 ;
    wire signal_16871 ;
    wire signal_16872 ;
    wire signal_16873 ;
    wire signal_16874 ;
    wire signal_16875 ;
    wire signal_16876 ;
    wire signal_16877 ;
    wire signal_16878 ;
    wire signal_16879 ;
    wire signal_16880 ;
    wire signal_16881 ;
    wire signal_16882 ;
    wire signal_16883 ;
    wire signal_16884 ;
    wire signal_16885 ;
    wire signal_16886 ;
    wire signal_16887 ;
    wire signal_16888 ;
    wire signal_16889 ;
    wire signal_16890 ;
    wire signal_16891 ;
    wire signal_16892 ;
    wire signal_16893 ;
    wire signal_16894 ;
    wire signal_16895 ;
    wire signal_16896 ;
    wire signal_16897 ;
    wire signal_16898 ;
    wire signal_16899 ;
    wire signal_16900 ;
    wire signal_16901 ;
    wire signal_16902 ;
    wire signal_16903 ;
    wire signal_16904 ;
    wire signal_16905 ;
    wire signal_16906 ;
    wire signal_16907 ;
    wire signal_16908 ;
    wire signal_16909 ;
    wire signal_16910 ;
    wire signal_16911 ;
    wire signal_16912 ;
    wire signal_16913 ;
    wire signal_16914 ;
    wire signal_16915 ;
    wire signal_16916 ;
    wire signal_16917 ;
    wire signal_16918 ;
    wire signal_16919 ;
    wire signal_16920 ;
    wire signal_16921 ;
    wire signal_16922 ;
    wire signal_16923 ;
    wire signal_16924 ;
    wire signal_16925 ;
    wire signal_16926 ;
    wire signal_16927 ;
    wire signal_16928 ;
    wire signal_16929 ;
    wire signal_16930 ;
    wire signal_16931 ;
    wire signal_16932 ;
    wire signal_16933 ;
    wire signal_16934 ;
    wire signal_16935 ;
    wire signal_16936 ;
    wire signal_16937 ;
    wire signal_16938 ;
    wire signal_16939 ;
    wire signal_16940 ;
    wire signal_16941 ;
    wire signal_16942 ;
    wire signal_16943 ;
    wire signal_16944 ;
    wire signal_16945 ;
    wire signal_16946 ;
    wire signal_16947 ;
    wire signal_16948 ;
    wire signal_16949 ;
    wire signal_16950 ;
    wire signal_16951 ;
    wire signal_16952 ;
    wire signal_16953 ;
    wire signal_16954 ;
    wire signal_16955 ;
    wire signal_16956 ;
    wire signal_16957 ;
    wire signal_16958 ;
    wire signal_16959 ;
    wire signal_16960 ;
    wire signal_16961 ;
    wire signal_16962 ;
    wire signal_16963 ;
    wire signal_16964 ;
    wire signal_16965 ;
    wire signal_16966 ;
    wire signal_16967 ;
    wire signal_16968 ;
    wire signal_16969 ;
    wire signal_16970 ;
    wire signal_16971 ;
    wire signal_16972 ;
    wire signal_16973 ;
    wire signal_16974 ;
    wire signal_16975 ;
    wire signal_16976 ;
    wire signal_16977 ;
    wire signal_16978 ;
    wire signal_16979 ;
    wire signal_16980 ;
    wire signal_16981 ;
    wire signal_16982 ;
    wire signal_16983 ;
    wire signal_16984 ;
    wire signal_16985 ;
    wire signal_16986 ;
    wire signal_16987 ;
    wire signal_16988 ;
    wire signal_16989 ;
    wire signal_16990 ;
    wire signal_16991 ;
    wire signal_16992 ;
    wire signal_16993 ;
    wire signal_16994 ;
    wire signal_16995 ;
    wire signal_16996 ;
    wire signal_16997 ;
    wire signal_16998 ;
    wire signal_16999 ;
    wire signal_17000 ;
    wire signal_17001 ;
    wire signal_17002 ;
    wire signal_17003 ;
    wire signal_17004 ;
    wire signal_17005 ;
    wire signal_17006 ;
    wire signal_17007 ;
    wire signal_17008 ;
    wire signal_17009 ;
    wire signal_17010 ;
    wire signal_17011 ;
    wire signal_17012 ;
    wire signal_17013 ;
    wire signal_17014 ;
    wire signal_17015 ;
    wire signal_17016 ;
    wire signal_17017 ;
    wire signal_17018 ;
    wire signal_17019 ;
    wire signal_17020 ;
    wire signal_17021 ;
    wire signal_17022 ;
    wire signal_17023 ;
    wire signal_17024 ;
    wire signal_17025 ;
    wire signal_17026 ;
    wire signal_17027 ;
    wire signal_17028 ;
    wire signal_17029 ;
    wire signal_17030 ;
    wire signal_17031 ;
    wire signal_17032 ;
    wire signal_17033 ;
    wire signal_17034 ;
    wire signal_17035 ;
    wire signal_17036 ;
    wire signal_17037 ;
    wire signal_17038 ;
    wire signal_17039 ;
    wire signal_17040 ;
    wire signal_17041 ;
    wire signal_17042 ;
    wire signal_17043 ;
    wire signal_17044 ;
    wire signal_17045 ;
    wire signal_17046 ;
    wire signal_17047 ;
    wire signal_17048 ;
    wire signal_17049 ;
    wire signal_17050 ;
    wire signal_17051 ;
    wire signal_17052 ;
    wire signal_17053 ;
    wire signal_17054 ;
    wire signal_17055 ;
    wire signal_17056 ;
    wire signal_17057 ;
    wire signal_17058 ;
    wire signal_17059 ;
    wire signal_17060 ;
    wire signal_17061 ;
    wire signal_17062 ;
    wire signal_17063 ;
    wire signal_17064 ;
    wire signal_17065 ;
    wire signal_17066 ;
    wire signal_17067 ;
    wire signal_17068 ;
    wire signal_17069 ;
    wire signal_17070 ;
    wire signal_17071 ;
    wire signal_17072 ;
    wire signal_17073 ;
    wire signal_17074 ;
    wire signal_17075 ;
    wire signal_17076 ;
    wire signal_17077 ;
    wire signal_17078 ;
    wire signal_17079 ;
    wire signal_17080 ;
    wire signal_17081 ;
    wire signal_17082 ;
    wire signal_17083 ;
    wire signal_17084 ;
    wire signal_17085 ;
    wire signal_17086 ;
    wire signal_17087 ;
    wire signal_17088 ;
    wire signal_17089 ;
    wire signal_17090 ;
    wire signal_17091 ;
    wire signal_17092 ;
    wire signal_17093 ;
    wire signal_17094 ;
    wire signal_17095 ;
    wire signal_17096 ;
    wire signal_17097 ;
    wire signal_17098 ;
    wire signal_17099 ;
    wire signal_17100 ;
    wire signal_17101 ;
    wire signal_17102 ;
    wire signal_17103 ;
    wire signal_17104 ;
    wire signal_17105 ;
    wire signal_17106 ;
    wire signal_17107 ;
    wire signal_17108 ;
    wire signal_17109 ;
    wire signal_17110 ;
    wire signal_17111 ;
    wire signal_17112 ;
    wire signal_17113 ;
    wire signal_17114 ;
    wire signal_17115 ;
    wire signal_17116 ;
    wire signal_17117 ;
    wire signal_17118 ;
    wire signal_17119 ;
    wire signal_17120 ;
    wire signal_17121 ;
    wire signal_17122 ;
    wire signal_17123 ;
    wire signal_17124 ;
    wire signal_17125 ;
    wire signal_17126 ;
    wire signal_17127 ;
    wire signal_17128 ;
    wire signal_17129 ;
    wire signal_17130 ;
    wire signal_17131 ;
    wire signal_17132 ;
    wire signal_17133 ;
    wire signal_17134 ;
    wire signal_17135 ;
    wire signal_17136 ;
    wire signal_17137 ;
    wire signal_17138 ;
    wire signal_17139 ;
    wire signal_17140 ;
    wire signal_17141 ;
    wire signal_17142 ;
    wire signal_17143 ;
    wire signal_17144 ;
    wire signal_17145 ;
    wire signal_17146 ;
    wire signal_17147 ;
    wire signal_17148 ;
    wire signal_17149 ;
    wire signal_17150 ;
    wire signal_17151 ;
    wire signal_17152 ;
    wire signal_17153 ;
    wire signal_17154 ;
    wire signal_17155 ;
    wire signal_17156 ;
    wire signal_17157 ;
    wire signal_17158 ;
    wire signal_17159 ;
    wire signal_17160 ;
    wire signal_17161 ;
    wire signal_17162 ;
    wire signal_17163 ;
    wire signal_17164 ;
    wire signal_17165 ;
    wire signal_17166 ;
    wire signal_17167 ;
    wire signal_17168 ;
    wire signal_17169 ;
    wire signal_17170 ;
    wire signal_17171 ;
    wire signal_17172 ;
    wire signal_17173 ;
    wire signal_17174 ;
    wire signal_17175 ;
    wire signal_17176 ;
    wire signal_17177 ;
    wire signal_17178 ;
    wire signal_17179 ;
    wire signal_17180 ;
    wire signal_17181 ;
    wire signal_17182 ;
    wire signal_17183 ;
    wire signal_17184 ;
    wire signal_17185 ;
    wire signal_17186 ;
    wire signal_17187 ;
    wire signal_17188 ;
    wire signal_17189 ;
    wire signal_17190 ;
    wire signal_17191 ;
    wire signal_17192 ;
    wire signal_17193 ;
    wire signal_17194 ;
    wire signal_17195 ;
    wire signal_17196 ;
    wire signal_17197 ;
    wire signal_17198 ;
    wire signal_17199 ;
    wire signal_17200 ;
    wire signal_17201 ;
    wire signal_17202 ;
    wire signal_17203 ;
    wire signal_17204 ;
    wire signal_17205 ;
    wire signal_17206 ;
    wire signal_17207 ;
    wire signal_17208 ;
    wire signal_17209 ;
    wire signal_17210 ;
    wire signal_17211 ;
    wire signal_17212 ;
    wire signal_17213 ;
    wire signal_17214 ;
    wire signal_17215 ;
    wire signal_17216 ;
    wire signal_17217 ;
    wire signal_17218 ;
    wire signal_17219 ;
    wire signal_17220 ;
    wire signal_17221 ;
    wire signal_17222 ;
    wire signal_17223 ;
    wire signal_17224 ;
    wire signal_17225 ;
    wire signal_17226 ;
    wire signal_17227 ;
    wire signal_17228 ;
    wire signal_17229 ;
    wire signal_17230 ;
    wire signal_17231 ;
    wire signal_17232 ;
    wire signal_17233 ;
    wire signal_17234 ;
    wire signal_17235 ;
    wire signal_17236 ;
    wire signal_17237 ;
    wire signal_17238 ;
    wire signal_17239 ;
    wire signal_17240 ;
    wire signal_17241 ;
    wire signal_17242 ;
    wire signal_17243 ;
    wire signal_17244 ;
    wire signal_17245 ;
    wire signal_17246 ;
    wire signal_17247 ;
    wire signal_17248 ;
    wire signal_17249 ;
    wire signal_17250 ;
    wire signal_17251 ;
    wire signal_17252 ;
    wire signal_17253 ;
    wire signal_17254 ;
    wire signal_17255 ;
    wire signal_17256 ;
    wire signal_17257 ;
    wire signal_17258 ;
    wire signal_17259 ;
    wire signal_17260 ;
    wire signal_17261 ;
    wire signal_17262 ;
    wire signal_17263 ;
    wire signal_17264 ;
    wire signal_17265 ;
    wire signal_17266 ;
    wire signal_17267 ;
    wire signal_17268 ;
    wire signal_17269 ;
    wire signal_17270 ;
    wire signal_17271 ;
    wire signal_17272 ;
    wire signal_17273 ;
    wire signal_17274 ;
    wire signal_17275 ;
    wire signal_17276 ;
    wire signal_17277 ;
    wire signal_17278 ;
    wire signal_17279 ;
    wire signal_17280 ;
    wire signal_17281 ;
    wire signal_17282 ;
    wire signal_17283 ;
    wire signal_17284 ;
    wire signal_17285 ;
    wire signal_17286 ;
    wire signal_17287 ;
    wire signal_17288 ;
    wire signal_17289 ;
    wire signal_17290 ;
    wire signal_17291 ;
    wire signal_17292 ;
    wire signal_17293 ;
    wire signal_17294 ;
    wire signal_17295 ;
    wire signal_17296 ;
    wire signal_17297 ;
    wire signal_17298 ;
    wire signal_17299 ;
    wire signal_17300 ;
    wire signal_17301 ;
    wire signal_17302 ;
    wire signal_17303 ;
    wire signal_17304 ;
    wire signal_17305 ;
    wire signal_17306 ;
    wire signal_17307 ;
    wire signal_17308 ;
    wire signal_17309 ;
    wire signal_17310 ;
    wire signal_17311 ;
    wire signal_17312 ;
    wire signal_17313 ;
    wire signal_17314 ;
    wire signal_17315 ;
    wire signal_17316 ;
    wire signal_17317 ;
    wire signal_17318 ;
    wire signal_17319 ;
    wire signal_17320 ;
    wire signal_17321 ;
    wire signal_17322 ;
    wire signal_17323 ;
    wire signal_17324 ;
    wire signal_17325 ;
    wire signal_17326 ;
    wire signal_17327 ;
    wire signal_17328 ;
    wire signal_17329 ;
    wire signal_17330 ;
    wire signal_17331 ;
    wire signal_17332 ;
    wire signal_17333 ;
    wire signal_17334 ;
    wire signal_17335 ;
    wire signal_17336 ;
    wire signal_17337 ;
    wire signal_17338 ;
    wire signal_17339 ;
    wire signal_17340 ;
    wire signal_17341 ;
    wire signal_17342 ;
    wire signal_17343 ;
    wire signal_17344 ;
    wire signal_17345 ;
    wire signal_17346 ;
    wire signal_17347 ;
    wire signal_17348 ;
    wire signal_17349 ;
    wire signal_17350 ;
    wire signal_17351 ;
    wire signal_17352 ;
    wire signal_17353 ;
    wire signal_17354 ;
    wire signal_17355 ;
    wire signal_17356 ;
    wire signal_17357 ;
    wire signal_17358 ;
    wire signal_17359 ;
    wire signal_17360 ;
    wire signal_17361 ;
    wire signal_17362 ;
    wire signal_17363 ;
    wire signal_17364 ;
    wire signal_17365 ;
    wire signal_17366 ;
    wire signal_17367 ;
    wire signal_17368 ;
    wire signal_17369 ;
    wire signal_17370 ;
    wire signal_17371 ;
    wire signal_17372 ;
    wire signal_17373 ;
    wire signal_17374 ;
    wire signal_17375 ;
    wire signal_17376 ;
    wire signal_17377 ;
    wire signal_17378 ;
    wire signal_17379 ;
    wire signal_17380 ;
    wire signal_17381 ;
    wire signal_17382 ;
    wire signal_17383 ;
    wire signal_17384 ;
    wire signal_17385 ;
    wire signal_17386 ;
    wire signal_17387 ;
    wire signal_17388 ;
    wire signal_17389 ;
    wire signal_17390 ;
    wire signal_17391 ;
    wire signal_17392 ;
    wire signal_17393 ;
    wire signal_17394 ;
    wire signal_17395 ;
    wire signal_17396 ;
    wire signal_17397 ;
    wire signal_17398 ;
    wire signal_17399 ;
    wire signal_17400 ;
    wire signal_17401 ;
    wire signal_17402 ;
    wire signal_17403 ;
    wire signal_17404 ;
    wire signal_17405 ;
    wire signal_17406 ;
    wire signal_17407 ;
    wire signal_17408 ;
    wire signal_17409 ;
    wire signal_17410 ;
    wire signal_17411 ;
    wire signal_17412 ;
    wire signal_17413 ;
    wire signal_17414 ;
    wire signal_17415 ;
    wire signal_17416 ;
    wire signal_17417 ;
    wire signal_17418 ;
    wire signal_17419 ;
    wire signal_17420 ;
    wire signal_17421 ;
    wire signal_17422 ;
    wire signal_17423 ;
    wire signal_17424 ;
    wire signal_17425 ;
    wire signal_17426 ;
    wire signal_17427 ;
    wire signal_17428 ;
    wire signal_17429 ;
    wire signal_17430 ;
    wire signal_17431 ;
    wire signal_17432 ;
    wire signal_17433 ;
    wire signal_17434 ;
    wire signal_17435 ;
    wire signal_17436 ;
    wire signal_17437 ;
    wire signal_17438 ;
    wire signal_17439 ;
    wire signal_17440 ;
    wire signal_17441 ;
    wire signal_17442 ;
    wire signal_17443 ;
    wire signal_17444 ;
    wire signal_17445 ;
    wire signal_17446 ;
    wire signal_17447 ;
    wire signal_17448 ;
    wire signal_17449 ;
    wire signal_17450 ;
    wire signal_17451 ;
    wire signal_17452 ;
    wire signal_17453 ;
    wire signal_17454 ;
    wire signal_17455 ;
    wire signal_17456 ;
    wire signal_17457 ;
    wire signal_17458 ;
    wire signal_17459 ;
    wire signal_17460 ;
    wire signal_17461 ;
    wire signal_17462 ;
    wire signal_17463 ;
    wire signal_17464 ;
    wire signal_17465 ;
    wire signal_17466 ;
    wire signal_17467 ;
    wire signal_17468 ;
    wire signal_17469 ;
    wire signal_17470 ;
    wire signal_17471 ;
    wire signal_17472 ;
    wire signal_17473 ;
    wire signal_17474 ;
    wire signal_17475 ;
    wire signal_17476 ;
    wire signal_17477 ;
    wire signal_17478 ;
    wire signal_17479 ;
    wire signal_17480 ;
    wire signal_17481 ;
    wire signal_17482 ;
    wire signal_17483 ;
    wire signal_17484 ;
    wire signal_17485 ;
    wire signal_17486 ;
    wire signal_17487 ;
    wire signal_17488 ;
    wire signal_17489 ;
    wire signal_17490 ;
    wire signal_17491 ;
    wire signal_17492 ;
    wire signal_17493 ;
    wire signal_17494 ;
    wire signal_17495 ;
    wire signal_17496 ;
    wire signal_17497 ;
    wire signal_17498 ;
    wire signal_17499 ;
    wire signal_17500 ;
    wire signal_17501 ;
    wire signal_17502 ;
    wire signal_17503 ;
    wire signal_17504 ;
    wire signal_17505 ;
    wire signal_17506 ;
    wire signal_17507 ;
    wire signal_17508 ;
    wire signal_17509 ;
    wire signal_17510 ;
    wire signal_17511 ;
    wire signal_17512 ;
    wire signal_17513 ;
    wire signal_17514 ;
    wire signal_17515 ;
    wire signal_17516 ;
    wire signal_17517 ;
    wire signal_17518 ;
    wire signal_17519 ;
    wire signal_17520 ;
    wire signal_17521 ;
    wire signal_17522 ;
    wire signal_17523 ;
    wire signal_17524 ;
    wire signal_17525 ;
    wire signal_17526 ;
    wire signal_17527 ;
    wire signal_17528 ;
    wire signal_17529 ;
    wire signal_17530 ;
    wire signal_17531 ;
    wire signal_17532 ;
    wire signal_17533 ;
    wire signal_17534 ;
    wire signal_17535 ;
    wire signal_17536 ;
    wire signal_17537 ;
    wire signal_17538 ;
    wire signal_17539 ;
    wire signal_17540 ;
    wire signal_17541 ;
    wire signal_17542 ;
    wire signal_17543 ;
    wire signal_17544 ;
    wire signal_17545 ;
    wire signal_17546 ;
    wire signal_17547 ;
    wire signal_17548 ;
    wire signal_17549 ;
    wire signal_17550 ;
    wire signal_17551 ;
    wire signal_17552 ;
    wire signal_17553 ;
    wire signal_17554 ;
    wire signal_17555 ;
    wire signal_17556 ;
    wire signal_17557 ;
    wire signal_17558 ;
    wire signal_17559 ;
    wire signal_17560 ;
    wire signal_17561 ;
    wire signal_17562 ;
    wire signal_17563 ;
    wire signal_17564 ;
    wire signal_17565 ;
    wire signal_17566 ;
    wire signal_17567 ;
    wire signal_17568 ;
    wire signal_17569 ;
    wire signal_17570 ;
    wire signal_17571 ;
    wire signal_17572 ;
    wire signal_17573 ;
    wire signal_17574 ;
    wire signal_17575 ;
    wire signal_17576 ;
    wire signal_17577 ;
    wire signal_17578 ;
    wire signal_17579 ;
    wire signal_17580 ;
    wire signal_17581 ;
    wire signal_17582 ;
    wire signal_17583 ;
    wire signal_17584 ;
    wire signal_17585 ;
    wire signal_17586 ;
    wire signal_17587 ;
    wire signal_17588 ;
    wire signal_17589 ;
    wire signal_17590 ;
    wire signal_17591 ;
    wire signal_17592 ;
    wire signal_17593 ;
    wire signal_17594 ;
    wire signal_17595 ;
    wire signal_17596 ;
    wire signal_17597 ;
    wire signal_17598 ;
    wire signal_17599 ;
    wire signal_17600 ;
    wire signal_17601 ;
    wire signal_17602 ;
    wire signal_17603 ;
    wire signal_17604 ;
    wire signal_17605 ;
    wire signal_17606 ;
    wire signal_17607 ;
    wire signal_17608 ;
    wire signal_17609 ;
    wire signal_17610 ;
    wire signal_17611 ;
    wire signal_17612 ;
    wire signal_17613 ;
    wire signal_17614 ;
    wire signal_17615 ;
    wire signal_17616 ;
    wire signal_17617 ;
    wire signal_17618 ;
    wire signal_17619 ;
    wire signal_17620 ;
    wire signal_17621 ;
    wire signal_17622 ;
    wire signal_17623 ;
    wire signal_17624 ;
    wire signal_17625 ;
    wire signal_17626 ;
    wire signal_17627 ;
    wire signal_17628 ;
    wire signal_17629 ;
    wire signal_17630 ;
    wire signal_17631 ;
    wire signal_17632 ;
    wire signal_17633 ;
    wire signal_17634 ;
    wire signal_17635 ;
    wire signal_17636 ;
    wire signal_17637 ;
    wire signal_17638 ;
    wire signal_17639 ;
    wire signal_17640 ;
    wire signal_17641 ;
    wire signal_17642 ;
    wire signal_17643 ;
    wire signal_17644 ;
    wire signal_17645 ;
    wire signal_17646 ;
    wire signal_17647 ;
    wire signal_17648 ;
    wire signal_17649 ;
    wire signal_17650 ;
    wire signal_17651 ;
    wire signal_17652 ;
    wire signal_17653 ;
    wire signal_17654 ;
    wire signal_17655 ;
    wire signal_17656 ;
    wire signal_17657 ;
    wire signal_17658 ;
    wire signal_17659 ;
    wire signal_17660 ;
    wire signal_17661 ;
    wire signal_17662 ;
    wire signal_17663 ;
    wire signal_17664 ;
    wire signal_17665 ;
    wire signal_17666 ;
    wire signal_17667 ;
    wire signal_17668 ;
    wire signal_17669 ;
    wire signal_17670 ;
    wire signal_17671 ;
    wire signal_17672 ;
    wire signal_17673 ;
    wire signal_17674 ;
    wire signal_17675 ;
    wire signal_17676 ;
    wire signal_17677 ;
    wire signal_17678 ;
    wire signal_17679 ;
    wire signal_17680 ;
    wire signal_17681 ;
    wire signal_17682 ;
    wire signal_17683 ;
    wire signal_17684 ;
    wire signal_17685 ;
    wire signal_17686 ;
    wire signal_17687 ;
    wire signal_17688 ;
    wire signal_17689 ;
    wire signal_17690 ;
    wire signal_17691 ;
    wire signal_17692 ;
    wire signal_17693 ;
    wire signal_17694 ;
    wire signal_17695 ;
    wire signal_17696 ;
    wire signal_17697 ;
    wire signal_17698 ;
    wire signal_17699 ;
    wire signal_17700 ;
    wire signal_17701 ;
    wire signal_17702 ;
    wire signal_17703 ;
    wire signal_17704 ;
    wire signal_17705 ;
    wire signal_17706 ;
    wire signal_17707 ;
    wire signal_17708 ;
    wire signal_17709 ;
    wire signal_17710 ;
    wire signal_17711 ;
    wire signal_17712 ;
    wire signal_17713 ;
    wire signal_17714 ;
    wire signal_17715 ;
    wire signal_17716 ;
    wire signal_17717 ;
    wire signal_17718 ;
    wire signal_17719 ;
    wire signal_17720 ;
    wire signal_17721 ;
    wire signal_17722 ;
    wire signal_17723 ;
    wire signal_17724 ;
    wire signal_17725 ;
    wire signal_17726 ;
    wire signal_17727 ;
    wire signal_17728 ;
    wire signal_17729 ;
    wire signal_17730 ;
    wire signal_17731 ;
    wire signal_17732 ;
    wire signal_17733 ;
    wire signal_17734 ;
    wire signal_17735 ;
    wire signal_17736 ;
    wire signal_17737 ;
    wire signal_17738 ;
    wire signal_17739 ;
    wire signal_17740 ;
    wire signal_17741 ;
    wire signal_17742 ;
    wire signal_17743 ;
    wire signal_17744 ;
    wire signal_17745 ;
    wire signal_17746 ;
    wire signal_17747 ;
    wire signal_17748 ;
    wire signal_17749 ;
    wire signal_17750 ;
    wire signal_17751 ;
    wire signal_17752 ;
    wire signal_17753 ;
    wire signal_17754 ;
    wire signal_17755 ;
    wire signal_17756 ;
    wire signal_17757 ;
    wire signal_17758 ;
    wire signal_17759 ;
    wire signal_17760 ;
    wire signal_17761 ;
    wire signal_17762 ;
    wire signal_17763 ;
    wire signal_17764 ;
    wire signal_17765 ;
    wire signal_17766 ;
    wire signal_17767 ;
    wire signal_17768 ;
    wire signal_17769 ;
    wire signal_17770 ;
    wire signal_17771 ;
    wire signal_17772 ;
    wire signal_17773 ;
    wire signal_17774 ;
    wire signal_17775 ;
    wire signal_17776 ;
    wire signal_17777 ;
    wire signal_17778 ;
    wire signal_17779 ;
    wire signal_17780 ;
    wire signal_17781 ;
    wire signal_17782 ;
    wire signal_17783 ;
    wire signal_17784 ;
    wire signal_17785 ;
    wire signal_17786 ;
    wire signal_17787 ;
    wire signal_17788 ;
    wire signal_17789 ;
    wire signal_17790 ;
    wire signal_17791 ;
    wire signal_17792 ;
    wire signal_17793 ;
    wire signal_17794 ;
    wire signal_17795 ;
    wire signal_17796 ;
    wire signal_17797 ;
    wire signal_17798 ;
    wire signal_17799 ;
    wire signal_17800 ;
    wire signal_17801 ;
    wire signal_17802 ;
    wire signal_17803 ;
    wire signal_17804 ;
    wire signal_17805 ;
    wire signal_17806 ;
    wire signal_17807 ;
    wire signal_17808 ;
    wire signal_17809 ;
    wire signal_17810 ;
    wire signal_17811 ;
    wire signal_17812 ;
    wire signal_17813 ;
    wire signal_17814 ;
    wire signal_17815 ;
    wire signal_17816 ;
    wire signal_17817 ;
    wire signal_17818 ;
    wire signal_17819 ;
    wire signal_17820 ;
    wire signal_17821 ;
    wire signal_17822 ;
    wire signal_17823 ;
    wire signal_17824 ;
    wire signal_17825 ;
    wire signal_17826 ;
    wire signal_17827 ;
    wire signal_17828 ;
    wire signal_17829 ;
    wire signal_17830 ;
    wire signal_17831 ;
    wire signal_17832 ;
    wire signal_17833 ;
    wire signal_17834 ;
    wire signal_17835 ;
    wire signal_17836 ;
    wire signal_17837 ;
    wire signal_17838 ;
    wire signal_17839 ;
    wire signal_17840 ;
    wire signal_17841 ;
    wire signal_17842 ;
    wire signal_17843 ;
    wire signal_17844 ;
    wire signal_17845 ;
    wire signal_17846 ;
    wire signal_17847 ;
    wire signal_17848 ;
    wire signal_17849 ;
    wire signal_17850 ;
    wire signal_17851 ;
    wire signal_17852 ;
    wire signal_17853 ;
    wire signal_17854 ;
    wire signal_17855 ;
    wire signal_17856 ;
    wire signal_17857 ;
    wire signal_17858 ;
    wire signal_17859 ;
    wire signal_17860 ;
    wire signal_17861 ;
    wire signal_17862 ;
    wire signal_17863 ;
    wire signal_17864 ;
    wire signal_17865 ;
    wire signal_17866 ;
    wire signal_17867 ;
    wire signal_17868 ;
    wire signal_17869 ;
    wire signal_17870 ;
    wire signal_17871 ;
    wire signal_17872 ;
    wire signal_17873 ;
    wire signal_17874 ;
    wire signal_17875 ;
    wire signal_17876 ;
    wire signal_17877 ;
    wire signal_17878 ;
    wire signal_17879 ;
    wire signal_17880 ;
    wire signal_17881 ;
    wire signal_17882 ;
    wire signal_17883 ;
    wire signal_17884 ;
    wire signal_17885 ;
    wire signal_17886 ;
    wire signal_17887 ;
    wire signal_17888 ;
    wire signal_17889 ;
    wire signal_17890 ;
    wire signal_17891 ;
    wire signal_17892 ;
    wire signal_17893 ;
    wire signal_17894 ;
    wire signal_17895 ;
    wire signal_17896 ;
    wire signal_17897 ;
    wire signal_17898 ;
    wire signal_17899 ;
    wire signal_17900 ;
    wire signal_17901 ;
    wire signal_17902 ;
    wire signal_17903 ;
    wire signal_17904 ;
    wire signal_17905 ;
    wire signal_17906 ;
    wire signal_17907 ;
    wire signal_17908 ;
    wire signal_17909 ;
    wire signal_17910 ;
    wire signal_17911 ;
    wire signal_17912 ;
    wire signal_17913 ;
    wire signal_17914 ;
    wire signal_17915 ;
    wire signal_17916 ;
    wire signal_17917 ;
    wire signal_17918 ;
    wire signal_17919 ;
    wire signal_17920 ;
    wire signal_17921 ;
    wire signal_17922 ;
    wire signal_17923 ;
    wire signal_17924 ;
    wire signal_17925 ;
    wire signal_17926 ;
    wire signal_17927 ;
    wire signal_17928 ;
    wire signal_17929 ;
    wire signal_17930 ;
    wire signal_17931 ;
    wire signal_17932 ;
    wire signal_17933 ;
    wire signal_17934 ;
    wire signal_17935 ;
    wire signal_17936 ;
    wire signal_17937 ;
    wire signal_17938 ;
    wire signal_17939 ;
    wire signal_17940 ;
    wire signal_17941 ;
    wire signal_17942 ;
    wire signal_17943 ;
    wire signal_17944 ;
    wire signal_17945 ;
    wire signal_17946 ;
    wire signal_17947 ;
    wire signal_17948 ;
    wire signal_17949 ;
    wire signal_17950 ;
    wire signal_17951 ;
    wire signal_17952 ;
    wire signal_17953 ;
    wire signal_17954 ;
    wire signal_17955 ;
    wire signal_17956 ;
    wire signal_17957 ;
    wire signal_17958 ;
    wire signal_17959 ;
    wire signal_17960 ;
    wire signal_17961 ;
    wire signal_17962 ;
    wire signal_17963 ;
    wire signal_17964 ;
    wire signal_17965 ;
    wire signal_17966 ;
    wire signal_17967 ;
    wire signal_17968 ;
    wire signal_17969 ;
    wire signal_17970 ;
    wire signal_17971 ;
    wire signal_17972 ;
    wire signal_17973 ;
    wire signal_17974 ;
    wire signal_17975 ;
    wire signal_17976 ;
    wire signal_17977 ;
    wire signal_17978 ;
    wire signal_17979 ;
    wire signal_17980 ;
    wire signal_17981 ;
    wire signal_17982 ;
    wire signal_17983 ;
    wire signal_17984 ;
    wire signal_17985 ;
    wire signal_17986 ;
    wire signal_17987 ;
    wire signal_17988 ;
    wire signal_17989 ;
    wire signal_17990 ;
    wire signal_17991 ;
    wire signal_17992 ;
    wire signal_17993 ;
    wire signal_17994 ;
    wire signal_17995 ;
    wire signal_17996 ;
    wire signal_17997 ;
    wire signal_17998 ;
    wire signal_17999 ;
    wire signal_18000 ;
    wire signal_18001 ;
    wire signal_18002 ;
    wire signal_18003 ;
    wire signal_18004 ;
    wire signal_18005 ;
    wire signal_18006 ;
    wire signal_18007 ;
    wire signal_18008 ;
    wire signal_18009 ;
    wire signal_18010 ;
    wire signal_18011 ;
    wire signal_18012 ;
    wire signal_18013 ;
    wire signal_18014 ;
    wire signal_18015 ;
    wire signal_18016 ;
    wire signal_18017 ;
    wire signal_18018 ;
    wire signal_18019 ;
    wire signal_18020 ;
    wire signal_18021 ;
    wire signal_18022 ;
    wire signal_18023 ;
    wire signal_18024 ;
    wire signal_18025 ;
    wire signal_18026 ;
    wire signal_18027 ;
    wire signal_18028 ;
    wire signal_18029 ;
    wire signal_18030 ;
    wire signal_18031 ;
    wire signal_18032 ;
    wire signal_18033 ;
    wire signal_18034 ;
    wire signal_18035 ;
    wire signal_18036 ;
    wire signal_18037 ;
    wire signal_18038 ;
    wire signal_18039 ;
    wire signal_18040 ;
    wire signal_18041 ;
    wire signal_18042 ;
    wire signal_18043 ;
    wire signal_18044 ;
    wire signal_18045 ;
    wire signal_18046 ;
    wire signal_18047 ;
    wire signal_18048 ;
    wire signal_18049 ;
    wire signal_18050 ;
    wire signal_18051 ;
    wire signal_18052 ;
    wire signal_18053 ;
    wire signal_18054 ;
    wire signal_18055 ;
    wire signal_18056 ;
    wire signal_18057 ;
    wire signal_18058 ;
    wire signal_18059 ;
    wire signal_18060 ;
    wire signal_18061 ;
    wire signal_18062 ;
    wire signal_18063 ;
    wire signal_18064 ;
    wire signal_18065 ;
    wire signal_18066 ;
    wire signal_18067 ;
    wire signal_18068 ;
    wire signal_18069 ;
    wire signal_18070 ;
    wire signal_18071 ;
    wire signal_18072 ;
    wire signal_18073 ;
    wire signal_18074 ;
    wire signal_18075 ;
    wire signal_18076 ;
    wire signal_18077 ;
    wire signal_18078 ;
    wire signal_18079 ;
    wire signal_18080 ;
    wire signal_18081 ;
    wire signal_18082 ;
    wire signal_18083 ;
    wire signal_18084 ;
    wire signal_18085 ;
    wire signal_18086 ;
    wire signal_18087 ;
    wire signal_18088 ;
    wire signal_18089 ;
    wire signal_18090 ;
    wire signal_18091 ;
    wire signal_18092 ;
    wire signal_18093 ;
    wire signal_18094 ;
    wire signal_18095 ;
    wire signal_18096 ;
    wire signal_18097 ;
    wire signal_18098 ;
    wire signal_18099 ;
    wire signal_18100 ;
    wire signal_18101 ;
    wire signal_18102 ;
    wire signal_18103 ;
    wire signal_18104 ;
    wire signal_18105 ;
    wire signal_18106 ;
    wire signal_18107 ;
    wire signal_18108 ;
    wire signal_18109 ;
    wire signal_18110 ;
    wire signal_18111 ;
    wire signal_18112 ;
    wire signal_18113 ;
    wire signal_18114 ;
    wire signal_18115 ;
    wire signal_18116 ;
    wire signal_18117 ;
    wire signal_18118 ;
    wire signal_18119 ;
    wire signal_18120 ;
    wire signal_18121 ;
    wire signal_18122 ;
    wire signal_18123 ;
    wire signal_18124 ;
    wire signal_18125 ;
    wire signal_18126 ;
    wire signal_18127 ;
    wire signal_18128 ;
    wire signal_18129 ;
    wire signal_18130 ;
    wire signal_18131 ;
    wire signal_18132 ;
    wire signal_18133 ;
    wire signal_18134 ;
    wire signal_18135 ;
    wire signal_18136 ;
    wire signal_18137 ;
    wire signal_18138 ;
    wire signal_18139 ;
    wire signal_18140 ;
    wire signal_18141 ;
    wire signal_18142 ;
    wire signal_18143 ;
    wire signal_18144 ;
    wire signal_18145 ;
    wire signal_18146 ;
    wire signal_18147 ;
    wire signal_18148 ;
    wire signal_18149 ;
    wire signal_18150 ;
    wire signal_18151 ;
    wire signal_18152 ;
    wire signal_18153 ;
    wire signal_18154 ;
    wire signal_18155 ;
    wire signal_18156 ;
    wire signal_18157 ;
    wire signal_18158 ;
    wire signal_18159 ;
    wire signal_18160 ;
    wire signal_18161 ;
    wire signal_18162 ;
    wire signal_18163 ;
    wire signal_18164 ;
    wire signal_18165 ;
    wire signal_18166 ;
    wire signal_18167 ;
    wire signal_18168 ;
    wire signal_18169 ;
    wire signal_18170 ;
    wire signal_18171 ;
    wire signal_18172 ;
    wire signal_18173 ;
    wire signal_18174 ;
    wire signal_18175 ;
    wire signal_18176 ;
    wire signal_18177 ;
    wire signal_18178 ;
    wire signal_18179 ;
    wire signal_18180 ;
    wire signal_18181 ;
    wire signal_18182 ;
    wire signal_18183 ;
    wire signal_18184 ;
    wire signal_18185 ;
    wire signal_18186 ;
    wire signal_18187 ;
    wire signal_18188 ;
    wire signal_18189 ;
    wire signal_18190 ;
    wire signal_18191 ;
    wire signal_18192 ;
    wire signal_18193 ;
    wire signal_18194 ;
    wire signal_18195 ;
    wire signal_18196 ;
    wire signal_18197 ;
    wire signal_18198 ;
    wire signal_18199 ;
    wire signal_18200 ;
    wire signal_18201 ;
    wire signal_18202 ;
    wire signal_18203 ;
    wire signal_18204 ;
    wire signal_18205 ;
    wire signal_18206 ;
    wire signal_18207 ;
    wire signal_18208 ;
    wire signal_18209 ;
    wire signal_18210 ;
    wire signal_18211 ;
    wire signal_18212 ;
    wire signal_18213 ;
    wire signal_18214 ;
    wire signal_18215 ;
    wire signal_18216 ;
    wire signal_18217 ;
    wire signal_18218 ;
    wire signal_18219 ;
    wire signal_18220 ;
    wire signal_18221 ;
    wire signal_18222 ;
    wire signal_18223 ;
    wire signal_18224 ;
    wire signal_18225 ;
    wire signal_18226 ;
    wire signal_18227 ;
    wire signal_18228 ;
    wire signal_18229 ;
    wire signal_18230 ;
    wire signal_18231 ;
    wire signal_18232 ;
    wire signal_18233 ;
    wire signal_18234 ;
    wire signal_18235 ;
    wire signal_18236 ;
    wire signal_18237 ;
    wire signal_18238 ;
    wire signal_18239 ;
    wire signal_18240 ;
    wire signal_18241 ;
    wire signal_18242 ;
    wire signal_18243 ;
    wire signal_18244 ;
    wire signal_18245 ;
    wire signal_18246 ;
    wire signal_18247 ;
    wire signal_18248 ;
    wire signal_18249 ;
    wire signal_18250 ;
    wire signal_18251 ;
    wire signal_18252 ;
    wire signal_18253 ;
    wire signal_18254 ;
    wire signal_18255 ;
    wire signal_18256 ;
    wire signal_18257 ;
    wire signal_18258 ;
    wire signal_18259 ;
    wire signal_18260 ;
    wire signal_18261 ;
    wire signal_18262 ;
    wire signal_18263 ;
    wire signal_18264 ;
    wire signal_18265 ;
    wire signal_18266 ;
    wire signal_18267 ;
    wire signal_18268 ;
    wire signal_18269 ;
    wire signal_18270 ;
    wire signal_18271 ;
    wire signal_18272 ;
    wire signal_18273 ;
    wire signal_18274 ;
    wire signal_18275 ;
    wire signal_18276 ;
    wire signal_18277 ;
    wire signal_18278 ;
    wire signal_18279 ;
    wire signal_18280 ;
    wire signal_18281 ;
    wire signal_18282 ;
    wire signal_18283 ;
    wire signal_18284 ;
    wire signal_18285 ;
    wire signal_18286 ;
    wire signal_18287 ;
    wire signal_18288 ;
    wire signal_18289 ;
    wire signal_18290 ;
    wire signal_18291 ;
    wire signal_18292 ;
    wire signal_18293 ;
    wire signal_18294 ;
    wire signal_18295 ;
    wire signal_18296 ;
    wire signal_18297 ;
    wire signal_18298 ;
    wire signal_18299 ;
    wire signal_18300 ;
    wire signal_18301 ;
    wire signal_18302 ;
    wire signal_18303 ;
    wire signal_18304 ;
    wire signal_18305 ;
    wire signal_18306 ;
    wire signal_18307 ;
    wire signal_18308 ;
    wire signal_18309 ;
    wire signal_18310 ;
    wire signal_18311 ;
    wire signal_18312 ;
    wire signal_18313 ;
    wire signal_18314 ;
    wire signal_18315 ;
    wire signal_18316 ;
    wire signal_18317 ;
    wire signal_18318 ;
    wire signal_18319 ;
    wire signal_18320 ;
    wire signal_18321 ;
    wire signal_18322 ;
    wire signal_18323 ;
    wire signal_18324 ;
    wire signal_18325 ;
    wire signal_18326 ;
    wire signal_18327 ;
    wire signal_18328 ;
    wire signal_18329 ;
    wire signal_18330 ;
    wire signal_18331 ;
    wire signal_18332 ;
    wire signal_18333 ;
    wire signal_18334 ;
    wire signal_18335 ;
    wire signal_18336 ;
    wire signal_18337 ;
    wire signal_18338 ;
    wire signal_18339 ;
    wire signal_18340 ;
    wire signal_18341 ;
    wire signal_18342 ;
    wire signal_18343 ;
    wire signal_18344 ;
    wire signal_18345 ;
    wire signal_18346 ;
    wire signal_18347 ;
    wire signal_18348 ;
    wire signal_18349 ;
    wire signal_18350 ;
    wire signal_18351 ;
    wire signal_18352 ;
    wire signal_18353 ;
    wire signal_18354 ;
    wire signal_18355 ;
    wire signal_18356 ;
    wire signal_18357 ;
    wire signal_18358 ;
    wire signal_18359 ;
    wire signal_18360 ;
    wire signal_18361 ;
    wire signal_18362 ;
    wire signal_18363 ;
    wire signal_18364 ;
    wire signal_18365 ;
    wire signal_18366 ;
    wire signal_18367 ;
    wire signal_18368 ;
    wire signal_18369 ;
    wire signal_18370 ;
    wire signal_18371 ;
    wire signal_18372 ;
    wire signal_18373 ;
    wire signal_18374 ;
    wire signal_18375 ;
    wire signal_18376 ;
    wire signal_18377 ;
    wire signal_18378 ;
    wire signal_18379 ;
    wire signal_18380 ;
    wire signal_18381 ;
    wire signal_18382 ;
    wire signal_18383 ;
    wire signal_18384 ;
    wire signal_18385 ;
    wire signal_18386 ;
    wire signal_18387 ;
    wire signal_18388 ;
    wire signal_18389 ;
    wire signal_18390 ;
    wire signal_18391 ;
    wire signal_18392 ;
    wire signal_18393 ;
    wire signal_18394 ;
    wire signal_18395 ;
    wire signal_18396 ;
    wire signal_18397 ;
    wire signal_18398 ;
    wire signal_18399 ;
    wire signal_18400 ;
    wire signal_18401 ;
    wire signal_18402 ;
    wire signal_18403 ;
    wire signal_18404 ;
    wire signal_18405 ;
    wire signal_18406 ;
    wire signal_18407 ;
    wire signal_18408 ;
    wire signal_18409 ;
    wire signal_18410 ;
    wire signal_18411 ;
    wire signal_18412 ;
    wire signal_18413 ;
    wire signal_18414 ;
    wire signal_18415 ;
    wire signal_18416 ;
    wire signal_18417 ;
    wire signal_18418 ;
    wire signal_18419 ;
    wire signal_18420 ;
    wire signal_18421 ;
    wire signal_18422 ;
    wire signal_18423 ;
    wire signal_18424 ;
    wire signal_18425 ;
    wire signal_18426 ;
    wire signal_18427 ;
    wire signal_18428 ;
    wire signal_18429 ;
    wire signal_18430 ;
    wire signal_18431 ;
    wire signal_18432 ;
    wire signal_18433 ;
    wire signal_18434 ;
    wire signal_18435 ;
    wire signal_18436 ;
    wire signal_18437 ;
    wire signal_18438 ;
    wire signal_18439 ;
    wire signal_18440 ;
    wire signal_18441 ;
    wire signal_18442 ;
    wire signal_18443 ;
    wire signal_18444 ;
    wire signal_18445 ;
    wire signal_18446 ;
    wire signal_18447 ;
    wire signal_18448 ;
    wire signal_18449 ;
    wire signal_18450 ;
    wire signal_18451 ;
    wire signal_18452 ;
    wire signal_18453 ;
    wire signal_18454 ;
    wire signal_18455 ;
    wire signal_18456 ;
    wire signal_18457 ;
    wire signal_18458 ;
    wire signal_18459 ;
    wire signal_18460 ;
    wire signal_18461 ;
    wire signal_18462 ;
    wire signal_18463 ;
    wire signal_18464 ;
    wire signal_18465 ;
    wire signal_18466 ;
    wire signal_18467 ;
    wire signal_18468 ;
    wire signal_18469 ;
    wire signal_18470 ;
    wire signal_18471 ;
    wire signal_18472 ;
    wire signal_18473 ;
    wire signal_18474 ;
    wire signal_18475 ;
    wire signal_18476 ;
    wire signal_18477 ;
    wire signal_18478 ;
    wire signal_18479 ;
    wire signal_18480 ;
    wire signal_18481 ;
    wire signal_18482 ;
    wire signal_18483 ;
    wire signal_18484 ;
    wire signal_18485 ;
    wire signal_18486 ;
    wire signal_18487 ;
    wire signal_18488 ;
    wire signal_18489 ;
    wire signal_18490 ;
    wire signal_18491 ;
    wire signal_18492 ;
    wire signal_18493 ;
    wire signal_18494 ;
    wire signal_18495 ;
    wire signal_18496 ;
    wire signal_18497 ;
    wire signal_18498 ;
    wire signal_18499 ;
    wire signal_18500 ;
    wire signal_18501 ;
    wire signal_18502 ;
    wire signal_18503 ;
    wire signal_18504 ;
    wire signal_18505 ;
    wire signal_18506 ;
    wire signal_18507 ;
    wire signal_18508 ;
    wire signal_18509 ;
    wire signal_18510 ;
    wire signal_18511 ;
    wire signal_18512 ;
    wire signal_18513 ;
    wire signal_18514 ;
    wire signal_18515 ;
    wire signal_18516 ;
    wire signal_18517 ;
    wire signal_18518 ;
    wire signal_18519 ;
    wire signal_18520 ;
    wire signal_18521 ;
    wire signal_18522 ;
    wire signal_18523 ;
    wire signal_18524 ;
    wire signal_18525 ;
    wire signal_18526 ;
    wire signal_18527 ;
    wire signal_18528 ;
    wire signal_18529 ;
    wire signal_18530 ;
    wire signal_18531 ;
    wire signal_18532 ;
    wire signal_18533 ;
    wire signal_18534 ;
    wire signal_18535 ;
    wire signal_18536 ;
    wire signal_18537 ;
    wire signal_18538 ;
    wire signal_18539 ;
    wire signal_18540 ;
    wire signal_18541 ;
    wire signal_18542 ;
    wire signal_18543 ;
    wire signal_18544 ;
    wire signal_18545 ;
    wire signal_18546 ;
    wire signal_18547 ;
    wire signal_18548 ;
    wire signal_18549 ;
    wire signal_18550 ;
    wire signal_18551 ;
    wire signal_18552 ;
    wire signal_18553 ;
    wire signal_18554 ;
    wire signal_18555 ;
    wire signal_18556 ;
    wire signal_18557 ;
    wire signal_18558 ;
    wire signal_18559 ;
    wire signal_18560 ;
    wire signal_18561 ;
    wire signal_18562 ;
    wire signal_18563 ;
    wire signal_18564 ;
    wire signal_18565 ;
    wire signal_18566 ;
    wire signal_18567 ;
    wire signal_18568 ;
    wire signal_18569 ;
    wire signal_18570 ;
    wire signal_18571 ;
    wire signal_18572 ;
    wire signal_18573 ;
    wire signal_18574 ;
    wire signal_18575 ;
    wire signal_18576 ;
    wire signal_18577 ;
    wire signal_18578 ;
    wire signal_18579 ;
    wire signal_18580 ;
    wire signal_18581 ;
    wire signal_18582 ;
    wire signal_18583 ;
    wire signal_18584 ;
    wire signal_18585 ;
    wire signal_18586 ;
    wire signal_18587 ;
    wire signal_18588 ;
    wire signal_18589 ;
    wire signal_18590 ;
    wire signal_18591 ;
    wire signal_18592 ;
    wire signal_18593 ;
    wire signal_18594 ;
    wire signal_18595 ;
    wire signal_18596 ;
    wire signal_18597 ;
    wire signal_18598 ;
    wire signal_18599 ;
    wire signal_18600 ;
    wire signal_18601 ;
    wire signal_18602 ;
    wire signal_18603 ;
    wire signal_18604 ;
    wire signal_18605 ;
    wire signal_18606 ;
    wire signal_18607 ;
    wire signal_18608 ;
    wire signal_18609 ;
    wire signal_18610 ;
    wire signal_18611 ;
    wire signal_18612 ;
    wire signal_18613 ;
    wire signal_18614 ;
    wire signal_18615 ;
    wire signal_18616 ;
    wire signal_18617 ;
    wire signal_18618 ;
    wire signal_18619 ;
    wire signal_18620 ;
    wire signal_18621 ;
    wire signal_18622 ;
    wire signal_18623 ;
    wire signal_18624 ;
    wire signal_18625 ;
    wire signal_18626 ;
    wire signal_18627 ;
    wire signal_18628 ;
    wire signal_18629 ;
    wire signal_18630 ;
    wire signal_18631 ;
    wire signal_18632 ;
    wire signal_18633 ;
    wire signal_18634 ;
    wire signal_18635 ;
    wire signal_18636 ;
    wire signal_18637 ;
    wire signal_18638 ;
    wire signal_18639 ;
    wire signal_18640 ;
    wire signal_18641 ;
    wire signal_18642 ;
    wire signal_18643 ;
    wire signal_18644 ;
    wire signal_18645 ;
    wire signal_18646 ;
    wire signal_18647 ;
    wire signal_18648 ;
    wire signal_18649 ;
    wire signal_18650 ;
    wire signal_18651 ;
    wire signal_18652 ;
    wire signal_18653 ;
    wire signal_18654 ;
    wire signal_18655 ;
    wire signal_18656 ;
    wire signal_18657 ;
    wire signal_18658 ;
    wire signal_18659 ;
    wire signal_18660 ;
    wire signal_18661 ;
    wire signal_18662 ;
    wire signal_18663 ;
    wire signal_18664 ;
    wire signal_18665 ;
    wire signal_18666 ;
    wire signal_18667 ;
    wire signal_18668 ;
    wire signal_18669 ;
    wire signal_18670 ;
    wire signal_18671 ;
    wire signal_18672 ;
    wire signal_18673 ;
    wire signal_18674 ;
    wire signal_18675 ;
    wire signal_18676 ;
    wire signal_18677 ;
    wire signal_18678 ;
    wire signal_18679 ;
    wire signal_18680 ;
    wire signal_18681 ;
    wire signal_18682 ;
    wire signal_18683 ;
    wire signal_18684 ;
    wire signal_18685 ;
    wire signal_18686 ;
    wire signal_18687 ;
    wire signal_18688 ;
    wire signal_18689 ;
    wire signal_18690 ;
    wire signal_18691 ;
    wire signal_18692 ;
    wire signal_18693 ;
    wire signal_18694 ;
    wire signal_18695 ;
    wire signal_18696 ;
    wire signal_18697 ;
    wire signal_18698 ;
    wire signal_18699 ;
    wire signal_18700 ;
    wire signal_18701 ;
    wire signal_18702 ;
    wire signal_18703 ;
    wire signal_18704 ;
    wire signal_18705 ;
    wire signal_18706 ;
    wire signal_18707 ;
    wire signal_18708 ;
    wire signal_18709 ;
    wire signal_18710 ;
    wire signal_18711 ;
    wire signal_18712 ;
    wire signal_18713 ;
    wire signal_18714 ;
    wire signal_18715 ;
    wire signal_18716 ;
    wire signal_18717 ;
    wire signal_18718 ;
    wire signal_18719 ;
    wire signal_18720 ;
    wire signal_18721 ;
    wire signal_18722 ;
    wire signal_18723 ;
    wire signal_18724 ;
    wire signal_18725 ;
    wire signal_18726 ;
    wire signal_18727 ;
    wire signal_18728 ;
    wire signal_18729 ;
    wire signal_18730 ;
    wire signal_18731 ;
    wire signal_18732 ;
    wire signal_18733 ;
    wire signal_18734 ;
    wire signal_18735 ;
    wire signal_18736 ;
    wire signal_18737 ;
    wire signal_18738 ;
    wire signal_18739 ;
    wire signal_18740 ;
    wire signal_18741 ;
    wire signal_18742 ;
    wire signal_18743 ;
    wire signal_18744 ;
    wire signal_18745 ;
    wire signal_18746 ;
    wire signal_18747 ;
    wire signal_18748 ;
    wire signal_18749 ;
    wire signal_18750 ;
    wire signal_18751 ;
    wire signal_18752 ;
    wire signal_18753 ;
    wire signal_18754 ;
    wire signal_18755 ;
    wire signal_18756 ;
    wire signal_18757 ;
    wire signal_18758 ;
    wire signal_18759 ;
    wire signal_18760 ;
    wire signal_18761 ;
    wire signal_18762 ;
    wire signal_18763 ;
    wire signal_18764 ;
    wire signal_18765 ;
    wire signal_18766 ;
    wire signal_18767 ;
    wire signal_18768 ;
    wire signal_18769 ;
    wire signal_18770 ;
    wire signal_18771 ;
    wire signal_18772 ;
    wire signal_18773 ;
    wire signal_18774 ;
    wire signal_18775 ;
    wire signal_18776 ;
    wire signal_18777 ;
    wire signal_18778 ;
    wire signal_18779 ;
    wire signal_18780 ;
    wire signal_18781 ;
    wire signal_18782 ;
    wire signal_18783 ;
    wire signal_18784 ;
    wire signal_18785 ;
    wire signal_18786 ;
    wire signal_18787 ;
    wire signal_18788 ;
    wire signal_18789 ;
    wire signal_18790 ;
    wire signal_18791 ;
    wire signal_18792 ;
    wire signal_18793 ;
    wire signal_18794 ;
    wire signal_18795 ;
    wire signal_18796 ;
    wire signal_18797 ;
    wire signal_18798 ;
    wire signal_18799 ;
    wire signal_18800 ;
    wire signal_18801 ;
    wire signal_18802 ;
    wire signal_18803 ;
    wire signal_18804 ;
    wire signal_18805 ;
    wire signal_18806 ;
    wire signal_18807 ;
    wire signal_18808 ;
    wire signal_18809 ;
    wire signal_18810 ;
    wire signal_18811 ;
    wire signal_18812 ;
    wire signal_18813 ;
    wire signal_18814 ;
    wire signal_18815 ;
    wire signal_18816 ;
    wire signal_18817 ;
    wire signal_18818 ;
    wire signal_18819 ;
    wire signal_18820 ;
    wire signal_18821 ;
    wire signal_18822 ;
    wire signal_18823 ;
    wire signal_18824 ;
    wire signal_18825 ;
    wire signal_18826 ;
    wire signal_18827 ;
    wire signal_18828 ;
    wire signal_18829 ;
    wire signal_18830 ;
    wire signal_18831 ;
    wire signal_18832 ;
    wire signal_18833 ;
    wire signal_18834 ;
    wire signal_18835 ;
    wire signal_18836 ;
    wire signal_18837 ;
    wire signal_18838 ;
    wire signal_18839 ;
    wire signal_18840 ;
    wire signal_18841 ;
    wire signal_18842 ;
    wire signal_18843 ;
    wire signal_18844 ;
    wire signal_18845 ;
    wire signal_18846 ;
    wire signal_18847 ;
    wire signal_18848 ;
    wire signal_18849 ;
    wire signal_18850 ;
    wire signal_18851 ;
    wire signal_18852 ;
    wire signal_18853 ;
    wire signal_18854 ;
    wire signal_18855 ;
    wire signal_18856 ;
    wire signal_18857 ;
    wire signal_18858 ;
    wire signal_18859 ;
    wire signal_18860 ;
    wire signal_18861 ;
    wire signal_18862 ;
    wire signal_18863 ;
    wire signal_18864 ;
    wire signal_18865 ;
    wire signal_18866 ;
    wire signal_18867 ;
    wire signal_18868 ;
    wire signal_18869 ;
    wire signal_18870 ;
    wire signal_18871 ;
    wire signal_18872 ;
    wire signal_18873 ;
    wire signal_18874 ;
    wire signal_18875 ;
    wire signal_18876 ;
    wire signal_18877 ;
    wire signal_18878 ;
    wire signal_18879 ;
    wire signal_18880 ;
    wire signal_18881 ;
    wire signal_18882 ;
    wire signal_18883 ;
    wire signal_18884 ;
    wire signal_18885 ;
    wire signal_18886 ;
    wire signal_18887 ;
    wire signal_18888 ;
    wire signal_18889 ;
    wire signal_18890 ;
    wire signal_18891 ;
    wire signal_18892 ;
    wire signal_18893 ;
    wire signal_18894 ;
    wire signal_18895 ;
    wire signal_18896 ;
    wire signal_18897 ;
    wire signal_18898 ;
    wire signal_18899 ;
    wire signal_18900 ;
    wire signal_18901 ;
    wire signal_18902 ;
    wire signal_18903 ;
    wire signal_18904 ;
    wire signal_18905 ;
    wire signal_18906 ;
    wire signal_18907 ;
    wire signal_18908 ;
    wire signal_18909 ;
    wire signal_18910 ;
    wire signal_18911 ;
    wire signal_18912 ;
    wire signal_18913 ;
    wire signal_18914 ;
    wire signal_18915 ;
    wire signal_18916 ;
    wire signal_18917 ;
    wire signal_18918 ;
    wire signal_18919 ;
    wire signal_18920 ;
    wire signal_18921 ;
    wire signal_18922 ;
    wire signal_18923 ;
    wire signal_18924 ;
    wire signal_18925 ;
    wire signal_18926 ;
    wire signal_18927 ;
    wire signal_18928 ;
    wire signal_18929 ;
    wire signal_18930 ;
    wire signal_18931 ;
    wire signal_18932 ;
    wire signal_18933 ;
    wire signal_18934 ;
    wire signal_18935 ;
    wire signal_18936 ;
    wire signal_18937 ;
    wire signal_18938 ;
    wire signal_18939 ;
    wire signal_18940 ;
    wire signal_18941 ;
    wire signal_18942 ;
    wire signal_18943 ;
    wire signal_18944 ;
    wire signal_18945 ;
    wire signal_18946 ;
    wire signal_18947 ;
    wire signal_18948 ;
    wire signal_18949 ;
    wire signal_18950 ;
    wire signal_18951 ;
    wire signal_18952 ;
    wire signal_18953 ;
    wire signal_18954 ;
    wire signal_18955 ;
    wire signal_18956 ;
    wire signal_18957 ;
    wire signal_18958 ;
    wire signal_18959 ;
    wire signal_18960 ;
    wire signal_18961 ;
    wire signal_18962 ;
    wire signal_18963 ;
    wire signal_18964 ;
    wire signal_18965 ;
    wire signal_18966 ;
    wire signal_18967 ;
    wire signal_18968 ;
    wire signal_18969 ;
    wire signal_18970 ;
    wire signal_18971 ;
    wire signal_18972 ;
    wire signal_18973 ;
    wire signal_18974 ;
    wire signal_18975 ;
    wire signal_18976 ;
    wire signal_18977 ;
    wire signal_18978 ;
    wire signal_18979 ;
    wire signal_18980 ;
    wire signal_18981 ;
    wire signal_18982 ;
    wire signal_18983 ;
    wire signal_18984 ;
    wire signal_18985 ;
    wire signal_18986 ;
    wire signal_18987 ;
    wire signal_18988 ;
    wire signal_18989 ;
    wire signal_18990 ;
    wire signal_18991 ;
    wire signal_18992 ;
    wire signal_18993 ;
    wire signal_18994 ;
    wire signal_18995 ;
    wire signal_18996 ;
    wire signal_18997 ;
    wire signal_18998 ;
    wire signal_18999 ;
    wire signal_19000 ;
    wire signal_19001 ;
    wire signal_19002 ;
    wire signal_19003 ;
    wire signal_19004 ;
    wire signal_19005 ;
    wire signal_19006 ;
    wire signal_19007 ;
    wire signal_19008 ;
    wire signal_19009 ;
    wire signal_19010 ;
    wire signal_19011 ;
    wire signal_19012 ;
    wire signal_19013 ;
    wire signal_19014 ;
    wire signal_19015 ;
    wire signal_19016 ;
    wire signal_19017 ;
    wire signal_19018 ;
    wire signal_19019 ;
    wire signal_19020 ;
    wire signal_19021 ;
    wire signal_19022 ;
    wire signal_19023 ;
    wire signal_19024 ;
    wire signal_19025 ;
    wire signal_19026 ;
    wire signal_19027 ;
    wire signal_19028 ;
    wire signal_19029 ;
    wire signal_19030 ;
    wire signal_19031 ;
    wire signal_19032 ;
    wire signal_19033 ;
    wire signal_19034 ;
    wire signal_19035 ;
    wire signal_19036 ;
    wire signal_19037 ;
    wire signal_19038 ;
    wire signal_19039 ;
    wire signal_19040 ;
    wire signal_19041 ;
    wire signal_19042 ;
    wire signal_19043 ;
    wire signal_19044 ;
    wire signal_19045 ;
    wire signal_19046 ;
    wire signal_19047 ;
    wire signal_19048 ;
    wire signal_19049 ;
    wire signal_19050 ;
    wire signal_19051 ;
    wire signal_19052 ;
    wire signal_19053 ;
    wire signal_19054 ;
    wire signal_19055 ;
    wire signal_19056 ;
    wire signal_19057 ;
    wire signal_19058 ;
    wire signal_19059 ;
    wire signal_19060 ;
    wire signal_19061 ;
    wire signal_19062 ;
    wire signal_19063 ;
    wire signal_19064 ;
    wire signal_19065 ;
    wire signal_19066 ;
    wire signal_19067 ;
    wire signal_19068 ;
    wire signal_19069 ;
    wire signal_19070 ;
    wire signal_19071 ;
    wire signal_19072 ;
    wire signal_19073 ;
    wire signal_19074 ;
    wire signal_19075 ;
    wire signal_19076 ;
    wire signal_19077 ;
    wire signal_19078 ;
    wire signal_19079 ;
    wire signal_19080 ;
    wire signal_19081 ;
    wire signal_19082 ;
    wire signal_19083 ;
    wire signal_19084 ;
    wire signal_19085 ;
    wire signal_19086 ;
    wire signal_19087 ;
    wire signal_19088 ;
    wire signal_19089 ;
    wire signal_19090 ;
    wire signal_19091 ;
    wire signal_19092 ;
    wire signal_19093 ;
    wire signal_19094 ;
    wire signal_19095 ;
    wire signal_19096 ;
    wire signal_19097 ;
    wire signal_19098 ;
    wire signal_19099 ;
    wire signal_19100 ;
    wire signal_19101 ;
    wire signal_19102 ;
    wire signal_19103 ;
    wire signal_19104 ;
    wire signal_19105 ;
    wire signal_19106 ;
    wire signal_19107 ;
    wire signal_19108 ;
    wire signal_19109 ;
    wire signal_19110 ;
    wire signal_19111 ;
    wire signal_19112 ;
    wire signal_19113 ;
    wire signal_19114 ;
    wire signal_19115 ;
    wire signal_19116 ;
    wire signal_19117 ;
    wire signal_19118 ;
    wire signal_19119 ;
    wire signal_19120 ;
    wire signal_19121 ;
    wire signal_19122 ;
    wire signal_19123 ;
    wire signal_19124 ;
    wire signal_19125 ;
    wire signal_19126 ;
    wire signal_19127 ;
    wire signal_19128 ;
    wire signal_19129 ;
    wire signal_19130 ;
    wire signal_19131 ;
    wire signal_19132 ;
    wire signal_19133 ;
    wire signal_19134 ;
    wire signal_19135 ;
    wire signal_19136 ;
    wire signal_19137 ;
    wire signal_19138 ;
    wire signal_19139 ;
    wire signal_19140 ;
    wire signal_19141 ;
    wire signal_19142 ;
    wire signal_19143 ;
    wire signal_19144 ;
    wire signal_19145 ;
    wire signal_19146 ;
    wire signal_19147 ;
    wire signal_19148 ;
    wire signal_19149 ;
    wire signal_19150 ;
    wire signal_19151 ;
    wire signal_19152 ;
    wire signal_19153 ;
    wire signal_19154 ;
    wire signal_19155 ;
    wire signal_19156 ;
    wire signal_19157 ;
    wire signal_19158 ;
    wire signal_19159 ;
    wire signal_19160 ;
    wire signal_19161 ;
    wire signal_19162 ;
    wire signal_19163 ;
    wire signal_19164 ;
    wire signal_19165 ;
    wire signal_19166 ;
    wire signal_19167 ;
    wire signal_19168 ;
    wire signal_19169 ;
    wire signal_19170 ;
    wire signal_19171 ;
    wire signal_19172 ;
    wire signal_19173 ;
    wire signal_19174 ;
    wire signal_19175 ;
    wire signal_19176 ;
    wire signal_19177 ;
    wire signal_19178 ;
    wire signal_19179 ;
    wire signal_19180 ;
    wire signal_19181 ;
    wire signal_19182 ;
    wire signal_19183 ;
    wire signal_19184 ;
    wire signal_19185 ;
    wire signal_19186 ;
    wire signal_19187 ;
    wire signal_19188 ;
    wire signal_19189 ;
    wire signal_19190 ;
    wire signal_19191 ;
    wire signal_19192 ;
    wire signal_19193 ;
    wire signal_19194 ;
    wire signal_19195 ;
    wire signal_19196 ;
    wire signal_19197 ;
    wire signal_19198 ;
    wire signal_19199 ;
    wire signal_19200 ;
    wire signal_19201 ;
    wire signal_19202 ;
    wire signal_19203 ;
    wire signal_19204 ;
    wire signal_19205 ;
    wire signal_19206 ;
    wire signal_19207 ;
    wire signal_19208 ;
    wire signal_19209 ;
    wire signal_19210 ;
    wire signal_19211 ;
    wire signal_19212 ;
    wire signal_19213 ;
    wire signal_19214 ;
    wire signal_19215 ;
    wire signal_19216 ;
    wire signal_19217 ;
    wire signal_19218 ;
    wire signal_19219 ;
    wire signal_19220 ;
    wire signal_19221 ;
    wire signal_19222 ;
    wire signal_19223 ;
    wire signal_19224 ;
    wire signal_19225 ;
    wire signal_19226 ;
    wire signal_19227 ;
    wire signal_19228 ;
    wire signal_19229 ;
    wire signal_19230 ;
    wire signal_19231 ;
    wire signal_19232 ;
    wire signal_19233 ;
    wire signal_19234 ;
    wire signal_19235 ;
    wire signal_19236 ;
    wire signal_19237 ;
    wire signal_19238 ;
    wire signal_19239 ;
    wire signal_19240 ;
    wire signal_19241 ;
    wire signal_19242 ;
    wire signal_19243 ;
    wire signal_19244 ;
    wire signal_19245 ;
    wire signal_19246 ;
    wire signal_19247 ;
    wire signal_19248 ;
    wire signal_19249 ;
    wire signal_19250 ;
    wire signal_19251 ;
    wire signal_19252 ;
    wire signal_19253 ;
    wire signal_19254 ;
    wire signal_19255 ;
    wire signal_19256 ;
    wire signal_19257 ;
    wire signal_19258 ;
    wire signal_19259 ;
    wire signal_19260 ;
    wire signal_19261 ;
    wire signal_19262 ;
    wire signal_19263 ;
    wire signal_19264 ;
    wire signal_19265 ;
    wire signal_19266 ;
    wire signal_19267 ;
    wire signal_19268 ;
    wire signal_19269 ;
    wire signal_19270 ;
    wire signal_19271 ;
    wire signal_19272 ;
    wire signal_19273 ;
    wire signal_19274 ;
    wire signal_19275 ;
    wire signal_19276 ;
    wire signal_19277 ;
    wire signal_19278 ;
    wire signal_19279 ;
    wire signal_19280 ;
    wire signal_19281 ;
    wire signal_19282 ;
    wire signal_19283 ;
    wire signal_19284 ;
    wire signal_19285 ;
    wire signal_19286 ;
    wire signal_19287 ;
    wire signal_19288 ;
    wire signal_19289 ;
    wire signal_19290 ;
    wire signal_19291 ;
    wire signal_19292 ;
    wire signal_19293 ;
    wire signal_19294 ;
    wire signal_19295 ;
    wire signal_19296 ;
    wire signal_19297 ;
    wire signal_19298 ;
    wire signal_19299 ;
    wire signal_19300 ;
    wire signal_19301 ;
    wire signal_19302 ;
    wire signal_19303 ;
    wire signal_19304 ;
    wire signal_19305 ;
    wire signal_19306 ;
    wire signal_19307 ;
    wire signal_19308 ;
    wire signal_19309 ;
    wire signal_19310 ;
    wire signal_19311 ;
    wire signal_19312 ;
    wire signal_19313 ;
    wire signal_19314 ;
    wire signal_19315 ;
    wire signal_19316 ;
    wire signal_19317 ;
    wire signal_19318 ;
    wire signal_19319 ;
    wire signal_19320 ;
    wire signal_19321 ;
    wire signal_19322 ;
    wire signal_19323 ;
    wire signal_19324 ;
    wire signal_19325 ;
    wire signal_19326 ;
    wire signal_19327 ;
    wire signal_19328 ;
    wire signal_19329 ;
    wire signal_19330 ;
    wire signal_19331 ;
    wire signal_19332 ;
    wire signal_19333 ;
    wire signal_19334 ;
    wire signal_19335 ;
    wire signal_19336 ;
    wire signal_19337 ;
    wire signal_19338 ;
    wire signal_19339 ;
    wire signal_19340 ;
    wire signal_19341 ;
    wire signal_19342 ;
    wire signal_19343 ;
    wire signal_19344 ;
    wire signal_19345 ;
    wire signal_19346 ;
    wire signal_19347 ;
    wire signal_19348 ;
    wire signal_19349 ;
    wire signal_19350 ;
    wire signal_19351 ;
    wire signal_19352 ;
    wire signal_19353 ;
    wire signal_19354 ;
    wire signal_19355 ;
    wire signal_19356 ;
    wire signal_19357 ;
    wire signal_19358 ;
    wire signal_19359 ;
    wire signal_19360 ;
    wire signal_19361 ;
    wire signal_19362 ;
    wire signal_19363 ;
    wire signal_19364 ;
    wire signal_19365 ;
    wire signal_19366 ;
    wire signal_19367 ;
    wire signal_19368 ;
    wire signal_19369 ;
    wire signal_19370 ;
    wire signal_19371 ;
    wire signal_19372 ;
    wire signal_19373 ;
    wire signal_19374 ;
    wire signal_19375 ;
    wire signal_19376 ;
    wire signal_19377 ;
    wire signal_19378 ;
    wire signal_19379 ;
    wire signal_19380 ;
    wire signal_19381 ;
    wire signal_19382 ;
    wire signal_19383 ;
    wire signal_19384 ;
    wire signal_19385 ;
    wire signal_19386 ;
    wire signal_19387 ;
    wire signal_19388 ;
    wire signal_19389 ;
    wire signal_19390 ;
    wire signal_19391 ;
    wire signal_19392 ;
    wire signal_19393 ;
    wire signal_19394 ;
    wire signal_19395 ;
    wire signal_19396 ;
    wire signal_19397 ;
    wire signal_19398 ;
    wire signal_19399 ;
    wire signal_19400 ;
    wire signal_19401 ;
    wire signal_19402 ;
    wire signal_19403 ;
    wire signal_19404 ;
    wire signal_19405 ;
    wire signal_19406 ;
    wire signal_19407 ;
    wire signal_19408 ;
    wire signal_19409 ;
    wire signal_19410 ;
    wire signal_19411 ;
    wire signal_19412 ;
    wire signal_19413 ;
    wire signal_19414 ;
    wire signal_19415 ;
    wire signal_19416 ;
    wire signal_19417 ;
    wire signal_19418 ;
    wire signal_19419 ;
    wire signal_19420 ;
    wire signal_19421 ;
    wire signal_19422 ;
    wire signal_19423 ;
    wire signal_19424 ;
    wire signal_19425 ;
    wire signal_19426 ;
    wire signal_19427 ;
    wire signal_19428 ;
    wire signal_19429 ;
    wire signal_19430 ;
    wire signal_19431 ;
    wire signal_19432 ;
    wire signal_19433 ;
    wire signal_19434 ;
    wire signal_19435 ;
    wire signal_19436 ;
    wire signal_19437 ;
    wire signal_19438 ;
    wire signal_19439 ;
    wire signal_19440 ;
    wire signal_19441 ;
    wire signal_19442 ;
    wire signal_19443 ;
    wire signal_19444 ;
    wire signal_19445 ;
    wire signal_19446 ;
    wire signal_19447 ;
    wire signal_19448 ;
    wire signal_19449 ;
    wire signal_19450 ;
    wire signal_19451 ;
    wire signal_19452 ;
    wire signal_19453 ;
    wire signal_19454 ;
    wire signal_19455 ;
    wire signal_19456 ;
    wire signal_19457 ;
    wire signal_19458 ;
    wire signal_19459 ;
    wire signal_19460 ;
    wire signal_19461 ;
    wire signal_19462 ;
    wire signal_19463 ;
    wire signal_19464 ;
    wire signal_19465 ;
    wire signal_19466 ;
    wire signal_19467 ;
    wire signal_19468 ;
    wire signal_19469 ;
    wire signal_19470 ;
    wire signal_19471 ;
    wire signal_19472 ;
    wire signal_19473 ;
    wire signal_19474 ;
    wire signal_19475 ;
    wire signal_19476 ;
    wire signal_19477 ;
    wire signal_19478 ;
    wire signal_19479 ;
    wire signal_19480 ;
    wire signal_19481 ;
    wire signal_19482 ;
    wire signal_19483 ;
    wire signal_19484 ;
    wire signal_19485 ;
    wire signal_19486 ;
    wire signal_19487 ;
    wire signal_19488 ;
    wire signal_19489 ;
    wire signal_19490 ;
    wire signal_19491 ;
    wire signal_19492 ;
    wire signal_19493 ;
    wire signal_19494 ;
    wire signal_19495 ;
    wire signal_19496 ;
    wire signal_19497 ;
    wire signal_19498 ;
    wire signal_19499 ;
    wire signal_19500 ;
    wire signal_19501 ;
    wire signal_19502 ;
    wire signal_19503 ;
    wire signal_19504 ;
    wire signal_19505 ;
    wire signal_19506 ;
    wire signal_19507 ;
    wire signal_19508 ;
    wire signal_19509 ;
    wire signal_19510 ;
    wire signal_19511 ;
    wire signal_19512 ;
    wire signal_19513 ;
    wire signal_19514 ;
    wire signal_19515 ;
    wire signal_19516 ;
    wire signal_19517 ;
    wire signal_19518 ;
    wire signal_19519 ;
    wire signal_19520 ;
    wire signal_19521 ;
    wire signal_19522 ;
    wire signal_19523 ;
    wire signal_19524 ;
    wire signal_19525 ;
    wire signal_19526 ;
    wire signal_19527 ;
    wire signal_19528 ;
    wire signal_19529 ;
    wire signal_19530 ;
    wire signal_19531 ;
    wire signal_19532 ;
    wire signal_19533 ;
    wire signal_19534 ;
    wire signal_19535 ;
    wire signal_19536 ;
    wire signal_19537 ;
    wire signal_19538 ;
    wire signal_19539 ;
    wire signal_19540 ;
    wire signal_19541 ;
    wire signal_19542 ;
    wire signal_19543 ;
    wire signal_19544 ;
    wire signal_19545 ;
    wire signal_19546 ;
    wire signal_19547 ;
    wire signal_19548 ;
    wire signal_19549 ;
    wire signal_19550 ;
    wire signal_19551 ;
    wire signal_19552 ;
    wire signal_19553 ;
    wire signal_19554 ;
    wire signal_19555 ;
    wire signal_19556 ;
    wire signal_19557 ;
    wire signal_19558 ;
    wire signal_19559 ;
    wire signal_19560 ;
    wire signal_19561 ;
    wire signal_19562 ;
    wire signal_19563 ;
    wire signal_19564 ;
    wire signal_19565 ;
    wire signal_19566 ;
    wire signal_19567 ;
    wire signal_19568 ;
    wire signal_19569 ;
    wire signal_19570 ;
    wire signal_19571 ;
    wire signal_19572 ;
    wire signal_19573 ;
    wire signal_19574 ;
    wire signal_19575 ;
    wire signal_19576 ;
    wire signal_19577 ;
    wire signal_19578 ;
    wire signal_19579 ;
    wire signal_19580 ;
    wire signal_19581 ;
    wire signal_19582 ;
    wire signal_19583 ;
    wire signal_19584 ;
    wire signal_19585 ;
    wire signal_19586 ;
    wire signal_19587 ;
    wire signal_19588 ;
    wire signal_19589 ;
    wire signal_19590 ;
    wire signal_19591 ;
    wire signal_19592 ;
    wire signal_19593 ;
    wire signal_19594 ;
    wire signal_19595 ;
    wire signal_19596 ;
    wire signal_19597 ;
    wire signal_19598 ;
    wire signal_19599 ;
    wire signal_19600 ;
    wire signal_19601 ;
    wire signal_19602 ;
    wire signal_19603 ;
    wire signal_19604 ;
    wire signal_19605 ;
    wire signal_19606 ;
    wire signal_19607 ;
    wire signal_19608 ;
    wire signal_19609 ;
    wire signal_19610 ;
    wire signal_19611 ;
    wire signal_19612 ;
    wire signal_19613 ;
    wire signal_19614 ;
    wire signal_19615 ;
    wire signal_19616 ;
    wire signal_19617 ;
    wire signal_19618 ;
    wire signal_19619 ;
    wire signal_19620 ;
    wire signal_19621 ;
    wire signal_19622 ;
    wire signal_19623 ;
    wire signal_19624 ;
    wire signal_19625 ;
    wire signal_19626 ;
    wire signal_19627 ;
    wire signal_19628 ;
    wire signal_19629 ;
    wire signal_19630 ;
    wire signal_19631 ;
    wire signal_19632 ;
    wire signal_19633 ;
    wire signal_19634 ;
    wire signal_19635 ;
    wire signal_19636 ;
    wire signal_19637 ;
    wire signal_19638 ;
    wire signal_19639 ;
    wire signal_19640 ;
    wire signal_19641 ;
    wire signal_19642 ;
    wire signal_19643 ;
    wire signal_19644 ;
    wire signal_19645 ;
    wire signal_19646 ;
    wire signal_19647 ;
    wire signal_19648 ;
    wire signal_19649 ;
    wire signal_19650 ;
    wire signal_19651 ;
    wire signal_19652 ;
    wire signal_19653 ;
    wire signal_19654 ;
    wire signal_19655 ;
    wire signal_19656 ;
    wire signal_19657 ;
    wire signal_19658 ;
    wire signal_19659 ;
    wire signal_19660 ;
    wire signal_19661 ;
    wire signal_19662 ;
    wire signal_19663 ;
    wire signal_19664 ;
    wire signal_19665 ;
    wire signal_19666 ;
    wire signal_19667 ;
    wire signal_19668 ;
    wire signal_19669 ;
    wire signal_19670 ;
    wire signal_19671 ;
    wire signal_19672 ;
    wire signal_19673 ;
    wire signal_19674 ;
    wire signal_19675 ;
    wire signal_19676 ;
    wire signal_19677 ;
    wire signal_19678 ;
    wire signal_19679 ;
    wire signal_19680 ;
    wire signal_19681 ;
    wire signal_19682 ;
    wire signal_19683 ;
    wire signal_19684 ;
    wire signal_19685 ;
    wire signal_19686 ;
    wire signal_19687 ;
    wire signal_19688 ;
    wire signal_19689 ;
    wire signal_19690 ;
    wire signal_19691 ;
    wire signal_19692 ;
    wire signal_19693 ;
    wire signal_19694 ;
    wire signal_19695 ;
    wire signal_19696 ;
    wire signal_19697 ;
    wire signal_19698 ;
    wire signal_19699 ;
    wire signal_19700 ;
    wire signal_19701 ;
    wire signal_19702 ;
    wire signal_19703 ;
    wire signal_19704 ;
    wire signal_19705 ;
    wire signal_19706 ;
    wire signal_19707 ;
    wire signal_19708 ;
    wire signal_19709 ;
    wire signal_19710 ;
    wire signal_19711 ;
    wire signal_19712 ;
    wire signal_19713 ;
    wire signal_19714 ;
    wire signal_19715 ;
    wire signal_19716 ;
    wire signal_19717 ;
    wire signal_19718 ;
    wire signal_19719 ;
    wire signal_19720 ;
    wire signal_19721 ;
    wire signal_19722 ;
    wire signal_19723 ;
    wire signal_19724 ;
    wire signal_19725 ;
    wire signal_19726 ;
    wire signal_19727 ;
    wire signal_19728 ;
    wire signal_19729 ;
    wire signal_19730 ;
    wire signal_19731 ;
    wire signal_19732 ;
    wire signal_19733 ;
    wire signal_19734 ;
    wire signal_19735 ;
    wire signal_19736 ;
    wire signal_19737 ;
    wire signal_19738 ;
    wire signal_19739 ;
    wire signal_19740 ;
    wire signal_19741 ;
    wire signal_19742 ;
    wire signal_19743 ;
    wire signal_19744 ;
    wire signal_19745 ;
    wire signal_19746 ;
    wire signal_19747 ;
    wire signal_19748 ;
    wire signal_19749 ;
    wire signal_19750 ;
    wire signal_19751 ;
    wire signal_19752 ;
    wire signal_19753 ;
    wire signal_19754 ;
    wire signal_19755 ;
    wire signal_19756 ;
    wire signal_19757 ;
    wire signal_19758 ;
    wire signal_19759 ;
    wire signal_19760 ;
    wire signal_19761 ;
    wire signal_19762 ;
    wire signal_19763 ;
    wire signal_19764 ;
    wire signal_19765 ;
    wire signal_19766 ;
    wire signal_19767 ;
    wire signal_19768 ;
    wire signal_19769 ;
    wire signal_19770 ;
    wire signal_19771 ;
    wire signal_19772 ;
    wire signal_19773 ;
    wire signal_19774 ;
    wire signal_19775 ;
    wire signal_19776 ;
    wire signal_19777 ;
    wire signal_19778 ;
    wire signal_19779 ;
    wire signal_19780 ;
    wire signal_19781 ;
    wire signal_19782 ;
    wire signal_19783 ;
    wire signal_19784 ;
    wire signal_19785 ;
    wire signal_19786 ;
    wire signal_19787 ;
    wire signal_19788 ;
    wire signal_19789 ;
    wire signal_19790 ;
    wire signal_19791 ;
    wire signal_19792 ;
    wire signal_19793 ;
    wire signal_19794 ;
    wire signal_19795 ;
    wire signal_19796 ;
    wire signal_19797 ;
    wire signal_19798 ;
    wire signal_19799 ;
    wire signal_19800 ;
    wire signal_19801 ;
    wire signal_19802 ;
    wire signal_19803 ;
    wire signal_19804 ;
    wire signal_19805 ;
    wire signal_19806 ;
    wire signal_19807 ;
    wire signal_19808 ;
    wire signal_19809 ;
    wire signal_19810 ;
    wire signal_19811 ;
    wire signal_19812 ;
    wire signal_19813 ;
    wire signal_19814 ;
    wire signal_19815 ;
    wire signal_19816 ;
    wire signal_19817 ;
    wire signal_19818 ;
    wire signal_19819 ;
    wire signal_19820 ;
    wire signal_19821 ;
    wire signal_19822 ;
    wire signal_19823 ;
    wire signal_19824 ;
    wire signal_19825 ;
    wire signal_19826 ;
    wire signal_19827 ;
    wire signal_19828 ;
    wire signal_19829 ;
    wire signal_19830 ;
    wire signal_19831 ;
    wire signal_19832 ;
    wire signal_19833 ;
    wire signal_19834 ;
    wire signal_19835 ;
    wire signal_19836 ;
    wire signal_19837 ;
    wire signal_19838 ;
    wire signal_19839 ;
    wire signal_19840 ;
    wire signal_19841 ;
    wire signal_19842 ;
    wire signal_19843 ;
    wire signal_19844 ;
    wire signal_19845 ;
    wire signal_19846 ;
    wire signal_19847 ;
    wire signal_19848 ;
    wire signal_19849 ;
    wire signal_19850 ;
    wire signal_19851 ;
    wire signal_19852 ;
    wire signal_19853 ;
    wire signal_19854 ;
    wire signal_19855 ;
    wire signal_19856 ;
    wire signal_19857 ;
    wire signal_19858 ;
    wire signal_19859 ;
    wire signal_19860 ;
    wire signal_19861 ;
    wire signal_19862 ;
    wire signal_19863 ;
    wire signal_19864 ;
    wire signal_19865 ;
    wire signal_19866 ;
    wire signal_19867 ;
    wire signal_19868 ;
    wire signal_19869 ;
    wire signal_19870 ;
    wire signal_19871 ;
    wire signal_19872 ;
    wire signal_19873 ;
    wire signal_19874 ;
    wire signal_19875 ;
    wire signal_19876 ;
    wire signal_19877 ;
    wire signal_19878 ;
    wire signal_19879 ;
    wire signal_19880 ;
    wire signal_19881 ;
    wire signal_19882 ;
    wire signal_19883 ;
    wire signal_19884 ;
    wire signal_19885 ;
    wire signal_19886 ;
    wire signal_19887 ;
    wire signal_19888 ;
    wire signal_19889 ;
    wire signal_19890 ;
    wire signal_19891 ;
    wire signal_19892 ;
    wire signal_19893 ;
    wire signal_19894 ;
    wire signal_19895 ;
    wire signal_19896 ;
    wire signal_19897 ;
    wire signal_19898 ;
    wire signal_19899 ;
    wire signal_19900 ;
    wire signal_19901 ;
    wire signal_19902 ;
    wire signal_19903 ;
    wire signal_19904 ;
    wire signal_19905 ;
    wire signal_19906 ;
    wire signal_19907 ;
    wire signal_19908 ;
    wire signal_19909 ;
    wire signal_19910 ;
    wire signal_19911 ;
    wire signal_19912 ;
    wire signal_19913 ;
    wire signal_19914 ;
    wire signal_19915 ;
    wire signal_19916 ;
    wire signal_19917 ;
    wire signal_19918 ;
    wire signal_19919 ;
    wire signal_19920 ;
    wire signal_19921 ;
    wire signal_19922 ;
    wire signal_19923 ;
    wire signal_19924 ;
    wire signal_19925 ;
    wire signal_19926 ;
    wire signal_19927 ;
    wire signal_19928 ;
    wire signal_19929 ;
    wire signal_19930 ;
    wire signal_19931 ;
    wire signal_19932 ;
    wire signal_19933 ;
    wire signal_19934 ;
    wire signal_19935 ;
    wire signal_19936 ;
    wire signal_19937 ;
    wire signal_19938 ;
    wire signal_19939 ;
    wire signal_19940 ;
    wire signal_19941 ;
    wire signal_19942 ;
    wire signal_19943 ;
    wire signal_19944 ;
    wire signal_19945 ;
    wire signal_19946 ;
    wire signal_19947 ;
    wire signal_19948 ;
    wire signal_19949 ;
    wire signal_19950 ;
    wire signal_19951 ;
    wire signal_19952 ;
    wire signal_19953 ;
    wire signal_19954 ;
    wire signal_19955 ;
    wire signal_19956 ;
    wire signal_19957 ;
    wire signal_19958 ;
    wire signal_19959 ;
    wire signal_19960 ;
    wire signal_19961 ;
    wire signal_19962 ;
    wire signal_19963 ;
    wire signal_19964 ;
    wire signal_19965 ;
    wire signal_19966 ;
    wire signal_19967 ;
    wire signal_19968 ;
    wire signal_19969 ;
    wire signal_19970 ;
    wire signal_19971 ;
    wire signal_19972 ;
    wire signal_19973 ;
    wire signal_19974 ;
    wire signal_19975 ;
    wire signal_19976 ;
    wire signal_19977 ;
    wire signal_19978 ;
    wire signal_19979 ;
    wire signal_19980 ;
    wire signal_19981 ;
    wire signal_19982 ;
    wire signal_19983 ;
    wire signal_19984 ;
    wire signal_19985 ;
    wire signal_19986 ;
    wire signal_19987 ;
    wire signal_19988 ;
    wire signal_19989 ;
    wire signal_19990 ;
    wire signal_19991 ;
    wire signal_19992 ;
    wire signal_19993 ;
    wire signal_19994 ;
    wire signal_19995 ;
    wire signal_19996 ;
    wire signal_19997 ;
    wire signal_19998 ;
    wire signal_19999 ;
    wire signal_20000 ;
    wire signal_20001 ;
    wire signal_20002 ;
    wire signal_20003 ;
    wire signal_20004 ;
    wire signal_20005 ;
    wire signal_20006 ;
    wire signal_20007 ;
    wire signal_20008 ;
    wire signal_20009 ;
    wire signal_20010 ;
    wire signal_20011 ;
    wire signal_20012 ;
    wire signal_20013 ;
    wire signal_20014 ;
    wire signal_20015 ;
    wire signal_20016 ;
    wire signal_20017 ;
    wire signal_20018 ;
    wire signal_20019 ;
    wire signal_20020 ;
    wire signal_20021 ;
    wire signal_20022 ;
    wire signal_20023 ;
    wire signal_20024 ;
    wire signal_20025 ;
    wire signal_20026 ;
    wire signal_20027 ;
    wire signal_20028 ;
    wire signal_20029 ;
    wire signal_20030 ;
    wire signal_20031 ;
    wire signal_20032 ;
    wire signal_20033 ;
    wire signal_20034 ;
    wire signal_20035 ;
    wire signal_20036 ;
    wire signal_20037 ;
    wire signal_20038 ;
    wire signal_20039 ;
    wire signal_20040 ;
    wire signal_20041 ;
    wire signal_20042 ;
    wire signal_20043 ;
    wire signal_20044 ;
    wire signal_20045 ;
    wire signal_20046 ;
    wire signal_20047 ;
    wire signal_20048 ;
    wire signal_20049 ;
    wire signal_20050 ;
    wire signal_20051 ;
    wire signal_20052 ;
    wire signal_20053 ;
    wire signal_20054 ;
    wire signal_20055 ;
    wire signal_20056 ;
    wire signal_20057 ;
    wire signal_20058 ;
    wire signal_20059 ;
    wire signal_20060 ;
    wire signal_20061 ;
    wire signal_20062 ;
    wire signal_20063 ;
    wire signal_20064 ;
    wire signal_20065 ;
    wire signal_20066 ;
    wire signal_20067 ;
    wire signal_20068 ;
    wire signal_20069 ;
    wire signal_20070 ;
    wire signal_20071 ;
    wire signal_20072 ;
    wire signal_20073 ;
    wire signal_20074 ;
    wire signal_20075 ;
    wire signal_20076 ;
    wire signal_20077 ;
    wire signal_20078 ;
    wire signal_20079 ;
    wire signal_20080 ;
    wire signal_20081 ;
    wire signal_20082 ;
    wire signal_20083 ;
    wire signal_20084 ;
    wire signal_20085 ;
    wire signal_20086 ;
    wire signal_20087 ;
    wire signal_20088 ;
    wire signal_20089 ;
    wire signal_20090 ;
    wire signal_20091 ;
    wire signal_20092 ;
    wire signal_20093 ;
    wire signal_20094 ;
    wire signal_20095 ;
    wire signal_20096 ;
    wire signal_20097 ;
    wire signal_20098 ;
    wire signal_20099 ;
    wire signal_20100 ;
    wire signal_20101 ;
    wire signal_20102 ;
    wire signal_20103 ;
    wire signal_20104 ;
    wire signal_20105 ;
    wire signal_20106 ;
    wire signal_20107 ;
    wire signal_20108 ;
    wire signal_20109 ;
    wire signal_20110 ;
    wire signal_20111 ;
    wire signal_20112 ;
    wire signal_20113 ;
    wire signal_20114 ;
    wire signal_20115 ;
    wire signal_20116 ;
    wire signal_20117 ;
    wire signal_20118 ;
    wire signal_20119 ;
    wire signal_20120 ;
    wire signal_20121 ;
    wire signal_20122 ;
    wire signal_20123 ;
    wire signal_20124 ;
    wire signal_20125 ;
    wire signal_20126 ;
    wire signal_20127 ;
    wire signal_20128 ;
    wire signal_20129 ;
    wire signal_20130 ;
    wire signal_20131 ;
    wire signal_20132 ;
    wire signal_20133 ;
    wire signal_20134 ;
    wire signal_20135 ;
    wire signal_20136 ;
    wire signal_20137 ;
    wire signal_20138 ;
    wire signal_20139 ;
    wire signal_20140 ;
    wire signal_20141 ;
    wire signal_20142 ;
    wire signal_20143 ;
    wire signal_20144 ;
    wire signal_20145 ;
    wire signal_20146 ;
    wire signal_20147 ;
    wire signal_20148 ;
    wire signal_20149 ;
    wire signal_20150 ;
    wire signal_20151 ;
    wire signal_20152 ;
    wire signal_20153 ;
    wire signal_20154 ;
    wire signal_20155 ;
    wire signal_20156 ;
    wire signal_20157 ;
    wire signal_20158 ;
    wire signal_20159 ;
    wire signal_20160 ;
    wire signal_20161 ;
    wire signal_20162 ;
    wire signal_20163 ;
    wire signal_20164 ;
    wire signal_20165 ;
    wire signal_20166 ;
    wire signal_20167 ;
    wire signal_20168 ;
    wire signal_20169 ;
    wire signal_20170 ;
    wire signal_20171 ;
    wire signal_20172 ;
    wire signal_20173 ;
    wire signal_20174 ;
    wire signal_20175 ;
    wire signal_20176 ;
    wire signal_20177 ;
    wire signal_20178 ;
    wire signal_20179 ;
    wire signal_20180 ;
    wire signal_20181 ;
    wire signal_20182 ;
    wire signal_20183 ;
    wire signal_20184 ;
    wire signal_20185 ;
    wire signal_20186 ;
    wire signal_20187 ;
    wire signal_20188 ;
    wire signal_20189 ;
    wire signal_20190 ;
    wire signal_20191 ;
    wire signal_20192 ;
    wire signal_20193 ;
    wire signal_20194 ;
    wire signal_20195 ;
    wire signal_20196 ;
    wire signal_20197 ;
    wire signal_20198 ;
    wire signal_20199 ;
    wire signal_20200 ;
    wire signal_20201 ;
    wire signal_20202 ;
    wire signal_20203 ;
    wire signal_20204 ;
    wire signal_20205 ;
    wire signal_20206 ;
    wire signal_20207 ;
    wire signal_20208 ;
    wire signal_20209 ;
    wire signal_20210 ;
    wire signal_20211 ;
    wire signal_20212 ;
    wire signal_20213 ;
    wire signal_20214 ;
    wire signal_20215 ;
    wire signal_20216 ;
    wire signal_20217 ;
    wire signal_20218 ;
    wire signal_20219 ;
    wire signal_20220 ;
    wire signal_20221 ;
    wire signal_20222 ;
    wire signal_20223 ;
    wire signal_20224 ;
    wire signal_20225 ;
    wire signal_20226 ;
    wire signal_20227 ;
    wire signal_20228 ;
    wire signal_20229 ;
    wire signal_20230 ;
    wire signal_20231 ;
    wire signal_20232 ;
    wire signal_20233 ;
    wire signal_20234 ;
    wire signal_20235 ;
    wire signal_20236 ;
    wire signal_20237 ;
    wire signal_20238 ;
    wire signal_20239 ;
    wire signal_20240 ;
    wire signal_20241 ;
    wire signal_20242 ;
    wire signal_20243 ;
    wire signal_20244 ;
    wire signal_20245 ;
    wire signal_20246 ;
    wire signal_20247 ;
    wire signal_20248 ;
    wire signal_20249 ;
    wire signal_20250 ;
    wire signal_20251 ;
    wire signal_20252 ;
    wire signal_20253 ;
    wire signal_20254 ;
    wire signal_20255 ;
    wire signal_20256 ;
    wire signal_20257 ;
    wire signal_20258 ;
    wire signal_20259 ;
    wire signal_20260 ;
    wire signal_20261 ;
    wire signal_20262 ;
    wire signal_20263 ;
    wire signal_20264 ;
    wire signal_20265 ;
    wire signal_20266 ;
    wire signal_20267 ;
    wire signal_20268 ;
    wire signal_20269 ;
    wire signal_20270 ;
    wire signal_20271 ;
    wire signal_20272 ;
    wire signal_20273 ;
    wire signal_20274 ;
    wire signal_20275 ;
    wire signal_20276 ;
    wire signal_20277 ;
    wire signal_20278 ;
    wire signal_20279 ;
    wire signal_20280 ;
    wire signal_20281 ;
    wire signal_20282 ;
    wire signal_20283 ;
    wire signal_20284 ;
    wire signal_20285 ;
    wire signal_20286 ;
    wire signal_20287 ;
    wire signal_20288 ;
    wire signal_20289 ;
    wire signal_20290 ;
    wire signal_20291 ;
    wire signal_20292 ;
    wire signal_20293 ;
    wire signal_20294 ;
    wire signal_20295 ;
    wire signal_20296 ;
    wire signal_20297 ;
    wire signal_20298 ;
    wire signal_20299 ;
    wire signal_20300 ;
    wire signal_20301 ;
    wire signal_20302 ;
    wire signal_20303 ;
    wire signal_20304 ;
    wire signal_20305 ;
    wire signal_20306 ;
    wire signal_20307 ;
    wire signal_20308 ;
    wire signal_20309 ;
    wire signal_20310 ;
    wire signal_20311 ;
    wire signal_20312 ;
    wire signal_20313 ;
    wire signal_20314 ;
    wire signal_20315 ;
    wire signal_20316 ;
    wire signal_20317 ;
    wire signal_20318 ;
    wire signal_20319 ;
    wire signal_20320 ;
    wire signal_20321 ;
    wire signal_20322 ;
    wire signal_20323 ;
    wire signal_20324 ;
    wire signal_20325 ;
    wire signal_20326 ;
    wire signal_20327 ;
    wire signal_20328 ;
    wire signal_20329 ;
    wire signal_20330 ;
    wire signal_20331 ;
    wire signal_20332 ;
    wire signal_20333 ;
    wire signal_20334 ;
    wire signal_20335 ;
    wire signal_20336 ;
    wire signal_20337 ;
    wire signal_20338 ;
    wire signal_20339 ;
    wire signal_20340 ;
    wire signal_20341 ;
    wire signal_20342 ;
    wire signal_20343 ;
    wire signal_20344 ;
    wire signal_20345 ;
    wire signal_20346 ;
    wire signal_20347 ;
    wire signal_20348 ;
    wire signal_20349 ;
    wire signal_20350 ;
    wire signal_20351 ;
    wire signal_20352 ;
    wire signal_20353 ;
    wire signal_20354 ;
    wire signal_20355 ;
    wire signal_20356 ;
    wire signal_20357 ;
    wire signal_20358 ;
    wire signal_20359 ;
    wire signal_20360 ;
    wire signal_20361 ;
    wire signal_20362 ;
    wire signal_20363 ;
    wire signal_20364 ;
    wire signal_20365 ;
    wire signal_20366 ;
    wire signal_20367 ;
    wire signal_20368 ;
    wire signal_20369 ;
    wire signal_20370 ;
    wire signal_20371 ;
    wire signal_20372 ;
    wire signal_20373 ;
    wire signal_20374 ;
    wire signal_20375 ;
    wire signal_20376 ;
    wire signal_20377 ;
    wire signal_20378 ;
    wire signal_20379 ;
    wire signal_20380 ;
    wire signal_20381 ;
    wire signal_20382 ;
    wire signal_20383 ;
    wire signal_20384 ;
    wire signal_20385 ;
    wire signal_20386 ;
    wire signal_20387 ;
    wire signal_20388 ;
    wire signal_20389 ;
    wire signal_20390 ;
    wire signal_20391 ;
    wire signal_20392 ;
    wire signal_20393 ;
    wire signal_20394 ;
    wire signal_20395 ;
    wire signal_20396 ;
    wire signal_20397 ;
    wire signal_20398 ;
    wire signal_20399 ;
    wire signal_20400 ;
    wire signal_20401 ;
    wire signal_20402 ;
    wire signal_20403 ;
    wire signal_20404 ;
    wire signal_20405 ;
    wire signal_20406 ;
    wire signal_20407 ;
    wire signal_20408 ;
    wire signal_20409 ;
    wire signal_20410 ;
    wire signal_20411 ;
    wire signal_20412 ;
    wire signal_20413 ;
    wire signal_20414 ;
    wire signal_20415 ;
    wire signal_20416 ;
    wire signal_20417 ;
    wire signal_20418 ;
    wire signal_20419 ;
    wire signal_20420 ;
    wire signal_20421 ;
    wire signal_20422 ;
    wire signal_20423 ;
    wire signal_20424 ;
    wire signal_20425 ;
    wire signal_20426 ;
    wire signal_20427 ;
    wire signal_20428 ;
    wire signal_20429 ;
    wire signal_20430 ;
    wire signal_20431 ;
    wire signal_20432 ;
    wire signal_20433 ;
    wire signal_20434 ;
    wire signal_20435 ;
    wire signal_20436 ;
    wire signal_20437 ;
    wire signal_20438 ;
    wire signal_20439 ;
    wire signal_20440 ;
    wire signal_20441 ;
    wire signal_20442 ;
    wire signal_20443 ;
    wire signal_20444 ;
    wire signal_20445 ;
    wire signal_20446 ;
    wire signal_20447 ;
    wire signal_20448 ;
    wire signal_20449 ;
    wire signal_20450 ;
    wire signal_20451 ;
    wire signal_20452 ;
    wire signal_20453 ;
    wire signal_20454 ;
    wire signal_20455 ;
    wire signal_20456 ;
    wire signal_20457 ;
    wire signal_20458 ;
    wire signal_20459 ;
    wire signal_20460 ;
    wire signal_20461 ;
    wire signal_20462 ;
    wire signal_20463 ;
    wire signal_20464 ;
    wire signal_20465 ;
    wire signal_20466 ;
    wire signal_20467 ;
    wire signal_20468 ;
    wire signal_20469 ;
    wire signal_20470 ;
    wire signal_20471 ;
    wire signal_20472 ;
    wire signal_20473 ;
    wire signal_20474 ;
    wire signal_20475 ;
    wire signal_20476 ;
    wire signal_20477 ;
    wire signal_20478 ;
    wire signal_20479 ;
    wire signal_20480 ;
    wire signal_20481 ;
    wire signal_20482 ;
    wire signal_20483 ;
    wire signal_20484 ;
    wire signal_20485 ;
    wire signal_20486 ;
    wire signal_20487 ;
    wire signal_20488 ;
    wire signal_20489 ;
    wire signal_20490 ;
    wire signal_20491 ;
    wire signal_20492 ;
    wire signal_20493 ;
    wire signal_20494 ;
    wire signal_20495 ;
    wire signal_20496 ;
    wire signal_20497 ;
    wire signal_20498 ;
    wire signal_20499 ;
    wire signal_20500 ;
    wire signal_20501 ;
    wire signal_20502 ;
    wire signal_20503 ;
    wire signal_20504 ;
    wire signal_20505 ;
    wire signal_20506 ;
    wire signal_20507 ;
    wire signal_20508 ;
    wire signal_20509 ;
    wire signal_20510 ;
    wire signal_20511 ;
    wire signal_20512 ;
    wire signal_20513 ;
    wire signal_20514 ;
    wire signal_20515 ;
    wire signal_20516 ;
    wire signal_20517 ;
    wire signal_20518 ;
    wire signal_20519 ;
    wire signal_20520 ;
    wire signal_20521 ;
    wire signal_20522 ;
    wire signal_20523 ;
    wire signal_20524 ;
    wire signal_20525 ;
    wire signal_20526 ;
    wire signal_20527 ;
    wire signal_20528 ;
    wire signal_20529 ;
    wire signal_20530 ;
    wire signal_20531 ;
    wire signal_20532 ;
    wire signal_20533 ;
    wire signal_20534 ;
    wire signal_20535 ;
    wire signal_20536 ;
    wire signal_20537 ;
    wire signal_20538 ;
    wire signal_20539 ;
    wire signal_20540 ;
    wire signal_20541 ;
    wire signal_20542 ;
    wire signal_20543 ;
    wire signal_20544 ;
    wire signal_20545 ;
    wire signal_20546 ;
    wire signal_20547 ;
    wire signal_20548 ;
    wire signal_20549 ;
    wire signal_20550 ;
    wire signal_20551 ;
    wire signal_20552 ;
    wire signal_20553 ;
    wire signal_20554 ;
    wire signal_20555 ;
    wire signal_20556 ;
    wire signal_20557 ;
    wire signal_20558 ;
    wire signal_20559 ;
    wire signal_20560 ;
    wire signal_20561 ;
    wire signal_20562 ;
    wire signal_20563 ;
    wire signal_20564 ;
    wire signal_20565 ;
    wire signal_20566 ;
    wire signal_20567 ;
    wire signal_20568 ;
    wire signal_20569 ;
    wire signal_20570 ;
    wire signal_20571 ;
    wire signal_20572 ;
    wire signal_20573 ;
    wire signal_20574 ;
    wire signal_20575 ;
    wire signal_20576 ;
    wire signal_20577 ;
    wire signal_20578 ;
    wire signal_20579 ;
    wire signal_20580 ;
    wire signal_20581 ;
    wire signal_20582 ;
    wire signal_20583 ;
    wire signal_20584 ;
    wire signal_20585 ;
    wire signal_20586 ;
    wire signal_20587 ;
    wire signal_20588 ;
    wire signal_20589 ;
    wire signal_20590 ;
    wire signal_20591 ;
    wire signal_20592 ;
    wire signal_20593 ;
    wire signal_20594 ;
    wire signal_20595 ;
    wire signal_20596 ;
    wire signal_20597 ;
    wire signal_20598 ;
    wire signal_20599 ;
    wire signal_20600 ;
    wire signal_20601 ;
    wire signal_20602 ;
    wire signal_20603 ;
    wire signal_20604 ;
    wire signal_20605 ;
    wire signal_20606 ;
    wire signal_20607 ;
    wire signal_20608 ;
    wire signal_20609 ;
    wire signal_20610 ;
    wire signal_20611 ;
    wire signal_20612 ;
    wire signal_20613 ;
    wire signal_20614 ;
    wire signal_20615 ;
    wire signal_20616 ;
    wire signal_20617 ;
    wire signal_20618 ;
    wire signal_20619 ;
    wire signal_20620 ;
    wire signal_20621 ;
    wire signal_20622 ;
    wire signal_20623 ;
    wire signal_20624 ;
    wire signal_20625 ;
    wire signal_20626 ;
    wire signal_20627 ;
    wire signal_20628 ;
    wire signal_20629 ;
    wire signal_20630 ;
    wire signal_20631 ;
    wire signal_20632 ;
    wire signal_20633 ;
    wire signal_20634 ;
    wire signal_20635 ;
    wire signal_20636 ;
    wire signal_20637 ;
    wire signal_20638 ;
    wire signal_20639 ;
    wire signal_20640 ;
    wire signal_20641 ;
    wire signal_20642 ;
    wire signal_20643 ;
    wire signal_20644 ;
    wire signal_20645 ;
    wire signal_20646 ;
    wire signal_20647 ;
    wire signal_20648 ;
    wire signal_20649 ;
    wire signal_20650 ;
    wire signal_20651 ;
    wire signal_20652 ;
    wire signal_20653 ;
    wire signal_20654 ;
    wire signal_20655 ;
    wire signal_20656 ;
    wire signal_20657 ;
    wire signal_20658 ;
    wire signal_20659 ;
    wire signal_20660 ;
    wire signal_20661 ;
    wire signal_20662 ;
    wire signal_20663 ;
    wire signal_20664 ;
    wire signal_20665 ;
    wire signal_20666 ;
    wire signal_20667 ;
    wire signal_20668 ;
    wire signal_20669 ;
    wire signal_20670 ;
    wire signal_20671 ;
    wire signal_20672 ;
    wire signal_20673 ;
    wire signal_20674 ;
    wire signal_20675 ;
    wire signal_20676 ;
    wire signal_20677 ;
    wire signal_20678 ;
    wire signal_20679 ;
    wire signal_20680 ;
    wire signal_20681 ;
    wire signal_20682 ;
    wire signal_20683 ;
    wire signal_20684 ;
    wire signal_20685 ;
    wire signal_20686 ;
    wire signal_20687 ;
    wire signal_20688 ;
    wire signal_20689 ;
    wire signal_20690 ;
    wire signal_20691 ;
    wire signal_20692 ;
    wire signal_20693 ;
    wire signal_20694 ;
    wire signal_20695 ;
    wire signal_20696 ;
    wire signal_20697 ;
    wire signal_20698 ;
    wire signal_20699 ;
    wire signal_20700 ;
    wire signal_20701 ;
    wire signal_20702 ;
    wire signal_20703 ;
    wire signal_20704 ;
    wire signal_20705 ;
    wire signal_20706 ;
    wire signal_20707 ;
    wire signal_20708 ;
    wire signal_20709 ;
    wire signal_20710 ;
    wire signal_20711 ;
    wire signal_20712 ;
    wire signal_20713 ;
    wire signal_20714 ;
    wire signal_20715 ;
    wire signal_20716 ;
    wire signal_20717 ;
    wire signal_20718 ;
    wire signal_20719 ;
    wire signal_20720 ;
    wire signal_20721 ;
    wire signal_20722 ;
    wire signal_20723 ;
    wire signal_20724 ;
    wire signal_20725 ;
    wire signal_20726 ;
    wire signal_20727 ;
    wire signal_20728 ;
    wire signal_20729 ;
    wire signal_20730 ;
    wire signal_20731 ;
    wire signal_20732 ;
    wire signal_20733 ;
    wire signal_20734 ;
    wire signal_20735 ;
    wire signal_20736 ;
    wire signal_20737 ;
    wire signal_20738 ;
    wire signal_20739 ;
    wire signal_20740 ;
    wire signal_20741 ;
    wire signal_20742 ;
    wire signal_20743 ;
    wire signal_20744 ;
    wire signal_20745 ;
    wire signal_20746 ;
    wire signal_20747 ;
    wire signal_20748 ;
    wire signal_20749 ;
    wire signal_20750 ;
    wire signal_20751 ;
    wire signal_20752 ;
    wire signal_20753 ;
    wire signal_20754 ;
    wire signal_20755 ;
    wire signal_20756 ;
    wire signal_20757 ;
    wire signal_20758 ;
    wire signal_20759 ;
    wire signal_20760 ;
    wire signal_20761 ;
    wire signal_20762 ;
    wire signal_20763 ;
    wire signal_20764 ;
    wire signal_20765 ;
    wire signal_20766 ;
    wire signal_20767 ;
    wire signal_20768 ;
    wire signal_20769 ;
    wire signal_20770 ;
    wire signal_20771 ;
    wire signal_20772 ;
    wire signal_20773 ;
    wire signal_20774 ;
    wire signal_20775 ;
    wire signal_20776 ;
    wire signal_20777 ;
    wire signal_20778 ;
    wire signal_20779 ;
    wire signal_20780 ;
    wire signal_20781 ;
    wire signal_20782 ;
    wire signal_20783 ;
    wire signal_20784 ;
    wire signal_20785 ;
    wire signal_20786 ;
    wire signal_20787 ;
    wire signal_20788 ;
    wire signal_20789 ;
    wire signal_20790 ;
    wire signal_20791 ;
    wire signal_20792 ;
    wire signal_20793 ;
    wire signal_20794 ;
    wire signal_20795 ;
    wire signal_20796 ;
    wire signal_20797 ;
    wire signal_20798 ;
    wire signal_20799 ;
    wire signal_20800 ;
    wire signal_20801 ;
    wire signal_20802 ;
    wire signal_20803 ;
    wire signal_20804 ;
    wire signal_20805 ;
    wire signal_20806 ;
    wire signal_20807 ;
    wire signal_20808 ;
    wire signal_20809 ;
    wire signal_20810 ;
    wire signal_20811 ;
    wire signal_20812 ;
    wire signal_20813 ;
    wire signal_20814 ;
    wire signal_20815 ;
    wire signal_20816 ;
    wire signal_20817 ;
    wire signal_20818 ;
    wire signal_20819 ;
    wire signal_20820 ;
    wire signal_20821 ;
    wire signal_20822 ;
    wire signal_20823 ;
    wire signal_20824 ;
    wire signal_20825 ;
    wire signal_20826 ;
    wire signal_20827 ;
    wire signal_20828 ;
    wire signal_20829 ;
    wire signal_20830 ;
    wire signal_20831 ;
    wire signal_20832 ;
    wire signal_20833 ;
    wire signal_20834 ;
    wire signal_20835 ;
    wire signal_20836 ;
    wire signal_20837 ;
    wire signal_20838 ;
    wire signal_20839 ;
    wire signal_20840 ;
    wire signal_20841 ;
    wire signal_20842 ;
    wire signal_20843 ;
    wire signal_20844 ;
    wire signal_20845 ;
    wire signal_20846 ;
    wire signal_20847 ;
    wire signal_20848 ;
    wire signal_20849 ;
    wire signal_20850 ;
    wire signal_20851 ;
    wire signal_20852 ;
    wire signal_20853 ;
    wire signal_20854 ;
    wire signal_20855 ;
    wire signal_20856 ;
    wire signal_20857 ;
    wire signal_20858 ;
    wire signal_20859 ;
    wire signal_20860 ;
    wire signal_20861 ;
    wire signal_20862 ;
    wire signal_20863 ;
    wire signal_20864 ;
    wire signal_20865 ;
    wire signal_20866 ;
    wire signal_20867 ;
    wire signal_20868 ;
    wire signal_20869 ;
    wire signal_20870 ;
    wire signal_20871 ;
    wire signal_20872 ;
    wire signal_20873 ;
    wire signal_20874 ;
    wire signal_20875 ;
    wire signal_20876 ;
    wire signal_20877 ;
    wire signal_20878 ;
    wire signal_20879 ;
    wire signal_20880 ;
    wire signal_20881 ;
    wire signal_20882 ;
    wire signal_20883 ;
    wire signal_20884 ;
    wire signal_20885 ;
    wire signal_20886 ;
    wire signal_20887 ;
    wire signal_20888 ;
    wire signal_20889 ;
    wire signal_20890 ;
    wire signal_20891 ;
    wire signal_20892 ;
    wire signal_20893 ;
    wire signal_20894 ;
    wire signal_20895 ;
    wire signal_20896 ;
    wire signal_20897 ;
    wire signal_20898 ;
    wire signal_20899 ;
    wire signal_20900 ;
    wire signal_20901 ;
    wire signal_20902 ;
    wire signal_20903 ;
    wire signal_20904 ;
    wire signal_20905 ;
    wire signal_20906 ;
    wire signal_20907 ;
    wire signal_20908 ;
    wire signal_20909 ;
    wire signal_20910 ;
    wire signal_20911 ;
    wire signal_20912 ;
    wire signal_20913 ;
    wire signal_20914 ;
    wire signal_20915 ;
    wire signal_20916 ;
    wire signal_20917 ;
    wire signal_20918 ;
    wire signal_20919 ;
    wire signal_20920 ;
    wire signal_20921 ;
    wire signal_20922 ;
    wire signal_20923 ;
    wire signal_20924 ;
    wire signal_20925 ;
    wire signal_20926 ;
    wire signal_20927 ;
    wire signal_20928 ;
    wire signal_20929 ;
    wire signal_20930 ;
    wire signal_20931 ;
    wire signal_20932 ;
    wire signal_20933 ;
    wire signal_20934 ;
    wire signal_20935 ;
    wire signal_20936 ;
    wire signal_20937 ;
    wire signal_20938 ;
    wire signal_20939 ;
    wire signal_20940 ;
    wire signal_20941 ;
    wire signal_20942 ;
    wire signal_20943 ;
    wire signal_20944 ;
    wire signal_20945 ;
    wire signal_20946 ;
    wire signal_20947 ;
    wire signal_20948 ;
    wire signal_20949 ;
    wire signal_20950 ;
    wire signal_20951 ;
    wire signal_20952 ;
    wire signal_20953 ;
    wire signal_20954 ;
    wire signal_20955 ;
    wire signal_20956 ;
    wire signal_20957 ;
    wire signal_20958 ;
    wire signal_20959 ;
    wire signal_20960 ;
    wire signal_20961 ;
    wire signal_20962 ;
    wire signal_20963 ;
    wire signal_20964 ;
    wire signal_20965 ;
    wire signal_20966 ;
    wire signal_20967 ;
    wire signal_20968 ;
    wire signal_20969 ;
    wire signal_20970 ;
    wire signal_20971 ;
    wire signal_20972 ;
    wire signal_20973 ;
    wire signal_20974 ;
    wire signal_20975 ;
    wire signal_20976 ;
    wire signal_20977 ;
    wire signal_20978 ;
    wire signal_20979 ;
    wire signal_20980 ;
    wire signal_20981 ;
    wire signal_20982 ;
    wire signal_20983 ;
    wire signal_20984 ;
    wire signal_20985 ;
    wire signal_20986 ;
    wire signal_20987 ;
    wire signal_20988 ;
    wire signal_20989 ;
    wire signal_20990 ;
    wire signal_20991 ;
    wire signal_20992 ;
    wire signal_20993 ;
    wire signal_20994 ;
    wire signal_20995 ;
    wire signal_20996 ;
    wire signal_20997 ;
    wire signal_20998 ;
    wire signal_20999 ;
    wire signal_21000 ;
    wire signal_21001 ;
    wire signal_21002 ;
    wire signal_21003 ;
    wire signal_21004 ;
    wire signal_21005 ;
    wire signal_21006 ;
    wire signal_21007 ;
    wire signal_21008 ;
    wire signal_21009 ;
    wire signal_21010 ;
    wire signal_21011 ;
    wire signal_21012 ;
    wire signal_21013 ;
    wire signal_21014 ;
    wire signal_21015 ;
    wire signal_21016 ;
    wire signal_21017 ;
    wire signal_21018 ;
    wire signal_21019 ;
    wire signal_21020 ;
    wire signal_21021 ;
    wire signal_21022 ;
    wire signal_21023 ;
    wire signal_21024 ;
    wire signal_21025 ;
    wire signal_21026 ;
    wire signal_21027 ;
    wire signal_21028 ;
    wire signal_21029 ;
    wire signal_21030 ;
    wire signal_21031 ;
    wire signal_21032 ;
    wire signal_21033 ;
    wire signal_21034 ;
    wire signal_21035 ;
    wire signal_21036 ;
    wire signal_21037 ;
    wire signal_21038 ;
    wire signal_21039 ;
    wire signal_21040 ;
    wire signal_21041 ;
    wire signal_21042 ;
    wire signal_21043 ;
    wire signal_21044 ;
    wire signal_21045 ;
    wire signal_21046 ;
    wire signal_21047 ;
    wire signal_21048 ;
    wire signal_21049 ;
    wire signal_21050 ;
    wire signal_21051 ;
    wire signal_21052 ;
    wire signal_21053 ;
    wire signal_21054 ;
    wire signal_21055 ;
    wire signal_21056 ;
    wire signal_21057 ;
    wire signal_21058 ;
    wire signal_21059 ;
    wire signal_21060 ;
    wire signal_21061 ;
    wire signal_21062 ;
    wire signal_21063 ;
    wire signal_21064 ;
    wire signal_21065 ;
    wire signal_21066 ;
    wire signal_21067 ;
    wire signal_21068 ;
    wire signal_21069 ;
    wire signal_21070 ;
    wire signal_21071 ;
    wire signal_21072 ;
    wire signal_21073 ;
    wire signal_21074 ;
    wire signal_21075 ;
    wire signal_21076 ;
    wire signal_21077 ;
    wire signal_21078 ;
    wire signal_21079 ;
    wire signal_21080 ;
    wire signal_21081 ;
    wire signal_21082 ;
    wire signal_21083 ;
    wire signal_21084 ;
    wire signal_21085 ;
    wire signal_21086 ;
    wire signal_21087 ;
    wire signal_21088 ;
    wire signal_21089 ;
    wire signal_21090 ;
    wire signal_21091 ;
    wire signal_21092 ;
    wire signal_21093 ;
    wire signal_21094 ;
    wire signal_21095 ;
    wire signal_21096 ;
    wire signal_21097 ;
    wire signal_21098 ;
    wire signal_21099 ;
    wire signal_21100 ;
    wire signal_21101 ;
    wire signal_21102 ;
    wire signal_21103 ;
    wire signal_21104 ;
    wire signal_21105 ;
    wire signal_21106 ;
    wire signal_21107 ;
    wire signal_21108 ;
    wire signal_21109 ;
    wire signal_21110 ;
    wire signal_21111 ;
    wire signal_21112 ;
    wire signal_21113 ;
    wire signal_21114 ;
    wire signal_21115 ;
    wire signal_21116 ;
    wire signal_21117 ;
    wire signal_21118 ;
    wire signal_21119 ;
    wire signal_21120 ;
    wire signal_21121 ;
    wire signal_21122 ;
    wire signal_21123 ;
    wire signal_21124 ;
    wire signal_21125 ;
    wire signal_21126 ;
    wire signal_21127 ;
    wire signal_21128 ;
    wire signal_21129 ;
    wire signal_21130 ;
    wire signal_21131 ;
    wire signal_21132 ;
    wire signal_21133 ;
    wire signal_21134 ;
    wire signal_21135 ;
    wire signal_21136 ;
    wire signal_21137 ;
    wire signal_21138 ;
    wire signal_21139 ;
    wire signal_21140 ;
    wire signal_21141 ;
    wire signal_21142 ;
    wire signal_21143 ;
    wire signal_21144 ;
    wire signal_21145 ;
    wire signal_21146 ;
    wire signal_21147 ;
    wire signal_21148 ;
    wire signal_21149 ;
    wire signal_21150 ;
    wire signal_21151 ;
    wire signal_21152 ;
    wire signal_21153 ;
    wire signal_21154 ;
    wire signal_21155 ;
    wire signal_21156 ;
    wire signal_21157 ;
    wire signal_21158 ;
    wire signal_21159 ;
    wire signal_21160 ;
    wire signal_21161 ;
    wire signal_21162 ;
    wire signal_21163 ;
    wire signal_21164 ;
    wire signal_21165 ;
    wire signal_21166 ;
    wire signal_21167 ;
    wire signal_21168 ;
    wire signal_21169 ;
    wire signal_21170 ;
    wire signal_21171 ;
    wire signal_21172 ;
    wire signal_21173 ;
    wire signal_21174 ;
    wire signal_21175 ;
    wire signal_21176 ;
    wire signal_21177 ;
    wire signal_21178 ;
    wire signal_21179 ;
    wire signal_21180 ;
    wire signal_21181 ;
    wire signal_21182 ;
    wire signal_21183 ;
    wire signal_21184 ;
    wire signal_21185 ;
    wire signal_21186 ;
    wire signal_21187 ;
    wire signal_21188 ;
    wire signal_21189 ;
    wire signal_21190 ;
    wire signal_21191 ;
    wire signal_21192 ;
    wire signal_21193 ;
    wire signal_21194 ;
    wire signal_21195 ;
    wire signal_21196 ;
    wire signal_21197 ;
    wire signal_21198 ;
    wire signal_21199 ;
    wire signal_21200 ;
    wire signal_21201 ;
    wire signal_21202 ;
    wire signal_21203 ;
    wire signal_21204 ;
    wire signal_21205 ;
    wire signal_21206 ;
    wire signal_21207 ;
    wire signal_21208 ;
    wire signal_21209 ;
    wire signal_21210 ;
    wire signal_21211 ;
    wire signal_21212 ;
    wire signal_21213 ;
    wire signal_21214 ;
    wire signal_21215 ;
    wire signal_21216 ;
    wire signal_21217 ;
    wire signal_21218 ;
    wire signal_21219 ;
    wire signal_21220 ;
    wire signal_21221 ;
    wire signal_21222 ;
    wire signal_21223 ;
    wire signal_21224 ;
    wire signal_21225 ;
    wire signal_21226 ;
    wire signal_21227 ;
    wire signal_21228 ;
    wire signal_21229 ;
    wire signal_21230 ;
    wire signal_21231 ;
    wire signal_21232 ;
    wire signal_21233 ;
    wire signal_21234 ;
    wire signal_21235 ;
    wire signal_21236 ;
    wire signal_21237 ;
    wire signal_21238 ;
    wire signal_21239 ;
    wire signal_21240 ;
    wire signal_21241 ;
    wire signal_21242 ;
    wire signal_21243 ;
    wire signal_21244 ;
    wire signal_21245 ;
    wire signal_21246 ;
    wire signal_21247 ;
    wire signal_21248 ;
    wire signal_21249 ;
    wire signal_21250 ;
    wire signal_21251 ;
    wire signal_21252 ;
    wire signal_21253 ;
    wire signal_21254 ;
    wire signal_21255 ;
    wire signal_21256 ;
    wire signal_21257 ;
    wire signal_21258 ;
    wire signal_21259 ;
    wire signal_21260 ;
    wire signal_21261 ;
    wire signal_21262 ;
    wire signal_21263 ;
    wire signal_21264 ;
    wire signal_21265 ;
    wire signal_21266 ;
    wire signal_21267 ;
    wire signal_21268 ;
    wire signal_21269 ;
    wire signal_21270 ;
    wire signal_21271 ;
    wire signal_21272 ;
    wire signal_21273 ;
    wire signal_21274 ;
    wire signal_21275 ;
    wire signal_21276 ;
    wire signal_21277 ;
    wire signal_21278 ;
    wire signal_21279 ;
    wire signal_21280 ;
    wire signal_21281 ;
    wire signal_21282 ;
    wire signal_21283 ;
    wire signal_21284 ;
    wire signal_21285 ;
    wire signal_21286 ;
    wire signal_21287 ;
    wire signal_21288 ;
    wire signal_21289 ;
    wire signal_21290 ;
    wire signal_21291 ;
    wire signal_21292 ;
    wire signal_21293 ;
    wire signal_21294 ;
    wire signal_21295 ;
    wire signal_21296 ;
    wire signal_21297 ;
    wire signal_21298 ;
    wire signal_21299 ;
    wire signal_21300 ;
    wire signal_21301 ;
    wire signal_21302 ;
    wire signal_21303 ;
    wire signal_21304 ;
    wire signal_21305 ;
    wire signal_21306 ;
    wire signal_21307 ;
    wire signal_21308 ;
    wire signal_21309 ;
    wire signal_21310 ;
    wire signal_21311 ;
    wire signal_21312 ;
    wire signal_21313 ;
    wire signal_21314 ;
    wire signal_21315 ;
    wire signal_21316 ;
    wire signal_21317 ;
    wire signal_21318 ;
    wire signal_21319 ;
    wire signal_21320 ;
    wire signal_21321 ;
    wire signal_21322 ;
    wire signal_21323 ;
    wire signal_21324 ;
    wire signal_21325 ;
    wire signal_21326 ;
    wire signal_21327 ;
    wire signal_21328 ;
    wire signal_21329 ;
    wire signal_21330 ;
    wire signal_21331 ;
    wire signal_21332 ;
    wire signal_21333 ;
    wire signal_21334 ;
    wire signal_21335 ;
    wire signal_21336 ;
    wire signal_21337 ;
    wire signal_21338 ;
    wire signal_21339 ;
    wire signal_21340 ;
    wire signal_21341 ;
    wire signal_21342 ;
    wire signal_21343 ;
    wire signal_21344 ;
    wire signal_21345 ;
    wire signal_21346 ;
    wire signal_21347 ;
    wire signal_21348 ;
    wire signal_21349 ;
    wire signal_21350 ;
    wire signal_21351 ;
    wire signal_21352 ;
    wire signal_21353 ;
    wire signal_21354 ;
    wire signal_21355 ;
    wire signal_21356 ;
    wire signal_21357 ;
    wire signal_21358 ;
    wire signal_21359 ;
    wire signal_21360 ;
    wire signal_21361 ;
    wire signal_21362 ;
    wire signal_21363 ;
    wire signal_21364 ;
    wire signal_21365 ;
    wire signal_21366 ;
    wire signal_21367 ;
    wire signal_21368 ;
    wire signal_21369 ;
    wire signal_21370 ;
    wire signal_21371 ;
    wire signal_21372 ;
    wire signal_21373 ;
    wire signal_21374 ;
    wire signal_21375 ;
    wire signal_21376 ;
    wire signal_21377 ;
    wire signal_21378 ;
    wire signal_21379 ;
    wire signal_21380 ;
    wire signal_21381 ;
    wire signal_21382 ;
    wire signal_21383 ;
    wire signal_21384 ;
    wire signal_21385 ;
    wire signal_21386 ;
    wire signal_21387 ;
    wire signal_21388 ;
    wire signal_21389 ;
    wire signal_21390 ;
    wire signal_21391 ;
    wire signal_21392 ;
    wire signal_21393 ;
    wire signal_21394 ;
    wire signal_21395 ;
    wire signal_21396 ;
    wire signal_21397 ;
    wire signal_21398 ;
    wire signal_21399 ;
    wire signal_21400 ;
    wire signal_21401 ;
    wire signal_21402 ;
    wire signal_21403 ;
    wire signal_21404 ;
    wire signal_21405 ;
    wire signal_21406 ;
    wire signal_21407 ;
    wire signal_21408 ;
    wire signal_21409 ;
    wire signal_21410 ;
    wire signal_21411 ;
    wire signal_21412 ;
    wire signal_21413 ;
    wire signal_21414 ;
    wire signal_21415 ;
    wire signal_21416 ;
    wire signal_21417 ;
    wire signal_21418 ;
    wire signal_21419 ;
    wire signal_21420 ;
    wire signal_21421 ;
    wire signal_21422 ;
    wire signal_21423 ;
    wire signal_21424 ;
    wire signal_21425 ;
    wire signal_21426 ;
    wire signal_21427 ;
    wire signal_21428 ;
    wire signal_21429 ;
    wire signal_21430 ;
    wire signal_21431 ;
    wire signal_21432 ;
    wire signal_21433 ;
    wire signal_21434 ;
    wire signal_21435 ;
    wire signal_21436 ;
    wire signal_21437 ;
    wire signal_21438 ;
    wire signal_21439 ;
    wire signal_21440 ;
    wire signal_21441 ;
    wire signal_21442 ;
    wire signal_21443 ;
    wire signal_21444 ;
    wire signal_21445 ;
    wire signal_21446 ;
    wire signal_21447 ;
    wire signal_21448 ;
    wire signal_21449 ;
    wire signal_21450 ;
    wire signal_21451 ;
    wire signal_21452 ;
    wire signal_21453 ;
    wire signal_21454 ;
    wire signal_21455 ;
    wire signal_21456 ;
    wire signal_21457 ;
    wire signal_21458 ;
    wire signal_21459 ;
    wire signal_21460 ;
    wire signal_21461 ;
    wire signal_21462 ;
    wire signal_21463 ;
    wire signal_21464 ;
    wire signal_21465 ;
    wire signal_21466 ;
    wire signal_21467 ;
    wire signal_21468 ;
    wire signal_21469 ;
    wire signal_21470 ;
    wire signal_21471 ;
    wire signal_21472 ;
    wire signal_21473 ;
    wire signal_21474 ;
    wire signal_21475 ;
    wire signal_21476 ;
    wire signal_21477 ;
    wire signal_21478 ;
    wire signal_21479 ;
    wire signal_21480 ;
    wire signal_21481 ;
    wire signal_21482 ;
    wire signal_21483 ;
    wire signal_21484 ;
    wire signal_21485 ;
    wire signal_21486 ;
    wire signal_21487 ;
    wire signal_21488 ;
    wire signal_21489 ;
    wire signal_21490 ;
    wire signal_21491 ;
    wire signal_21492 ;
    wire signal_21493 ;
    wire signal_21494 ;
    wire signal_21495 ;
    wire signal_21496 ;
    wire signal_21497 ;
    wire signal_21498 ;
    wire signal_21499 ;
    wire signal_21500 ;
    wire signal_21501 ;
    wire signal_21502 ;
    wire signal_21503 ;
    wire signal_21504 ;
    wire signal_21505 ;
    wire signal_21506 ;
    wire signal_21507 ;
    wire signal_21508 ;
    wire signal_21509 ;
    wire signal_21510 ;
    wire signal_21511 ;
    wire signal_21512 ;
    wire signal_21513 ;
    wire signal_21514 ;
    wire signal_21515 ;
    wire signal_21516 ;
    wire signal_21517 ;
    wire signal_21518 ;
    wire signal_21519 ;
    wire signal_21520 ;
    wire signal_21521 ;
    wire signal_21522 ;
    wire signal_21523 ;
    wire signal_21524 ;
    wire signal_21525 ;
    wire signal_21526 ;
    wire signal_21527 ;
    wire signal_21528 ;
    wire signal_21529 ;
    wire signal_21530 ;
    wire signal_21531 ;
    wire signal_21532 ;
    wire signal_21533 ;
    wire signal_21534 ;
    wire signal_21535 ;
    wire signal_21536 ;
    wire signal_21537 ;
    wire signal_21538 ;
    wire signal_21539 ;
    wire signal_21540 ;
    wire signal_21541 ;
    wire signal_21542 ;
    wire signal_21543 ;
    wire signal_21544 ;
    wire signal_21545 ;
    wire signal_21546 ;
    wire signal_21547 ;
    wire signal_21548 ;
    wire signal_21549 ;
    wire signal_21550 ;
    wire signal_21551 ;
    wire signal_21552 ;
    wire signal_21553 ;
    wire signal_21554 ;
    wire signal_21555 ;
    wire signal_21556 ;
    wire signal_21557 ;
    wire signal_21558 ;
    wire signal_21559 ;
    wire signal_21560 ;
    wire signal_21561 ;
    wire signal_21562 ;
    wire signal_21563 ;
    wire signal_21564 ;
    wire signal_21565 ;
    wire signal_21566 ;
    wire signal_21567 ;
    wire signal_21568 ;
    wire signal_21569 ;
    wire signal_21570 ;
    wire signal_21571 ;
    wire signal_21572 ;
    wire signal_21573 ;
    wire signal_21574 ;
    wire signal_21575 ;
    wire signal_21576 ;
    wire signal_21577 ;
    wire signal_21578 ;
    wire signal_21579 ;
    wire signal_21580 ;
    wire signal_21581 ;
    wire signal_21582 ;
    wire signal_21583 ;
    wire signal_21584 ;
    wire signal_21585 ;
    wire signal_21586 ;
    wire signal_21587 ;
    wire signal_21588 ;
    wire signal_21589 ;
    wire signal_21590 ;
    wire signal_21591 ;
    wire signal_21592 ;
    wire signal_21593 ;
    wire signal_21594 ;
    wire signal_21595 ;
    wire signal_21596 ;
    wire signal_21597 ;
    wire signal_21598 ;
    wire signal_21599 ;
    wire signal_21600 ;
    wire signal_21601 ;
    wire signal_21602 ;
    wire signal_21603 ;
    wire signal_21604 ;
    wire signal_21605 ;
    wire signal_21606 ;
    wire signal_21607 ;
    wire signal_21608 ;
    wire signal_21609 ;
    wire signal_21610 ;
    wire signal_21611 ;
    wire signal_21612 ;
    wire signal_21613 ;
    wire signal_21614 ;
    wire signal_21615 ;
    wire signal_21616 ;
    wire signal_21617 ;
    wire signal_21618 ;
    wire signal_21619 ;
    wire signal_21620 ;
    wire signal_21621 ;
    wire signal_21622 ;
    wire signal_21623 ;
    wire signal_21624 ;
    wire signal_21625 ;
    wire signal_21626 ;
    wire signal_21627 ;
    wire signal_21628 ;
    wire signal_21629 ;
    wire signal_21630 ;
    wire signal_21631 ;
    wire signal_21632 ;
    wire signal_21633 ;
    wire signal_21634 ;
    wire signal_21635 ;
    wire signal_21636 ;
    wire signal_21637 ;
    wire signal_21638 ;
    wire signal_21639 ;
    wire signal_21640 ;
    wire signal_21641 ;
    wire signal_21642 ;
    wire signal_21643 ;
    wire signal_21644 ;
    wire signal_21645 ;
    wire signal_21646 ;
    wire signal_21647 ;
    wire signal_21648 ;
    wire signal_21649 ;
    wire signal_21650 ;
    wire signal_21651 ;
    wire signal_21652 ;
    wire signal_21653 ;
    wire signal_21654 ;
    wire signal_21655 ;
    wire signal_21656 ;
    wire signal_21657 ;
    wire signal_21658 ;
    wire signal_21659 ;
    wire signal_21660 ;
    wire signal_21661 ;
    wire signal_21662 ;
    wire signal_21663 ;
    wire signal_21664 ;
    wire signal_21665 ;
    wire signal_21666 ;
    wire signal_21667 ;
    wire signal_21668 ;
    wire signal_21669 ;
    wire signal_21670 ;
    wire signal_21671 ;
    wire signal_21672 ;
    wire signal_21673 ;
    wire signal_21674 ;
    wire signal_21675 ;
    wire signal_21676 ;
    wire signal_21677 ;
    wire signal_21678 ;
    wire signal_21679 ;
    wire signal_21680 ;
    wire signal_21681 ;
    wire signal_21682 ;
    wire signal_21683 ;
    wire signal_21684 ;
    wire signal_21685 ;
    wire signal_21686 ;
    wire signal_21687 ;
    wire signal_21688 ;
    wire signal_21689 ;
    wire signal_21690 ;
    wire signal_21691 ;
    wire signal_21692 ;
    wire signal_21693 ;
    wire signal_21694 ;
    wire signal_21695 ;
    wire signal_21696 ;
    wire signal_21697 ;
    wire signal_21698 ;
    wire signal_21699 ;
    wire signal_21700 ;
    wire signal_21701 ;
    wire signal_21702 ;
    wire signal_21703 ;
    wire signal_21704 ;
    wire signal_21705 ;
    wire signal_21706 ;
    wire signal_21707 ;
    wire signal_21708 ;
    wire signal_21709 ;
    wire signal_21710 ;
    wire signal_21711 ;
    wire signal_21712 ;
    wire signal_21713 ;
    wire signal_21714 ;
    wire signal_21715 ;
    wire signal_21716 ;
    wire signal_21717 ;
    wire signal_21718 ;
    wire signal_21719 ;
    wire signal_21720 ;
    wire signal_21721 ;
    wire signal_21722 ;
    wire signal_21723 ;
    wire signal_21724 ;
    wire signal_21725 ;
    wire signal_21726 ;
    wire signal_21727 ;
    wire signal_21728 ;
    wire signal_21729 ;
    wire signal_21730 ;
    wire signal_21731 ;
    wire signal_21732 ;
    wire signal_21733 ;
    wire signal_21734 ;
    wire signal_21735 ;
    wire signal_21736 ;
    wire signal_21737 ;
    wire signal_21738 ;
    wire signal_21739 ;
    wire signal_21740 ;
    wire signal_21741 ;
    wire signal_21742 ;
    wire signal_21743 ;
    wire signal_21744 ;
    wire signal_21745 ;
    wire signal_21746 ;
    wire signal_21747 ;
    wire signal_21748 ;
    wire signal_21749 ;
    wire signal_21750 ;
    wire signal_21751 ;
    wire signal_21752 ;
    wire signal_21753 ;
    wire signal_21754 ;
    wire signal_21755 ;
    wire signal_21756 ;
    wire signal_21757 ;
    wire signal_21758 ;
    wire signal_21759 ;
    wire signal_21760 ;
    wire signal_21761 ;
    wire signal_21762 ;
    wire signal_21763 ;
    wire signal_21764 ;
    wire signal_21765 ;
    wire signal_21766 ;
    wire signal_21767 ;
    wire signal_21768 ;
    wire signal_21769 ;
    wire signal_21770 ;
    wire signal_21771 ;
    wire signal_21772 ;
    wire signal_21773 ;
    wire signal_21774 ;
    wire signal_21775 ;
    wire signal_21776 ;
    wire signal_21777 ;
    wire signal_21778 ;
    wire signal_21779 ;
    wire signal_21780 ;
    wire signal_21781 ;
    wire signal_21782 ;
    wire signal_21783 ;
    wire signal_21784 ;
    wire signal_21785 ;
    wire signal_21786 ;
    wire signal_21787 ;
    wire signal_21788 ;
    wire signal_21789 ;
    wire signal_21790 ;
    wire signal_21791 ;
    wire signal_21792 ;
    wire signal_21793 ;
    wire signal_21794 ;
    wire signal_21795 ;
    wire signal_21796 ;
    wire signal_21797 ;
    wire signal_21798 ;
    wire signal_21799 ;
    wire signal_21800 ;
    wire signal_21801 ;
    wire signal_21802 ;
    wire signal_21803 ;
    wire signal_21804 ;
    wire signal_21805 ;
    wire signal_21806 ;
    wire signal_21807 ;
    wire signal_21808 ;
    wire signal_21809 ;
    wire signal_21810 ;
    wire signal_21811 ;
    wire signal_21812 ;
    wire signal_21813 ;
    wire signal_21814 ;
    wire signal_21815 ;
    wire signal_21816 ;
    wire signal_21817 ;
    wire signal_21818 ;
    wire signal_21819 ;
    wire signal_21820 ;
    wire signal_21821 ;
    wire signal_21822 ;
    wire signal_21823 ;
    wire signal_21824 ;
    wire signal_21825 ;
    wire signal_21826 ;
    wire signal_21827 ;
    wire signal_21828 ;
    wire signal_21829 ;
    wire signal_21830 ;
    wire signal_21831 ;
    wire signal_21832 ;
    wire signal_21833 ;
    wire signal_21834 ;
    wire signal_21835 ;
    wire signal_21836 ;
    wire signal_21837 ;
    wire signal_21838 ;
    wire signal_21839 ;
    wire signal_21840 ;
    wire signal_21841 ;
    wire signal_21842 ;
    wire signal_21843 ;
    wire signal_21844 ;
    wire signal_21845 ;
    wire signal_21846 ;
    wire signal_21847 ;
    wire signal_21848 ;
    wire signal_21849 ;
    wire signal_21850 ;
    wire signal_21851 ;
    wire signal_21852 ;
    wire signal_21853 ;
    wire signal_21854 ;
    wire signal_21855 ;
    wire signal_21856 ;
    wire signal_21857 ;
    wire signal_21858 ;
    wire signal_21859 ;
    wire signal_21860 ;
    wire signal_21861 ;
    wire signal_21862 ;
    wire signal_21863 ;
    wire signal_21864 ;
    wire signal_21865 ;
    wire signal_21866 ;
    wire signal_21867 ;
    wire signal_21868 ;
    wire signal_21869 ;
    wire signal_21870 ;
    wire signal_21871 ;
    wire signal_21872 ;
    wire signal_21873 ;
    wire signal_21874 ;
    wire signal_21875 ;
    wire signal_21876 ;
    wire signal_21877 ;
    wire signal_21878 ;
    wire signal_21879 ;
    wire signal_21880 ;
    wire signal_21881 ;
    wire signal_21882 ;
    wire signal_21883 ;
    wire signal_21884 ;
    wire signal_21885 ;
    wire signal_21886 ;
    wire signal_21887 ;
    wire signal_21888 ;
    wire signal_21889 ;
    wire signal_21890 ;
    wire signal_21891 ;
    wire signal_21892 ;
    wire signal_21893 ;
    wire signal_21894 ;
    wire signal_21895 ;
    wire signal_21896 ;
    wire signal_21897 ;
    wire signal_21898 ;
    wire signal_21899 ;
    wire signal_21900 ;
    wire signal_21901 ;
    wire signal_21902 ;
    wire signal_21903 ;
    wire signal_21904 ;
    wire signal_21905 ;
    wire signal_21906 ;
    wire signal_21907 ;
    wire signal_21908 ;
    wire signal_21909 ;
    wire signal_21910 ;
    wire signal_21911 ;
    wire signal_21912 ;
    wire signal_21913 ;
    wire signal_21914 ;
    wire signal_21915 ;
    wire signal_21916 ;
    wire signal_21917 ;
    wire signal_21918 ;
    wire signal_21919 ;
    wire signal_21920 ;
    wire signal_21921 ;
    wire signal_21922 ;
    wire signal_21923 ;
    wire signal_21924 ;
    wire signal_21925 ;
    wire signal_21926 ;
    wire signal_21927 ;
    wire signal_21928 ;
    wire signal_21929 ;
    wire signal_21930 ;
    wire signal_21931 ;
    wire signal_21932 ;
    wire signal_21933 ;
    wire signal_21934 ;
    wire signal_21935 ;
    wire signal_21936 ;
    wire signal_21937 ;
    wire signal_21938 ;
    wire signal_21939 ;
    wire signal_21940 ;
    wire signal_21941 ;
    wire signal_21942 ;
    wire signal_21943 ;
    wire signal_21944 ;
    wire signal_21945 ;
    wire signal_21946 ;
    wire signal_21947 ;
    wire signal_21948 ;
    wire signal_21949 ;
    wire signal_21950 ;
    wire signal_21951 ;
    wire signal_21952 ;
    wire signal_21953 ;
    wire signal_21954 ;
    wire signal_21955 ;
    wire signal_21956 ;
    wire signal_21957 ;
    wire signal_21958 ;
    wire signal_21959 ;
    wire signal_21960 ;
    wire signal_21961 ;
    wire signal_21962 ;
    wire signal_21963 ;
    wire signal_21964 ;
    wire signal_21965 ;
    wire signal_21966 ;
    wire signal_21967 ;
    wire signal_21968 ;
    wire signal_21969 ;
    wire signal_21970 ;
    wire signal_21971 ;
    wire signal_21972 ;
    wire signal_21973 ;
    wire signal_21974 ;
    wire signal_21975 ;
    wire signal_21976 ;
    wire signal_21977 ;
    wire signal_21978 ;
    wire signal_21979 ;
    wire signal_21980 ;
    wire signal_21981 ;
    wire signal_21982 ;
    wire signal_21983 ;
    wire signal_21984 ;
    wire signal_21985 ;
    wire signal_21986 ;
    wire signal_21987 ;
    wire signal_21988 ;
    wire signal_21989 ;
    wire signal_21990 ;
    wire signal_21991 ;
    wire signal_21992 ;
    wire signal_21993 ;
    wire signal_21994 ;
    wire signal_21995 ;
    wire signal_21996 ;
    wire signal_21997 ;
    wire signal_21998 ;
    wire signal_21999 ;
    wire signal_22000 ;
    wire signal_22001 ;
    wire signal_22002 ;
    wire signal_22003 ;
    wire signal_22004 ;
    wire signal_22005 ;
    wire signal_22006 ;
    wire signal_22007 ;
    wire signal_22008 ;
    wire signal_22009 ;
    wire signal_22010 ;
    wire signal_22011 ;
    wire signal_22012 ;
    wire signal_22013 ;
    wire signal_22014 ;
    wire signal_22015 ;
    wire signal_22016 ;
    wire signal_22017 ;
    wire signal_22018 ;
    wire signal_22019 ;
    wire signal_22020 ;
    wire signal_22021 ;
    wire signal_22022 ;
    wire signal_22023 ;
    wire signal_22024 ;
    wire signal_22025 ;
    wire signal_22026 ;
    wire signal_22027 ;
    wire signal_22028 ;
    wire signal_22029 ;
    wire signal_22030 ;
    wire signal_22031 ;
    wire signal_22032 ;
    wire signal_22033 ;
    wire signal_22034 ;
    wire signal_22035 ;
    wire signal_22036 ;
    wire signal_22037 ;
    wire signal_22038 ;
    wire signal_22039 ;
    wire signal_22040 ;
    wire signal_22041 ;
    wire signal_22042 ;
    wire signal_22043 ;
    wire signal_22044 ;
    wire signal_22045 ;
    wire signal_22046 ;
    wire signal_22047 ;
    wire signal_22048 ;
    wire signal_22049 ;
    wire signal_22050 ;
    wire signal_22051 ;
    wire signal_22052 ;
    wire signal_22053 ;
    wire signal_22054 ;
    wire signal_22055 ;
    wire signal_22056 ;
    wire signal_22057 ;
    wire signal_22058 ;
    wire signal_22059 ;
    wire signal_22060 ;
    wire signal_22061 ;
    wire signal_22062 ;
    wire signal_22063 ;
    wire signal_22064 ;
    wire signal_22065 ;
    wire signal_22066 ;
    wire signal_22067 ;
    wire signal_22068 ;
    wire signal_22069 ;
    wire signal_22070 ;
    wire signal_22071 ;
    wire signal_22072 ;
    wire signal_22073 ;
    wire signal_22074 ;
    wire signal_22075 ;
    wire signal_22076 ;
    wire signal_22077 ;
    wire signal_22078 ;
    wire signal_22079 ;
    wire signal_22080 ;
    wire signal_22081 ;
    wire signal_22082 ;
    wire signal_22083 ;
    wire signal_22084 ;
    wire signal_22085 ;
    wire signal_22086 ;
    wire signal_22087 ;
    wire signal_22088 ;
    wire signal_22089 ;
    wire signal_22090 ;
    wire signal_22091 ;
    wire signal_22092 ;
    wire signal_22093 ;
    wire signal_22094 ;
    wire signal_22095 ;
    wire signal_22096 ;
    wire signal_22097 ;
    wire signal_22098 ;
    wire signal_22099 ;
    wire signal_22100 ;
    wire signal_22101 ;
    wire signal_22102 ;
    wire signal_22103 ;
    wire signal_22104 ;
    wire signal_22105 ;
    wire signal_22106 ;
    wire signal_22107 ;
    wire signal_22108 ;
    wire signal_22109 ;
    wire signal_22110 ;
    wire signal_22111 ;
    wire signal_22112 ;
    wire signal_22113 ;
    wire signal_22114 ;
    wire signal_22115 ;
    wire signal_22116 ;
    wire signal_22117 ;
    wire signal_22118 ;
    wire signal_22119 ;
    wire signal_22120 ;
    wire signal_22121 ;
    wire signal_22122 ;
    wire signal_22123 ;
    wire signal_22124 ;
    wire signal_22125 ;
    wire signal_22126 ;
    wire signal_22127 ;
    wire signal_22128 ;
    wire signal_22129 ;
    wire signal_22130 ;
    wire signal_22131 ;
    wire signal_22132 ;
    wire signal_22133 ;
    wire signal_22134 ;
    wire signal_22135 ;
    wire signal_22136 ;
    wire signal_22137 ;
    wire signal_22138 ;
    wire signal_22139 ;
    wire signal_22140 ;
    wire signal_22141 ;
    wire signal_22142 ;
    wire signal_22143 ;
    wire signal_22144 ;
    wire signal_22145 ;
    wire signal_22146 ;
    wire signal_22147 ;
    wire signal_22148 ;
    wire signal_22149 ;
    wire signal_22150 ;
    wire signal_22151 ;
    wire signal_22152 ;
    wire signal_22153 ;
    wire signal_22154 ;
    wire signal_22155 ;
    wire signal_22156 ;
    wire signal_22157 ;
    wire signal_22158 ;
    wire signal_22159 ;
    wire signal_22160 ;
    wire signal_22161 ;
    wire signal_22162 ;
    wire signal_22163 ;
    wire signal_22164 ;
    wire signal_22165 ;
    wire signal_22166 ;
    wire signal_22167 ;
    wire signal_22168 ;
    wire signal_22169 ;
    wire signal_22170 ;
    wire signal_22171 ;
    wire signal_22172 ;
    wire signal_22173 ;
    wire signal_22174 ;
    wire signal_22175 ;
    wire signal_22176 ;
    wire signal_22177 ;
    wire signal_22178 ;
    wire signal_22179 ;
    wire signal_22180 ;
    wire signal_22181 ;
    wire signal_22182 ;
    wire signal_22183 ;
    wire signal_22184 ;
    wire signal_22185 ;
    wire signal_22186 ;
    wire signal_22187 ;
    wire signal_22188 ;
    wire signal_22189 ;
    wire signal_22190 ;
    wire signal_22191 ;
    wire signal_22192 ;
    wire signal_22193 ;
    wire signal_22194 ;
    wire signal_22195 ;
    wire signal_22196 ;
    wire signal_22197 ;
    wire signal_22198 ;
    wire signal_22199 ;
    wire signal_22200 ;
    wire signal_22201 ;
    wire signal_22202 ;
    wire signal_22203 ;
    wire signal_22204 ;
    wire signal_22205 ;
    wire signal_22206 ;
    wire signal_22207 ;
    wire signal_22208 ;
    wire signal_22209 ;
    wire signal_22210 ;
    wire signal_22211 ;
    wire signal_22212 ;
    wire signal_22213 ;
    wire signal_22214 ;
    wire signal_22215 ;
    wire signal_22216 ;
    wire signal_22217 ;
    wire signal_22218 ;
    wire signal_22219 ;
    wire signal_22220 ;
    wire signal_22221 ;
    wire signal_22222 ;
    wire signal_22223 ;
    wire signal_22224 ;
    wire signal_22225 ;
    wire signal_22226 ;
    wire signal_22227 ;
    wire signal_22228 ;
    wire signal_22229 ;
    wire signal_22230 ;
    wire signal_22231 ;
    wire signal_22232 ;
    wire signal_22233 ;
    wire signal_22234 ;
    wire signal_22235 ;
    wire signal_22236 ;
    wire signal_22237 ;
    wire signal_22238 ;
    wire signal_22239 ;
    wire signal_22240 ;
    wire signal_22241 ;
    wire signal_22242 ;
    wire signal_22243 ;
    wire signal_22244 ;
    wire signal_22245 ;
    wire signal_22246 ;
    wire signal_22247 ;
    wire signal_22248 ;
    wire signal_22249 ;
    wire signal_22250 ;
    wire signal_22251 ;
    wire signal_22252 ;
    wire signal_22253 ;
    wire signal_22254 ;
    wire signal_22255 ;
    wire signal_22256 ;
    wire signal_22257 ;
    wire signal_22258 ;
    wire signal_22259 ;
    wire signal_22260 ;
    wire signal_22261 ;
    wire signal_22262 ;
    wire signal_22263 ;
    wire signal_22264 ;
    wire signal_22265 ;
    wire signal_22266 ;
    wire signal_22267 ;
    wire signal_22268 ;
    wire signal_22269 ;
    wire signal_22270 ;
    wire signal_22271 ;
    wire signal_22272 ;
    wire signal_22273 ;
    wire signal_22274 ;
    wire signal_22275 ;
    wire signal_22276 ;
    wire signal_22277 ;
    wire signal_22278 ;
    wire signal_22279 ;
    wire signal_22280 ;
    wire signal_22281 ;
    wire signal_22282 ;
    wire signal_22283 ;
    wire signal_22284 ;
    wire signal_22285 ;
    wire signal_22286 ;
    wire signal_22287 ;
    wire signal_22288 ;
    wire signal_22289 ;
    wire signal_22290 ;
    wire signal_22291 ;
    wire signal_22292 ;
    wire signal_22293 ;
    wire signal_22294 ;
    wire signal_22295 ;
    wire signal_22296 ;
    wire signal_22297 ;
    wire signal_22298 ;
    wire signal_22299 ;
    wire signal_22300 ;
    wire signal_22301 ;
    wire signal_22302 ;
    wire signal_22303 ;
    wire signal_22304 ;
    wire signal_22305 ;
    wire signal_22306 ;
    wire signal_22307 ;
    wire signal_22308 ;
    wire signal_22309 ;
    wire signal_22310 ;
    wire signal_22311 ;
    wire signal_22312 ;
    wire signal_22313 ;
    wire signal_22314 ;
    wire signal_22315 ;
    wire signal_22316 ;
    wire signal_22317 ;
    wire signal_22318 ;
    wire signal_22319 ;
    wire signal_22320 ;
    wire signal_22321 ;
    wire signal_22322 ;
    wire signal_22323 ;
    wire signal_22324 ;
    wire signal_22325 ;
    wire signal_22326 ;
    wire signal_22327 ;
    wire signal_22328 ;
    wire signal_22329 ;
    wire signal_22330 ;
    wire signal_22331 ;
    wire signal_22332 ;
    wire signal_22333 ;
    wire signal_22334 ;
    wire signal_22335 ;
    wire signal_22336 ;
    wire signal_22337 ;
    wire signal_22338 ;
    wire signal_22339 ;
    wire signal_22340 ;
    wire signal_22341 ;
    wire signal_22342 ;
    wire signal_22343 ;
    wire signal_22344 ;
    wire signal_22345 ;
    wire signal_22346 ;
    wire signal_22347 ;
    wire signal_22348 ;
    wire signal_22349 ;
    wire signal_22350 ;
    wire signal_22351 ;
    wire signal_22352 ;
    wire signal_22353 ;
    wire signal_22354 ;
    wire signal_22355 ;
    wire signal_22356 ;
    wire signal_22357 ;
    wire signal_22358 ;
    wire signal_22359 ;
    wire signal_22360 ;
    wire signal_22361 ;
    wire signal_22362 ;
    wire signal_22363 ;
    wire signal_22364 ;
    wire signal_22365 ;
    wire signal_22366 ;
    wire signal_22367 ;
    wire signal_22368 ;
    wire signal_22369 ;
    wire signal_22370 ;
    wire signal_22371 ;
    wire signal_22372 ;
    wire signal_22373 ;
    wire signal_22374 ;
    wire signal_22375 ;
    wire signal_22376 ;
    wire signal_22377 ;
    wire signal_22378 ;
    wire signal_22379 ;
    wire signal_22380 ;
    wire signal_22381 ;
    wire signal_22382 ;
    wire signal_22383 ;
    wire signal_22384 ;
    wire signal_22385 ;
    wire signal_22386 ;
    wire signal_22387 ;
    wire signal_22388 ;
    wire signal_22389 ;
    wire signal_22390 ;
    wire signal_22391 ;
    wire signal_22392 ;
    wire signal_22393 ;
    wire signal_22394 ;
    wire signal_22395 ;
    wire signal_22396 ;
    wire signal_22397 ;
    wire signal_22398 ;
    wire signal_22399 ;
    wire signal_22400 ;
    wire signal_22401 ;
    wire signal_22402 ;
    wire signal_22403 ;
    wire signal_22404 ;
    wire signal_22405 ;
    wire signal_22406 ;
    wire signal_22407 ;
    wire signal_22408 ;
    wire signal_22409 ;
    wire signal_22410 ;
    wire signal_22411 ;
    wire signal_22412 ;
    wire signal_22413 ;
    wire signal_22414 ;
    wire signal_22415 ;
    wire signal_22416 ;
    wire signal_22417 ;
    wire signal_22418 ;
    wire signal_22419 ;
    wire signal_22420 ;
    wire signal_22421 ;
    wire signal_22422 ;
    wire signal_22423 ;
    wire signal_22424 ;
    wire signal_22425 ;
    wire signal_22426 ;
    wire signal_22427 ;
    wire signal_22428 ;
    wire signal_22429 ;
    wire signal_22430 ;
    wire signal_22431 ;
    wire signal_22432 ;
    wire signal_22433 ;
    wire signal_22434 ;
    wire signal_22435 ;
    wire signal_22436 ;
    wire signal_22437 ;
    wire signal_22438 ;
    wire signal_22439 ;
    wire signal_22440 ;
    wire signal_22441 ;
    wire signal_22442 ;
    wire signal_22443 ;
    wire signal_22444 ;
    wire signal_22445 ;
    wire signal_22446 ;
    wire signal_22447 ;
    wire signal_22448 ;
    wire signal_22449 ;
    wire signal_22450 ;
    wire signal_22451 ;
    wire signal_22452 ;
    wire signal_22453 ;
    wire signal_22454 ;
    wire signal_22455 ;
    wire signal_22456 ;
    wire signal_22457 ;
    wire signal_22458 ;
    wire signal_22459 ;
    wire signal_22460 ;
    wire signal_22461 ;
    wire signal_22462 ;
    wire signal_22463 ;
    wire signal_22464 ;
    wire signal_22465 ;
    wire signal_22466 ;
    wire signal_22467 ;
    wire signal_22468 ;
    wire signal_22469 ;
    wire signal_22470 ;
    wire signal_22471 ;
    wire signal_22472 ;
    wire signal_22473 ;
    wire signal_22474 ;
    wire signal_22475 ;
    wire signal_22476 ;
    wire signal_22477 ;
    wire signal_22478 ;
    wire signal_22479 ;
    wire signal_22480 ;
    wire signal_22481 ;
    wire signal_22482 ;
    wire signal_22483 ;
    wire signal_22484 ;
    wire signal_22485 ;
    wire signal_22486 ;
    wire signal_22487 ;
    wire signal_22488 ;
    wire signal_22489 ;
    wire signal_22490 ;
    wire signal_22491 ;
    wire signal_22492 ;
    wire signal_22493 ;
    wire signal_22494 ;
    wire signal_22495 ;
    wire signal_22496 ;
    wire signal_22497 ;
    wire signal_22498 ;
    wire signal_22499 ;
    wire signal_22500 ;
    wire signal_22501 ;
    wire signal_22502 ;
    wire signal_22503 ;
    wire signal_22504 ;
    wire signal_22505 ;
    wire signal_22506 ;
    wire signal_22507 ;
    wire signal_22508 ;
    wire signal_22509 ;
    wire signal_22510 ;
    wire signal_22511 ;
    wire signal_22512 ;
    wire signal_22513 ;
    wire signal_22514 ;
    wire signal_22515 ;
    wire signal_22516 ;
    wire signal_22517 ;
    wire signal_22518 ;
    wire signal_22519 ;
    wire signal_22520 ;
    wire signal_22521 ;
    wire signal_22522 ;
    wire signal_22523 ;
    wire signal_22524 ;
    wire signal_22525 ;
    wire signal_22526 ;
    wire signal_22527 ;
    wire signal_22528 ;
    wire signal_22529 ;
    wire signal_22530 ;
    wire signal_22531 ;
    wire signal_22532 ;
    wire signal_22533 ;
    wire signal_22534 ;
    wire signal_22535 ;
    wire signal_22536 ;
    wire signal_22537 ;
    wire signal_22538 ;
    wire signal_22539 ;
    wire signal_22540 ;
    wire signal_22541 ;
    wire signal_22542 ;
    wire signal_22543 ;
    wire signal_22544 ;
    wire signal_22545 ;
    wire signal_22546 ;
    wire signal_22547 ;
    wire signal_22548 ;
    wire signal_22549 ;
    wire signal_22550 ;
    wire signal_22551 ;
    wire signal_22552 ;
    wire signal_22553 ;
    wire signal_22554 ;
    wire signal_22555 ;
    wire signal_22556 ;
    wire signal_22557 ;
    wire signal_22558 ;
    wire signal_22559 ;
    wire signal_22560 ;
    wire signal_22561 ;
    wire signal_22562 ;
    wire signal_22563 ;
    wire signal_22564 ;
    wire signal_22565 ;
    wire signal_22566 ;
    wire signal_22567 ;
    wire signal_22568 ;
    wire signal_22569 ;
    wire signal_22570 ;
    wire signal_22571 ;
    wire signal_22572 ;
    wire signal_22573 ;
    wire signal_22574 ;
    wire signal_22575 ;
    wire signal_22576 ;
    wire signal_22577 ;
    wire signal_22578 ;
    wire signal_22579 ;
    wire signal_22580 ;
    wire signal_22581 ;
    wire signal_22582 ;
    wire signal_22583 ;
    wire signal_22584 ;
    wire signal_22585 ;
    wire signal_22586 ;
    wire signal_22587 ;
    wire signal_22588 ;
    wire signal_22589 ;
    wire signal_22590 ;
    wire signal_22591 ;
    wire signal_22592 ;
    wire signal_22593 ;
    wire signal_22594 ;
    wire signal_22595 ;
    wire signal_22596 ;
    wire signal_22597 ;
    wire signal_22598 ;
    wire signal_22599 ;
    wire signal_22600 ;
    wire signal_22601 ;
    wire signal_22602 ;
    wire signal_22603 ;
    wire signal_22604 ;
    wire signal_22605 ;
    wire signal_22606 ;
    wire signal_22607 ;
    wire signal_22608 ;
    wire signal_22609 ;
    wire signal_22610 ;
    wire signal_22611 ;
    wire signal_22612 ;
    wire signal_22613 ;
    wire signal_22614 ;
    wire signal_22615 ;
    wire signal_22616 ;
    wire signal_22617 ;
    wire signal_22618 ;
    wire signal_22619 ;
    wire signal_22620 ;
    wire signal_22621 ;
    wire signal_22622 ;
    wire signal_22623 ;
    wire signal_22624 ;
    wire signal_22625 ;
    wire signal_22626 ;
    wire signal_22627 ;
    wire signal_22628 ;
    wire signal_22629 ;
    wire signal_22630 ;
    wire signal_22631 ;
    wire signal_22632 ;
    wire signal_22633 ;
    wire signal_22634 ;
    wire signal_22635 ;
    wire signal_22636 ;
    wire signal_22637 ;
    wire signal_22638 ;
    wire signal_22639 ;
    wire signal_22640 ;
    wire signal_22641 ;
    wire signal_22642 ;
    wire signal_22643 ;
    wire signal_22644 ;
    wire signal_22645 ;
    wire signal_22646 ;
    wire signal_22647 ;
    wire signal_22648 ;
    wire signal_22649 ;
    wire signal_22650 ;
    wire signal_22651 ;
    wire signal_22652 ;
    wire signal_22653 ;
    wire signal_22654 ;
    wire signal_22655 ;
    wire signal_22656 ;
    wire signal_22657 ;
    wire signal_22658 ;
    wire signal_22659 ;
    wire signal_22660 ;
    wire signal_22661 ;
    wire signal_22662 ;
    wire signal_22663 ;
    wire signal_22664 ;
    wire signal_22665 ;
    wire signal_22666 ;
    wire signal_22667 ;
    wire signal_22668 ;
    wire signal_22669 ;
    wire signal_22670 ;
    wire signal_22671 ;
    wire signal_22672 ;
    wire signal_22673 ;
    wire signal_22674 ;
    wire signal_22675 ;
    wire signal_22676 ;
    wire signal_22677 ;
    wire signal_22678 ;
    wire signal_22679 ;
    wire signal_22680 ;
    wire signal_22681 ;
    wire signal_22682 ;
    wire signal_22683 ;
    wire signal_22684 ;
    wire signal_22685 ;
    wire signal_22686 ;
    wire signal_22687 ;
    wire signal_22688 ;
    wire signal_22689 ;
    wire signal_22690 ;
    wire signal_22691 ;
    wire signal_22692 ;
    wire signal_22693 ;
    wire signal_22694 ;
    wire signal_22695 ;
    wire signal_22696 ;
    wire signal_22697 ;
    wire signal_22698 ;
    wire signal_22699 ;
    wire signal_22700 ;
    wire signal_22701 ;
    wire signal_22702 ;
    wire signal_22703 ;
    wire signal_22704 ;
    wire signal_22705 ;
    wire signal_22706 ;
    wire signal_22707 ;
    wire signal_22708 ;
    wire signal_22709 ;
    wire signal_22710 ;
    wire signal_22711 ;
    wire signal_22712 ;
    wire signal_22713 ;
    wire signal_22714 ;
    wire signal_22715 ;
    wire signal_22716 ;
    wire signal_22717 ;
    wire signal_22718 ;
    wire signal_22719 ;
    wire signal_22720 ;
    wire signal_22721 ;
    wire signal_22722 ;
    wire signal_22723 ;
    wire signal_22724 ;
    wire signal_22725 ;
    wire signal_22726 ;
    wire signal_22727 ;
    wire signal_22728 ;
    wire signal_22729 ;
    wire signal_22730 ;
    wire signal_22731 ;
    wire signal_22732 ;
    wire signal_22733 ;
    wire signal_22734 ;
    wire signal_22735 ;
    wire signal_22736 ;
    wire signal_22737 ;
    wire signal_22738 ;
    wire signal_22739 ;
    wire signal_22740 ;
    wire signal_22741 ;
    wire signal_22742 ;
    wire signal_22743 ;
    wire signal_22744 ;
    wire signal_22745 ;
    wire signal_22746 ;
    wire signal_22747 ;
    wire signal_22748 ;
    wire signal_22749 ;
    wire signal_22750 ;
    wire signal_22751 ;
    wire signal_22752 ;
    wire signal_22753 ;
    wire signal_22754 ;
    wire signal_22755 ;
    wire signal_22756 ;
    wire signal_22757 ;
    wire signal_22758 ;
    wire signal_22759 ;
    wire signal_22760 ;
    wire signal_22761 ;
    wire signal_22762 ;
    wire signal_22763 ;
    wire signal_22764 ;
    wire signal_22765 ;
    wire signal_22766 ;
    wire signal_22767 ;
    wire signal_22768 ;
    wire signal_22769 ;
    wire signal_22770 ;
    wire signal_22771 ;
    wire signal_22772 ;
    wire signal_22773 ;
    wire signal_22774 ;
    wire signal_22775 ;
    wire signal_22776 ;
    wire signal_22777 ;
    wire signal_22778 ;
    wire signal_22779 ;
    wire signal_22780 ;
    wire signal_22781 ;
    wire signal_22782 ;
    wire signal_22783 ;
    wire signal_22784 ;
    wire signal_22785 ;
    wire signal_22786 ;
    wire signal_22787 ;
    wire signal_22788 ;
    wire signal_22789 ;
    wire signal_22790 ;
    wire signal_22791 ;
    wire signal_22792 ;
    wire signal_22793 ;
    wire signal_22794 ;
    wire signal_22795 ;
    wire signal_22796 ;
    wire signal_22797 ;
    wire signal_22798 ;
    wire signal_22799 ;
    wire signal_22800 ;
    wire signal_22801 ;
    wire signal_22802 ;
    wire signal_22803 ;
    wire signal_22804 ;
    wire signal_22805 ;
    wire signal_22806 ;
    wire signal_22807 ;
    wire signal_22808 ;
    wire signal_22809 ;
    wire signal_22810 ;
    wire signal_22811 ;
    wire signal_22812 ;
    wire signal_22813 ;
    wire signal_22814 ;
    wire signal_22815 ;
    wire signal_22816 ;
    wire signal_22817 ;
    wire signal_22818 ;
    wire signal_22819 ;
    wire signal_22820 ;
    wire signal_22821 ;
    wire signal_22822 ;
    wire signal_22823 ;
    wire signal_22824 ;
    wire signal_22825 ;
    wire signal_22826 ;
    wire signal_22827 ;
    wire signal_22828 ;
    wire signal_22829 ;
    wire signal_22830 ;
    wire signal_22831 ;
    wire signal_22832 ;
    wire signal_22833 ;
    wire signal_22834 ;
    wire signal_22835 ;
    wire signal_22836 ;
    wire signal_22837 ;
    wire signal_22838 ;
    wire signal_22839 ;
    wire signal_22840 ;
    wire signal_22841 ;
    wire signal_22842 ;
    wire signal_22843 ;
    wire signal_22844 ;
    wire signal_22845 ;
    wire signal_22846 ;
    wire signal_22847 ;
    wire signal_22848 ;
    wire signal_22849 ;
    wire signal_22850 ;
    wire signal_22851 ;
    wire signal_22852 ;
    wire signal_22853 ;
    wire signal_22854 ;
    wire signal_22855 ;
    wire signal_22856 ;
    wire signal_22857 ;
    wire signal_22858 ;
    wire signal_22859 ;
    wire signal_22860 ;
    wire signal_22861 ;
    wire signal_22862 ;
    wire signal_22863 ;
    wire signal_22864 ;
    wire signal_22865 ;
    wire signal_22866 ;
    wire signal_22867 ;
    wire signal_22868 ;
    wire signal_22869 ;
    wire signal_22870 ;
    wire signal_22871 ;
    wire signal_22872 ;
    wire signal_22873 ;
    wire signal_22874 ;
    wire signal_22875 ;
    wire signal_22876 ;
    wire signal_22877 ;
    wire signal_22878 ;
    wire signal_22879 ;
    wire signal_22880 ;
    wire signal_22881 ;
    wire signal_22882 ;
    wire signal_22883 ;
    wire signal_22884 ;
    wire signal_22885 ;
    wire signal_22886 ;
    wire signal_22887 ;
    wire signal_22888 ;
    wire signal_22889 ;
    wire signal_22890 ;
    wire signal_22891 ;
    wire signal_22892 ;
    wire signal_22893 ;
    wire signal_22894 ;
    wire signal_22895 ;
    wire signal_22896 ;
    wire signal_22897 ;
    wire signal_22898 ;
    wire signal_22899 ;
    wire signal_22900 ;
    wire signal_22901 ;
    wire signal_22902 ;
    wire signal_22903 ;
    wire signal_22904 ;
    wire signal_22905 ;
    wire signal_22906 ;
    wire signal_22907 ;
    wire signal_22908 ;
    wire signal_22909 ;
    wire signal_22910 ;
    wire signal_22911 ;
    wire signal_22912 ;
    wire signal_22913 ;
    wire signal_22914 ;
    wire signal_22915 ;
    wire signal_22916 ;
    wire signal_22917 ;
    wire signal_22918 ;
    wire signal_22919 ;
    wire signal_22920 ;
    wire signal_22921 ;
    wire signal_22922 ;
    wire signal_22923 ;
    wire signal_22924 ;
    wire signal_22925 ;
    wire signal_22926 ;
    wire signal_22927 ;
    wire signal_22928 ;
    wire signal_22929 ;
    wire signal_22930 ;
    wire signal_22931 ;
    wire signal_22932 ;
    wire signal_22933 ;
    wire signal_22934 ;
    wire signal_22935 ;
    wire signal_22936 ;
    wire signal_22937 ;
    wire signal_22938 ;
    wire signal_22939 ;
    wire signal_22940 ;
    wire signal_22941 ;
    wire signal_22942 ;
    wire signal_22943 ;
    wire signal_22944 ;
    wire signal_22945 ;
    wire signal_22946 ;
    wire signal_22947 ;
    wire signal_22948 ;
    wire signal_22949 ;
    wire signal_22950 ;
    wire signal_22951 ;
    wire signal_22952 ;
    wire signal_22953 ;
    wire signal_22954 ;
    wire signal_22955 ;
    wire signal_22956 ;
    wire signal_22957 ;
    wire signal_22958 ;
    wire signal_22959 ;
    wire signal_22960 ;
    wire signal_22961 ;
    wire signal_22962 ;
    wire signal_22963 ;
    wire signal_22964 ;
    wire signal_22965 ;
    wire signal_22966 ;
    wire signal_22967 ;
    wire signal_22968 ;
    wire signal_22969 ;
    wire signal_22970 ;
    wire signal_22971 ;
    wire signal_22972 ;
    wire signal_22973 ;
    wire signal_22974 ;
    wire signal_22975 ;
    wire signal_22976 ;
    wire signal_22977 ;
    wire signal_22978 ;
    wire signal_22979 ;
    wire signal_22980 ;
    wire signal_22981 ;
    wire signal_22982 ;
    wire signal_22983 ;
    wire signal_22984 ;
    wire signal_22985 ;
    wire signal_22986 ;
    wire signal_22987 ;
    wire signal_22988 ;
    wire signal_22989 ;
    wire signal_22990 ;
    wire signal_22991 ;
    wire signal_22992 ;
    wire signal_22993 ;
    wire signal_22994 ;
    wire signal_22995 ;
    wire signal_22996 ;
    wire signal_22997 ;
    wire signal_22998 ;
    wire signal_22999 ;
    wire signal_23000 ;
    wire signal_23001 ;
    wire signal_23002 ;
    wire signal_23003 ;
    wire signal_23004 ;
    wire signal_23005 ;
    wire signal_23006 ;
    wire signal_23007 ;
    wire signal_23008 ;
    wire signal_23009 ;
    wire signal_23010 ;
    wire signal_23011 ;
    wire signal_23012 ;
    wire signal_23013 ;
    wire signal_23014 ;
    wire signal_23015 ;
    wire signal_23016 ;
    wire signal_23017 ;
    wire signal_23018 ;
    wire signal_23019 ;
    wire signal_23020 ;
    wire signal_23021 ;
    wire signal_23022 ;
    wire signal_23023 ;
    wire signal_23024 ;
    wire signal_23025 ;
    wire signal_23026 ;
    wire signal_23027 ;
    wire signal_23028 ;
    wire signal_23029 ;
    wire signal_23030 ;
    wire signal_23031 ;
    wire signal_23032 ;
    wire signal_23033 ;
    wire signal_23034 ;
    wire signal_23035 ;
    wire signal_23036 ;
    wire signal_23037 ;
    wire signal_23038 ;
    wire signal_23039 ;
    wire signal_23040 ;
    wire signal_23041 ;
    wire signal_23042 ;
    wire signal_23043 ;
    wire signal_23044 ;
    wire signal_23045 ;
    wire signal_23046 ;
    wire signal_23047 ;
    wire signal_23048 ;
    wire signal_23049 ;
    wire signal_23050 ;
    wire signal_23051 ;
    wire signal_23052 ;
    wire signal_23053 ;
    wire signal_23054 ;
    wire signal_23055 ;
    wire signal_23056 ;
    wire signal_23057 ;
    wire signal_23058 ;
    wire signal_23059 ;
    wire signal_23060 ;
    wire signal_23061 ;
    wire signal_23062 ;
    wire signal_23063 ;
    wire signal_23064 ;
    wire signal_23065 ;
    wire signal_23066 ;
    wire signal_23067 ;
    wire signal_23068 ;
    wire signal_23069 ;
    wire signal_23070 ;
    wire signal_23071 ;
    wire signal_23072 ;
    wire signal_23073 ;
    wire signal_23074 ;
    wire signal_23075 ;
    wire signal_23076 ;
    wire signal_23077 ;
    wire signal_23078 ;
    wire signal_23079 ;
    wire signal_23080 ;
    wire signal_23081 ;
    wire signal_23082 ;
    wire signal_23083 ;
    wire signal_23084 ;
    wire signal_23085 ;
    wire signal_23086 ;
    wire signal_23087 ;
    wire signal_23088 ;
    wire signal_23089 ;
    wire signal_23090 ;
    wire signal_23091 ;
    wire signal_23092 ;
    wire signal_23093 ;
    wire signal_23094 ;
    wire signal_23095 ;
    wire signal_23096 ;
    wire signal_23097 ;
    wire signal_23098 ;
    wire signal_23099 ;
    wire signal_23100 ;
    wire signal_23101 ;
    wire signal_23102 ;
    wire signal_23103 ;
    wire signal_23104 ;
    wire signal_23105 ;
    wire signal_23106 ;
    wire signal_23107 ;
    wire signal_23108 ;
    wire signal_23109 ;
    wire signal_23110 ;
    wire signal_23111 ;
    wire signal_23112 ;
    wire signal_23113 ;
    wire signal_23114 ;
    wire signal_23115 ;
    wire signal_23116 ;
    wire signal_23117 ;
    wire signal_23118 ;
    wire signal_23119 ;
    wire signal_23120 ;
    wire signal_23121 ;
    wire signal_23122 ;
    wire signal_23123 ;
    wire signal_23124 ;
    wire signal_23125 ;
    wire signal_23126 ;
    wire signal_23127 ;
    wire signal_23128 ;
    wire signal_23129 ;
    wire signal_23130 ;
    wire signal_23131 ;
    wire signal_23132 ;
    wire signal_23133 ;
    wire signal_23134 ;
    wire signal_23135 ;
    wire signal_23136 ;
    wire signal_23137 ;
    wire signal_23138 ;
    wire signal_23139 ;
    wire signal_23140 ;
    wire signal_23141 ;
    wire signal_23142 ;
    wire signal_23143 ;
    wire signal_23144 ;
    wire signal_23145 ;
    wire signal_23146 ;
    wire signal_23147 ;
    wire signal_23148 ;
    wire signal_23149 ;
    wire signal_23150 ;
    wire signal_23151 ;
    wire signal_23152 ;
    wire signal_23153 ;
    wire signal_23154 ;
    wire signal_23155 ;
    wire signal_23156 ;
    wire signal_23157 ;
    wire signal_23158 ;
    wire signal_23159 ;
    wire signal_23160 ;
    wire signal_23161 ;
    wire signal_23162 ;
    wire signal_23163 ;
    wire signal_23164 ;
    wire signal_23165 ;
    wire signal_23166 ;
    wire signal_23167 ;
    wire signal_23168 ;
    wire signal_23169 ;
    wire signal_23170 ;
    wire signal_23171 ;
    wire signal_23172 ;
    wire signal_23173 ;
    wire signal_23174 ;
    wire signal_23175 ;
    wire signal_23176 ;
    wire signal_23177 ;
    wire signal_23178 ;
    wire signal_23179 ;
    wire signal_23180 ;
    wire signal_23181 ;
    wire signal_23182 ;
    wire signal_23183 ;
    wire signal_23184 ;
    wire signal_23185 ;
    wire signal_23186 ;
    wire signal_23187 ;
    wire signal_23188 ;
    wire signal_23189 ;
    wire signal_23190 ;
    wire signal_23191 ;
    wire signal_23192 ;
    wire signal_23193 ;
    wire signal_23194 ;
    wire signal_23195 ;
    wire signal_23196 ;
    wire signal_23197 ;
    wire signal_23198 ;
    wire signal_23199 ;
    wire signal_23200 ;
    wire signal_23201 ;
    wire signal_23202 ;
    wire signal_23203 ;
    wire signal_23204 ;
    wire signal_23205 ;
    wire signal_23206 ;
    wire signal_23207 ;
    wire signal_23208 ;
    wire signal_23209 ;
    wire signal_23210 ;
    wire signal_23211 ;
    wire signal_23212 ;
    wire signal_23213 ;
    wire signal_23214 ;
    wire signal_23215 ;
    wire signal_23216 ;
    wire signal_23217 ;
    wire signal_23218 ;
    wire signal_23219 ;
    wire signal_23220 ;
    wire signal_23221 ;
    wire signal_23222 ;
    wire signal_23223 ;
    wire signal_23224 ;
    wire signal_23225 ;
    wire signal_23226 ;
    wire signal_23227 ;
    wire signal_23228 ;
    wire signal_23229 ;
    wire signal_23230 ;
    wire signal_23231 ;
    wire signal_23232 ;
    wire signal_23233 ;
    wire signal_23234 ;
    wire signal_23235 ;
    wire signal_23236 ;
    wire signal_23237 ;
    wire signal_23238 ;
    wire signal_23239 ;
    wire signal_23240 ;
    wire signal_23241 ;
    wire signal_23242 ;
    wire signal_23243 ;
    wire signal_23244 ;
    wire signal_23245 ;
    wire signal_23246 ;
    wire signal_23247 ;
    wire signal_23248 ;
    wire signal_23249 ;
    wire signal_23250 ;
    wire signal_23251 ;
    wire signal_23252 ;
    wire signal_23253 ;
    wire signal_23254 ;
    wire signal_23255 ;
    wire signal_23256 ;
    wire signal_23257 ;
    wire signal_23258 ;
    wire signal_23259 ;
    wire signal_23260 ;
    wire signal_23261 ;
    wire signal_23262 ;
    wire signal_23263 ;
    wire signal_23264 ;
    wire signal_23265 ;
    wire signal_23266 ;
    wire signal_23267 ;
    wire signal_23268 ;
    wire signal_23269 ;
    wire signal_23270 ;
    wire signal_23271 ;
    wire signal_23272 ;
    wire signal_23273 ;
    wire signal_23274 ;
    wire signal_23275 ;
    wire signal_23276 ;
    wire signal_23277 ;
    wire signal_23278 ;
    wire signal_23279 ;
    wire signal_23280 ;
    wire signal_23281 ;
    wire signal_23282 ;
    wire signal_23283 ;
    wire signal_23284 ;
    wire signal_23285 ;
    wire signal_23286 ;
    wire signal_23287 ;
    wire signal_23288 ;
    wire signal_23289 ;
    wire signal_23290 ;
    wire signal_23291 ;
    wire signal_23292 ;
    wire signal_23293 ;
    wire signal_23294 ;
    wire signal_23295 ;
    wire signal_23296 ;
    wire signal_23297 ;
    wire signal_23298 ;
    wire signal_23299 ;
    wire signal_23300 ;
    wire signal_23301 ;
    wire signal_23302 ;
    wire signal_23303 ;
    wire signal_23304 ;
    wire signal_23305 ;
    wire signal_23306 ;
    wire signal_23307 ;
    wire signal_23308 ;
    wire signal_23309 ;
    wire signal_23310 ;
    wire signal_23311 ;
    wire signal_23312 ;
    wire signal_23313 ;
    wire signal_23314 ;
    wire signal_23315 ;
    wire signal_23316 ;
    wire signal_23317 ;
    wire signal_23318 ;
    wire signal_23319 ;
    wire signal_23320 ;
    wire signal_23321 ;
    wire signal_23322 ;
    wire signal_23323 ;
    wire signal_23324 ;
    wire signal_23325 ;
    wire signal_23326 ;
    wire signal_23327 ;
    wire signal_23328 ;
    wire signal_23329 ;
    wire signal_23330 ;
    wire signal_23331 ;
    wire signal_23332 ;
    wire signal_23333 ;
    wire signal_23334 ;
    wire signal_23335 ;
    wire signal_23336 ;
    wire signal_23337 ;
    wire signal_23338 ;
    wire signal_23339 ;
    wire signal_23340 ;
    wire signal_23341 ;
    wire signal_23342 ;
    wire signal_23343 ;
    wire signal_23344 ;
    wire signal_23345 ;
    wire signal_23346 ;
    wire signal_23347 ;
    wire signal_23348 ;
    wire signal_23349 ;
    wire signal_23350 ;
    wire signal_23351 ;
    wire signal_23352 ;
    wire signal_23353 ;
    wire signal_23354 ;
    wire signal_23355 ;
    wire signal_23356 ;
    wire signal_23357 ;
    wire signal_23358 ;
    wire signal_23359 ;
    wire signal_23360 ;
    wire signal_23361 ;
    wire signal_23362 ;
    wire signal_23363 ;
    wire signal_23364 ;
    wire signal_23365 ;
    wire signal_23366 ;
    wire signal_23367 ;
    wire signal_23368 ;
    wire signal_23369 ;
    wire signal_23370 ;
    wire signal_23371 ;
    wire signal_23372 ;
    wire signal_23373 ;
    wire signal_23374 ;
    wire signal_23375 ;
    wire signal_23376 ;
    wire signal_23377 ;
    wire signal_23378 ;
    wire signal_23379 ;
    wire signal_23380 ;
    wire signal_23381 ;
    wire signal_23382 ;
    wire signal_23383 ;
    wire signal_23384 ;
    wire signal_23385 ;
    wire signal_23386 ;
    wire signal_23387 ;
    wire signal_23388 ;
    wire signal_23389 ;
    wire signal_23390 ;
    wire signal_23391 ;
    wire signal_23392 ;
    wire signal_23393 ;
    wire signal_23394 ;
    wire signal_23395 ;
    wire signal_23396 ;
    wire signal_23397 ;
    wire signal_23398 ;
    wire signal_23399 ;
    wire signal_23400 ;
    wire signal_23401 ;
    wire signal_23402 ;
    wire signal_23403 ;
    wire signal_23404 ;
    wire signal_23405 ;
    wire signal_23406 ;
    wire signal_23407 ;
    wire signal_23408 ;
    wire signal_23409 ;
    wire signal_23410 ;
    wire signal_23411 ;
    wire signal_23412 ;
    wire signal_23413 ;
    wire signal_23414 ;
    wire signal_23415 ;
    wire signal_23416 ;
    wire signal_23417 ;
    wire signal_23418 ;
    wire signal_23419 ;
    wire signal_23420 ;
    wire signal_23421 ;
    wire signal_23422 ;
    wire signal_23423 ;
    wire signal_23424 ;
    wire signal_23425 ;
    wire signal_23426 ;
    wire signal_23427 ;
    wire signal_23428 ;
    wire signal_23429 ;
    wire signal_23430 ;
    wire signal_23431 ;
    wire signal_23432 ;
    wire signal_23433 ;
    wire signal_23434 ;
    wire signal_23435 ;
    wire signal_23436 ;
    wire signal_23437 ;
    wire signal_23438 ;
    wire signal_23439 ;
    wire signal_23440 ;
    wire signal_23441 ;
    wire signal_23442 ;
    wire signal_23443 ;
    wire signal_23444 ;
    wire signal_23445 ;
    wire signal_23446 ;
    wire signal_23447 ;
    wire signal_23448 ;
    wire signal_23449 ;
    wire signal_23450 ;
    wire signal_23451 ;
    wire signal_23452 ;
    wire signal_23453 ;
    wire signal_23454 ;
    wire signal_23455 ;
    wire signal_23456 ;
    wire signal_23457 ;
    wire signal_23458 ;
    wire signal_23459 ;
    wire signal_23460 ;
    wire signal_23461 ;
    wire signal_23462 ;
    wire signal_23463 ;
    wire signal_23464 ;
    wire signal_23465 ;
    wire signal_23466 ;
    wire signal_23467 ;
    wire signal_23468 ;
    wire signal_23469 ;
    wire signal_23470 ;
    wire signal_23471 ;
    wire signal_23472 ;
    wire signal_23473 ;
    wire signal_23474 ;
    wire signal_23475 ;
    wire signal_23476 ;
    wire signal_23477 ;
    wire signal_23478 ;
    wire signal_23479 ;
    wire signal_23480 ;
    wire signal_23481 ;
    wire signal_23482 ;
    wire signal_23483 ;
    wire signal_23484 ;
    wire signal_23485 ;
    wire signal_23486 ;
    wire signal_23487 ;
    wire signal_23488 ;
    wire signal_23489 ;
    wire signal_23490 ;
    wire signal_23491 ;
    wire signal_23492 ;
    wire signal_23493 ;
    wire signal_23494 ;
    wire signal_23495 ;
    wire signal_23496 ;
    wire signal_23497 ;
    wire signal_23498 ;
    wire signal_23499 ;
    wire signal_23500 ;
    wire signal_23501 ;
    wire signal_23502 ;
    wire signal_23503 ;
    wire signal_23504 ;
    wire signal_23505 ;
    wire signal_23506 ;
    wire signal_23507 ;
    wire signal_23508 ;
    wire signal_23509 ;
    wire signal_23510 ;
    wire signal_23511 ;
    wire signal_23512 ;
    wire signal_23513 ;
    wire signal_23514 ;
    wire signal_23515 ;
    wire signal_23516 ;
    wire signal_23517 ;
    wire signal_23518 ;
    wire signal_23519 ;
    wire signal_23520 ;
    wire signal_23521 ;
    wire signal_23522 ;
    wire signal_23523 ;
    wire signal_23524 ;
    wire signal_23525 ;
    wire signal_23526 ;
    wire signal_23527 ;
    wire signal_23528 ;
    wire signal_23529 ;
    wire signal_23530 ;
    wire signal_23531 ;
    wire signal_23532 ;
    wire signal_23533 ;
    wire signal_23534 ;
    wire signal_23535 ;
    wire signal_23536 ;
    wire signal_23537 ;
    wire signal_23538 ;
    wire signal_23539 ;
    wire signal_23540 ;
    wire signal_23541 ;
    wire signal_23542 ;
    wire signal_23543 ;
    wire signal_23544 ;
    wire signal_23545 ;
    wire signal_23546 ;
    wire signal_23547 ;
    wire signal_23548 ;
    wire signal_23549 ;
    wire signal_23550 ;
    wire signal_23551 ;
    wire signal_23552 ;
    wire signal_23553 ;
    wire signal_23554 ;
    wire signal_23555 ;
    wire signal_23556 ;
    wire signal_23557 ;
    wire signal_23558 ;
    wire signal_23559 ;
    wire signal_23560 ;
    wire signal_23561 ;
    wire signal_23562 ;
    wire signal_23563 ;
    wire signal_23564 ;
    wire signal_23565 ;
    wire signal_23566 ;
    wire signal_23567 ;
    wire signal_23568 ;
    wire signal_23569 ;
    wire signal_23570 ;
    wire signal_23571 ;
    wire signal_23572 ;
    wire signal_23573 ;
    wire signal_23574 ;
    wire signal_23575 ;
    wire signal_23576 ;
    wire signal_23577 ;
    wire signal_23578 ;
    wire signal_23579 ;
    wire signal_23580 ;
    wire signal_23581 ;
    wire signal_23582 ;
    wire signal_23583 ;
    wire signal_23584 ;
    wire signal_23585 ;
    wire signal_23586 ;
    wire signal_23587 ;
    wire signal_23588 ;
    wire signal_23589 ;
    wire signal_23590 ;
    wire signal_23591 ;
    wire signal_23592 ;
    wire signal_23593 ;
    wire signal_23594 ;
    wire signal_23595 ;
    wire signal_23596 ;
    wire signal_23597 ;
    wire signal_23598 ;
    wire signal_23599 ;
    wire signal_23600 ;
    wire signal_23601 ;
    wire signal_23602 ;
    wire signal_23603 ;
    wire signal_23604 ;
    wire signal_23605 ;
    wire signal_23606 ;
    wire signal_23607 ;
    wire signal_23608 ;
    wire signal_23609 ;
    wire signal_23610 ;
    wire signal_23611 ;
    wire signal_23612 ;
    wire signal_23613 ;
    wire signal_23614 ;
    wire signal_23615 ;
    wire signal_23616 ;
    wire signal_23617 ;
    wire signal_23618 ;
    wire signal_23619 ;
    wire signal_23620 ;
    wire signal_23621 ;
    wire signal_23622 ;
    wire signal_23623 ;
    wire signal_23624 ;
    wire signal_23625 ;
    wire signal_23626 ;
    wire signal_23627 ;
    wire signal_23628 ;
    wire signal_23629 ;
    wire signal_23630 ;
    wire signal_23631 ;
    wire signal_23632 ;
    wire signal_23633 ;
    wire signal_23634 ;
    wire signal_23635 ;
    wire signal_23636 ;
    wire signal_23637 ;
    wire signal_23638 ;
    wire signal_23639 ;
    wire signal_23640 ;
    wire signal_23641 ;
    wire signal_23642 ;
    wire signal_23643 ;
    wire signal_23644 ;
    wire signal_23645 ;
    wire signal_23646 ;
    wire signal_23647 ;
    wire signal_23648 ;
    wire signal_23649 ;
    wire signal_23650 ;
    wire signal_23651 ;
    wire signal_23652 ;
    wire signal_23653 ;
    wire signal_23654 ;
    wire signal_23655 ;
    wire signal_23656 ;
    wire signal_23657 ;
    wire signal_23658 ;
    wire signal_23659 ;
    wire signal_23660 ;
    wire signal_23661 ;
    wire signal_23662 ;
    wire signal_23663 ;
    wire signal_23664 ;
    wire signal_23665 ;
    wire signal_23666 ;
    wire signal_23667 ;
    wire signal_23668 ;
    wire signal_23669 ;
    wire signal_23670 ;
    wire signal_23671 ;
    wire signal_23672 ;
    wire signal_23673 ;
    wire signal_23674 ;
    wire signal_23675 ;
    wire signal_23676 ;
    wire signal_23677 ;
    wire signal_23678 ;
    wire signal_23679 ;
    wire signal_23680 ;
    wire signal_23681 ;
    wire signal_23682 ;
    wire signal_23683 ;
    wire signal_23684 ;
    wire signal_23685 ;
    wire signal_23686 ;
    wire signal_23687 ;
    wire signal_23688 ;
    wire signal_23689 ;
    wire signal_23690 ;
    wire signal_23691 ;
    wire signal_23692 ;
    wire signal_23693 ;
    wire signal_23694 ;
    wire signal_23695 ;
    wire signal_23696 ;
    wire signal_23697 ;
    wire signal_23698 ;
    wire signal_23699 ;
    wire signal_23700 ;
    wire signal_23701 ;
    wire signal_23702 ;
    wire signal_23703 ;
    wire signal_23704 ;
    wire signal_23705 ;
    wire signal_23706 ;
    wire signal_23707 ;
    wire signal_23708 ;
    wire signal_23709 ;
    wire signal_23710 ;
    wire signal_23711 ;
    wire signal_23712 ;
    wire signal_23713 ;
    wire signal_23714 ;
    wire signal_23715 ;
    wire signal_23716 ;
    wire signal_23717 ;
    wire signal_23718 ;
    wire signal_23719 ;
    wire signal_23720 ;
    wire signal_23721 ;
    wire signal_23722 ;
    wire signal_23723 ;
    wire signal_23724 ;
    wire signal_23725 ;
    wire signal_23726 ;
    wire signal_23727 ;
    wire signal_23728 ;
    wire signal_23729 ;
    wire signal_23730 ;
    wire signal_23731 ;
    wire signal_23732 ;
    wire signal_23733 ;
    wire signal_23734 ;
    wire signal_23735 ;
    wire signal_23736 ;
    wire signal_23737 ;
    wire signal_23738 ;
    wire signal_23739 ;
    wire signal_23740 ;
    wire signal_23741 ;
    wire signal_23742 ;
    wire signal_23743 ;
    wire signal_23744 ;
    wire signal_23745 ;
    wire signal_23746 ;
    wire signal_23747 ;
    wire signal_23748 ;
    wire signal_23749 ;
    wire signal_23750 ;
    wire signal_23751 ;
    wire signal_23752 ;
    wire signal_23753 ;
    wire signal_23754 ;
    wire signal_23755 ;
    wire signal_23756 ;
    wire signal_23757 ;
    wire signal_23758 ;
    wire signal_23759 ;
    wire signal_23760 ;
    wire signal_23761 ;
    wire signal_23762 ;
    wire signal_23763 ;
    wire signal_23764 ;
    wire signal_23765 ;
    wire signal_23766 ;
    wire signal_23767 ;
    wire signal_23768 ;
    wire signal_23769 ;
    wire signal_23770 ;
    wire signal_23771 ;
    wire signal_23772 ;
    wire signal_23773 ;
    wire signal_23774 ;
    wire signal_23775 ;
    wire signal_23776 ;
    wire signal_23777 ;
    wire signal_23778 ;
    wire signal_23779 ;
    wire signal_23780 ;
    wire signal_23781 ;
    wire signal_23782 ;
    wire signal_23783 ;
    wire signal_23784 ;
    wire signal_23785 ;
    wire signal_23786 ;
    wire signal_23787 ;
    wire signal_23788 ;
    wire signal_23789 ;
    wire signal_23790 ;
    wire signal_23791 ;
    wire signal_23792 ;
    wire signal_23793 ;
    wire signal_23794 ;
    wire signal_23795 ;
    wire signal_23796 ;
    wire signal_23797 ;
    wire signal_23798 ;
    wire signal_23799 ;
    wire signal_23800 ;
    wire signal_23801 ;
    wire signal_23802 ;
    wire signal_23803 ;
    wire signal_23804 ;
    wire signal_23805 ;
    wire signal_23806 ;
    wire signal_23807 ;
    wire signal_23808 ;
    wire signal_23809 ;
    wire signal_23810 ;
    wire signal_23811 ;
    wire signal_23812 ;
    wire signal_23813 ;
    wire signal_23814 ;
    wire signal_23815 ;
    wire signal_23816 ;
    wire signal_23817 ;
    wire signal_23818 ;
    wire signal_23819 ;
    wire signal_23820 ;
    wire signal_23821 ;
    wire signal_23822 ;
    wire signal_23823 ;
    wire signal_23824 ;
    wire signal_23825 ;
    wire signal_23826 ;
    wire signal_23827 ;
    wire signal_23828 ;
    wire signal_23829 ;
    wire signal_23830 ;
    wire signal_23831 ;
    wire signal_23832 ;
    wire signal_23833 ;
    wire signal_23834 ;
    wire signal_23835 ;
    wire signal_23836 ;
    wire signal_23837 ;
    wire signal_23838 ;
    wire signal_23839 ;
    wire signal_23840 ;
    wire signal_23841 ;
    wire signal_23842 ;
    wire signal_23843 ;
    wire signal_23844 ;
    wire signal_23845 ;
    wire signal_23846 ;
    wire signal_23847 ;
    wire signal_23848 ;
    wire signal_23849 ;
    wire signal_23850 ;
    wire signal_23851 ;
    wire signal_23852 ;
    wire signal_23853 ;
    wire signal_23854 ;
    wire signal_23855 ;
    wire signal_23856 ;
    wire signal_23857 ;
    wire signal_23858 ;
    wire signal_23859 ;
    wire signal_23860 ;
    wire signal_23861 ;
    wire signal_23862 ;
    wire signal_23863 ;
    wire signal_23864 ;
    wire signal_23865 ;
    wire signal_23866 ;
    wire signal_23867 ;
    wire signal_23868 ;
    wire signal_23869 ;
    wire signal_23870 ;
    wire signal_23871 ;
    wire signal_23872 ;
    wire signal_23873 ;
    wire signal_23874 ;
    wire signal_23875 ;
    wire signal_23876 ;
    wire signal_23877 ;
    wire signal_23878 ;
    wire signal_23879 ;
    wire signal_23880 ;
    wire signal_23881 ;
    wire signal_23882 ;
    wire signal_23883 ;
    wire signal_23884 ;
    wire signal_23885 ;
    wire signal_23886 ;
    wire signal_23887 ;
    wire signal_23888 ;
    wire signal_23889 ;
    wire signal_23890 ;
    wire signal_23891 ;
    wire signal_23892 ;
    wire signal_23893 ;
    wire signal_23894 ;
    wire signal_23895 ;
    wire signal_23896 ;
    wire signal_23897 ;
    wire signal_23898 ;
    wire signal_23899 ;
    wire signal_23900 ;
    wire signal_23901 ;
    wire signal_23902 ;
    wire signal_23903 ;
    wire signal_23904 ;
    wire signal_23905 ;
    wire signal_23906 ;
    wire signal_23907 ;
    wire signal_23908 ;
    wire signal_23909 ;
    wire signal_23910 ;
    wire signal_23911 ;
    wire signal_23912 ;
    wire signal_23913 ;
    wire signal_23914 ;
    wire signal_23915 ;
    wire signal_23916 ;
    wire signal_23917 ;
    wire signal_23918 ;
    wire signal_23919 ;
    wire signal_23920 ;
    wire signal_23921 ;
    wire signal_23922 ;
    wire signal_23923 ;
    wire signal_23924 ;
    wire signal_23925 ;
    wire signal_23926 ;
    wire signal_23927 ;
    wire signal_23928 ;
    wire signal_23929 ;
    wire signal_23930 ;
    wire signal_23931 ;
    wire signal_23932 ;
    wire signal_23933 ;
    wire signal_23934 ;
    wire signal_23935 ;
    wire signal_23936 ;
    wire signal_23937 ;
    wire signal_23938 ;
    wire signal_23939 ;
    wire signal_23940 ;
    wire signal_23941 ;
    wire signal_23942 ;
    wire signal_23943 ;
    wire signal_23944 ;
    wire signal_23945 ;
    wire signal_23946 ;
    wire signal_23947 ;
    wire signal_23948 ;
    wire signal_23949 ;
    wire signal_23950 ;
    wire signal_23951 ;
    wire signal_23952 ;
    wire signal_23953 ;
    wire signal_23954 ;
    wire signal_23955 ;
    wire signal_23956 ;
    wire signal_23957 ;
    wire signal_23958 ;
    wire signal_23959 ;
    wire signal_23960 ;
    wire signal_23961 ;
    wire signal_23962 ;
    wire signal_23963 ;
    wire signal_23964 ;
    wire signal_23965 ;
    wire signal_23966 ;
    wire signal_23967 ;
    wire signal_23968 ;
    wire signal_23969 ;
    wire signal_23970 ;
    wire signal_23971 ;
    wire signal_23972 ;
    wire signal_23973 ;
    wire signal_23974 ;
    wire signal_23975 ;
    wire signal_23976 ;
    wire signal_23977 ;
    wire signal_23978 ;
    wire signal_23979 ;
    wire signal_23980 ;
    wire signal_23981 ;
    wire signal_23982 ;
    wire signal_23983 ;
    wire signal_23984 ;
    wire signal_23985 ;
    wire signal_23986 ;
    wire signal_23987 ;
    wire signal_23988 ;
    wire signal_23989 ;
    wire signal_23990 ;
    wire signal_23991 ;
    wire signal_23992 ;
    wire signal_23993 ;
    wire signal_23994 ;
    wire signal_23995 ;
    wire signal_23996 ;
    wire signal_23997 ;
    wire signal_23998 ;
    wire signal_23999 ;
    wire signal_24000 ;
    wire signal_24001 ;
    wire signal_24002 ;
    wire signal_24003 ;
    wire signal_24004 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_400) ) ;
    INV_X1 cell_1 ( .A (signal_395), .ZN (signal_401) ) ;
    INV_X1 cell_2 ( .A (signal_395), .ZN (signal_398) ) ;
    INV_X1 cell_3 ( .A (signal_395), .ZN (signal_396) ) ;
    INV_X1 cell_4 ( .A (signal_395), .ZN (signal_397) ) ;
    INV_X1 cell_5 ( .A (signal_395), .ZN (signal_399) ) ;
    NOR2_X1 cell_6 ( .A1 (signal_406), .A2 (signal_411), .ZN (signal_395) ) ;
    INV_X1 cell_7 ( .A (signal_4388), .ZN (signal_406) ) ;
    INV_X1 cell_8 ( .A (signal_395), .ZN (signal_402) ) ;
    NOR2_X1 cell_9 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_404) ) ;
    INV_X1 cell_10 ( .A (signal_404), .ZN (signal_403) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_4388), .A2 (signal_403), .ZN (signal_4384) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_4388), .A2 (signal_4385), .ZN (signal_418) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_418), .A2 (signal_403), .ZN (signal_4383) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_4385), .A2 (signal_404), .ZN (signal_411) ) ;
    INV_X1 cell_15 ( .A (signal_4386), .ZN (signal_409) ) ;
    AND2_X1 cell_16 ( .A1 (signal_409), .A2 (signal_4387), .ZN (signal_414) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_418), .A2 (signal_414), .ZN (signal_405) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_402), .A2 (signal_405), .ZN (signal_4382) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_4385), .A2 (signal_406), .ZN (signal_416) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_414), .A2 (signal_416), .ZN (signal_408) ) ;
    NAND2_X1 cell_21 ( .A1 (signal_4385), .A2 (signal_4384), .ZN (signal_407) ) ;
    NAND2_X1 cell_22 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_4381) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_4387), .A2 (signal_409), .ZN (signal_412) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_418), .A2 (signal_412), .ZN (signal_410) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_411), .A2 (signal_410), .ZN (signal_4380) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_416), .A2 (signal_412), .ZN (signal_413) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_402), .A2 (signal_413), .ZN (signal_4379) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .a ({signal_7457, signal_3750}), .b ({signal_7458, signal_4258}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .a ({signal_7460, signal_3749}), .b ({signal_7461, signal_4257}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .a ({signal_7463, signal_3748}), .b ({signal_7464, signal_4256}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .a ({signal_7466, signal_3747}), .b ({signal_7467, signal_4255}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .a ({signal_7469, signal_3746}), .b ({signal_7470, signal_4254}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .a ({signal_7472, signal_3745}), .b ({signal_7473, signal_4253}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .a ({signal_7475, signal_3744}), .b ({signal_7476, signal_4252}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .a ({signal_7478, signal_3743}), .b ({signal_7479, signal_4251}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({signal_7481, signal_3814}), .b ({signal_7482, signal_4322}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({signal_7484, signal_3813}), .b ({signal_7485, signal_4321}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({signal_7487, signal_3812}), .b ({signal_7488, signal_4320}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({signal_7490, signal_3811}), .b ({signal_7491, signal_4319}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({signal_7493, signal_3810}), .b ({signal_7494, signal_4318}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({signal_7496, signal_3809}), .b ({signal_7497, signal_4317}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({signal_7499, signal_3808}), .b ({signal_7500, signal_4316}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({signal_7502, signal_3807}), .b ({signal_7503, signal_4315}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({signal_7505, signal_3782}), .b ({signal_7506, signal_4290}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({signal_7508, signal_3781}), .b ({signal_7509, signal_4289}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({signal_7511, signal_3780}), .b ({signal_7512, signal_4288}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({signal_7514, signal_3779}), .b ({signal_7515, signal_4287}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({signal_7517, signal_3778}), .b ({signal_7518, signal_4286}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({signal_7520, signal_3777}), .b ({signal_7521, signal_4285}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({signal_7523, signal_3776}), .b ({signal_7524, signal_4284}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({signal_7526, signal_3775}), .b ({signal_7527, signal_4283}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    NAND2_X1 cell_284 ( .A1 (signal_4385), .A2 (signal_414), .ZN (signal_415) ) ;
    NOR2_X1 cell_285 ( .A1 (signal_4388), .A2 (signal_415), .ZN (done) ) ;
    INV_X1 cell_286 ( .A (signal_416), .ZN (signal_417) ) ;
    NAND2_X1 cell_287 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_419) ) ;
    NOR2_X1 cell_288 ( .A1 (signal_417), .A2 (signal_419), .ZN (signal_393) ) ;
    INV_X1 cell_289 ( .A (signal_418), .ZN (signal_420) ) ;
    NOR2_X1 cell_290 ( .A1 (signal_420), .A2 (signal_419), .ZN (signal_394) ) ;
    INV_X1 cell_4187 ( .A (signal_3597), .ZN (signal_3607) ) ;
    MUX2_X1 cell_4188 ( .S (signal_3609), .A (signal_3598), .B (signal_3599), .Z (signal_3597) ) ;
    NOR2_X1 cell_4189 ( .A1 (reset), .A2 (signal_3600), .ZN (signal_3610) ) ;
    XNOR2_X1 cell_4190 ( .A (signal_4388), .B (signal_4387), .ZN (signal_3600) ) ;
    MUX2_X1 cell_4191 ( .S (signal_4385), .A (signal_3601), .B (signal_3602), .Z (signal_3608) ) ;
    NAND2_X1 cell_4192 ( .A1 (signal_3598), .A2 (signal_3603), .ZN (signal_3602) ) ;
    NAND2_X1 cell_4193 ( .A1 (signal_3609), .A2 (signal_3606), .ZN (signal_3603) ) ;
    NOR2_X1 cell_4194 ( .A1 (signal_3604), .A2 (signal_3612), .ZN (signal_3598) ) ;
    NOR2_X1 cell_4195 ( .A1 (signal_4387), .A2 (reset), .ZN (signal_3604) ) ;
    NOR2_X1 cell_4196 ( .A1 (signal_3609), .A2 (signal_3599), .ZN (signal_3601) ) ;
    NAND2_X1 cell_4197 ( .A1 (signal_4387), .A2 (signal_3605), .ZN (signal_3599) ) ;
    NOR2_X1 cell_4198 ( .A1 (reset), .A2 (signal_3611), .ZN (signal_3605) ) ;
    NOR2_X1 cell_4199 ( .A1 (reset), .A2 (signal_4388), .ZN (signal_3612) ) ;
    INV_X1 cell_4200 ( .A (reset), .ZN (signal_3606) ) ;
    INV_X1 cell_4201 ( .A (signal_4388), .ZN (signal_3611) ) ;
    INV_X1 cell_4205 ( .A (signal_4386), .ZN (signal_3609) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4209 ( .a ({signal_7529, signal_4378}), .b ({signal_7530, signal_3870}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4210 ( .a ({signal_7532, signal_4278}), .b ({signal_7533, signal_3770}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4211 ( .a ({signal_7535, signal_4277}), .b ({signal_7536, signal_3769}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4212 ( .a ({signal_7538, signal_4276}), .b ({signal_7539, signal_3768}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4213 ( .a ({signal_7541, signal_4275}), .b ({signal_7542, signal_3767}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4214 ( .a ({signal_7544, signal_4274}), .b ({signal_7545, signal_3766}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4215 ( .a ({signal_7547, signal_4273}), .b ({signal_7548, signal_3765}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4216 ( .a ({signal_7550, signal_4272}), .b ({signal_7551, signal_3764}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4217 ( .a ({signal_7553, signal_4271}), .b ({signal_7554, signal_3763}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4218 ( .a ({signal_7556, signal_4270}), .b ({signal_7557, signal_3762}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4219 ( .a ({signal_7559, signal_4269}), .b ({signal_7560, signal_3761}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4220 ( .a ({signal_7562, signal_4368}), .b ({signal_7563, signal_3860}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4221 ( .a ({signal_7565, signal_4268}), .b ({signal_7566, signal_3760}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4222 ( .a ({signal_7568, signal_4267}), .b ({signal_7569, signal_3759}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4223 ( .a ({signal_7571, signal_4266}), .b ({signal_7572, signal_3758}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4224 ( .a ({signal_7574, signal_4265}), .b ({signal_7575, signal_3757}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4225 ( .a ({signal_7577, signal_4264}), .b ({signal_7578, signal_3756}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4226 ( .a ({signal_7580, signal_4263}), .b ({signal_7581, signal_3755}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4227 ( .a ({signal_7583, signal_4262}), .b ({signal_7584, signal_3754}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4228 ( .a ({signal_7586, signal_4261}), .b ({signal_7587, signal_3753}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4229 ( .a ({signal_7589, signal_4260}), .b ({signal_7590, signal_3752}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4230 ( .a ({signal_7592, signal_4259}), .b ({signal_7593, signal_3751}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4231 ( .a ({signal_7595, signal_4367}), .b ({signal_7596, signal_3859}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4232 ( .a ({signal_7598, signal_4366}), .b ({signal_7599, signal_3858}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4233 ( .a ({signal_7601, signal_4365}), .b ({signal_7602, signal_3857}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4234 ( .a ({signal_7604, signal_4364}), .b ({signal_7605, signal_3856}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4235 ( .a ({signal_7607, signal_4363}), .b ({signal_7608, signal_3855}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4236 ( .a ({signal_7610, signal_4362}), .b ({signal_7611, signal_3854}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4237 ( .a ({signal_7613, signal_4361}), .b ({signal_7614, signal_3853}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4238 ( .a ({signal_7616, signal_4360}), .b ({signal_7617, signal_3852}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4239 ( .a ({signal_7619, signal_4359}), .b ({signal_7620, signal_3851}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4240 ( .a ({signal_7622, signal_4377}), .b ({signal_7623, signal_3869}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4241 ( .a ({signal_7625, signal_4358}), .b ({signal_7626, signal_3850}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4242 ( .a ({signal_7628, signal_4357}), .b ({signal_7629, signal_3849}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4243 ( .a ({signal_7631, signal_4356}), .b ({signal_7632, signal_3848}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4244 ( .a ({signal_7634, signal_4355}), .b ({signal_7635, signal_3847}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4245 ( .a ({signal_7637, signal_4354}), .b ({signal_7638, signal_3846}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4246 ( .a ({signal_7640, signal_4353}), .b ({signal_7641, signal_3845}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4247 ( .a ({signal_7643, signal_4352}), .b ({signal_7644, signal_3844}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4248 ( .a ({signal_7646, signal_4351}), .b ({signal_7647, signal_3843}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4249 ( .a ({signal_7649, signal_4350}), .b ({signal_7650, signal_3842}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4250 ( .a ({signal_7652, signal_4349}), .b ({signal_7653, signal_3841}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4251 ( .a ({signal_7655, signal_4376}), .b ({signal_7656, signal_3868}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4252 ( .a ({signal_7658, signal_4348}), .b ({signal_7659, signal_3840}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4253 ( .a ({signal_7661, signal_4347}), .b ({signal_7662, signal_3839}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4254 ( .a ({signal_7664, signal_4346}), .b ({signal_7665, signal_3838}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4255 ( .a ({signal_7667, signal_4345}), .b ({signal_7668, signal_3837}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4256 ( .a ({signal_7670, signal_4344}), .b ({signal_7671, signal_3836}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4257 ( .a ({signal_7673, signal_4343}), .b ({signal_7674, signal_3835}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4258 ( .a ({signal_7676, signal_4342}), .b ({signal_7677, signal_3834}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4259 ( .a ({signal_7679, signal_4341}), .b ({signal_7680, signal_3833}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4260 ( .a ({signal_7682, signal_4340}), .b ({signal_7683, signal_3832}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4261 ( .a ({signal_7685, signal_4339}), .b ({signal_7686, signal_3831}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4262 ( .a ({signal_7688, signal_4375}), .b ({signal_7689, signal_3867}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4263 ( .a ({signal_7691, signal_4338}), .b ({signal_7692, signal_3830}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4264 ( .a ({signal_7694, signal_4337}), .b ({signal_7695, signal_3829}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4265 ( .a ({signal_7697, signal_4336}), .b ({signal_7698, signal_3828}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4266 ( .a ({signal_7700, signal_4335}), .b ({signal_7701, signal_3827}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4267 ( .a ({signal_7703, signal_4334}), .b ({signal_7704, signal_3826}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4268 ( .a ({signal_7706, signal_4333}), .b ({signal_7707, signal_3825}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4269 ( .a ({signal_7709, signal_4332}), .b ({signal_7710, signal_3824}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4270 ( .a ({signal_7712, signal_4331}), .b ({signal_7713, signal_3823}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4271 ( .a ({signal_7715, signal_4330}), .b ({signal_7716, signal_3822}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4272 ( .a ({signal_7718, signal_4329}), .b ({signal_7719, signal_3821}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4273 ( .a ({signal_7721, signal_4374}), .b ({signal_7722, signal_3866}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4274 ( .a ({signal_7724, signal_4328}), .b ({signal_7725, signal_3820}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4275 ( .a ({signal_7727, signal_4327}), .b ({signal_7728, signal_3819}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4276 ( .a ({signal_7730, signal_4326}), .b ({signal_7731, signal_3818}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4277 ( .a ({signal_7733, signal_4325}), .b ({signal_7734, signal_3817}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4278 ( .a ({signal_7736, signal_4324}), .b ({signal_7737, signal_3816}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4279 ( .a ({signal_7739, signal_4323}), .b ({signal_7740, signal_3815}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4280 ( .a ({signal_7742, signal_4373}), .b ({signal_7743, signal_3865}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4281 ( .a ({signal_7745, signal_4314}), .b ({signal_7746, signal_3806}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4282 ( .a ({signal_7748, signal_4313}), .b ({signal_7749, signal_3805}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4283 ( .a ({signal_7751, signal_4312}), .b ({signal_7752, signal_3804}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4284 ( .a ({signal_7754, signal_4311}), .b ({signal_7755, signal_3803}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4285 ( .a ({signal_7757, signal_4310}), .b ({signal_7758, signal_3802}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4286 ( .a ({signal_7760, signal_4309}), .b ({signal_7761, signal_3801}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4287 ( .a ({signal_7763, signal_4372}), .b ({signal_7764, signal_3864}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4288 ( .a ({signal_7766, signal_4308}), .b ({signal_7767, signal_3800}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4289 ( .a ({signal_7769, signal_4307}), .b ({signal_7770, signal_3799}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4290 ( .a ({signal_7772, signal_4306}), .b ({signal_7773, signal_3798}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4291 ( .a ({signal_7775, signal_4305}), .b ({signal_7776, signal_3797}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4292 ( .a ({signal_7778, signal_4304}), .b ({signal_7779, signal_3796}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4293 ( .a ({signal_7781, signal_4303}), .b ({signal_7782, signal_3795}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4294 ( .a ({signal_7784, signal_4302}), .b ({signal_7785, signal_3794}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4295 ( .a ({signal_7787, signal_4301}), .b ({signal_7788, signal_3793}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4296 ( .a ({signal_7790, signal_4300}), .b ({signal_7791, signal_3792}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4297 ( .a ({signal_7793, signal_4299}), .b ({signal_7794, signal_3791}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4298 ( .a ({signal_7796, signal_4371}), .b ({signal_7797, signal_3863}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4299 ( .a ({signal_7799, signal_4298}), .b ({signal_7800, signal_3790}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4300 ( .a ({signal_7802, signal_4297}), .b ({signal_7803, signal_3789}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4301 ( .a ({signal_7805, signal_4296}), .b ({signal_7806, signal_3788}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4302 ( .a ({signal_7808, signal_4295}), .b ({signal_7809, signal_3787}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4303 ( .a ({signal_7811, signal_4294}), .b ({signal_7812, signal_3786}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4304 ( .a ({signal_7814, signal_4293}), .b ({signal_7815, signal_3785}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4305 ( .a ({signal_7817, signal_4292}), .b ({signal_7818, signal_3784}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4306 ( .a ({signal_7820, signal_4291}), .b ({signal_7821, signal_3783}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4307 ( .a ({signal_7823, signal_4370}), .b ({signal_7824, signal_3862}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4308 ( .a ({signal_7826, signal_4282}), .b ({signal_7827, signal_3774}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4309 ( .a ({signal_7829, signal_4281}), .b ({signal_7830, signal_3773}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4310 ( .a ({signal_7832, signal_4280}), .b ({signal_7833, signal_3772}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4311 ( .a ({signal_7835, signal_4279}), .b ({signal_7836, signal_3771}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4312 ( .a ({signal_7838, signal_4369}), .b ({signal_7839, signal_3861}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4313 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7881, signal_4549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4314 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7882, signal_4550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4315 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7883, signal_4551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4316 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_7884, signal_4552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4317 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_7885, signal_4553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4318 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_7886, signal_4554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4319 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_7887, signal_4555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4320 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_7888, signal_4556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4321 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_7889, signal_4557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4322 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_7890, signal_4558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4323 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7891, signal_4559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4324 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7892, signal_4560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4325 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7893, signal_4561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4326 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_7894, signal_4562}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4327 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_7895, signal_4563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4328 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_7896, signal_4564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4329 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_7897, signal_4565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4330 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_7898, signal_4566}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4331 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_7899, signal_4567}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4332 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_7900, signal_4568}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4333 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7901, signal_4569}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4334 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7902, signal_4570}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4335 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7903, signal_4571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4336 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_7904, signal_4572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4337 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_7905, signal_4573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4338 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_7906, signal_4574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4339 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_7907, signal_4575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4340 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_7908, signal_4576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4341 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_7909, signal_4577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4342 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_7910, signal_4578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4343 ( .a ({signal_7634, signal_4355}), .b ({signal_7625, signal_4358}), .c ({signal_7841, signal_4579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4344 ( .a ({signal_7634, signal_4355}), .b ({signal_7616, signal_4360}), .c ({signal_7842, signal_4580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4345 ( .a ({signal_7634, signal_4355}), .b ({signal_7613, signal_4361}), .c ({signal_7843, signal_4581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4346 ( .a ({signal_7625, signal_4358}), .b ({signal_7616, signal_4360}), .c ({signal_7844, signal_4582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4347 ( .a ({signal_7619, signal_4359}), .b ({signal_7613, signal_4361}), .c ({signal_7845, signal_4583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4348 ( .a ({signal_7631, signal_4356}), .b ({signal_7628, signal_4357}), .c ({signal_7846, signal_4584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4349 ( .a ({signal_7631, signal_4356}), .b ({signal_7616, signal_4360}), .c ({signal_7847, signal_4585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4350 ( .a ({signal_7628, signal_4357}), .b ({signal_7616, signal_4360}), .c ({signal_7848, signal_4586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4351 ( .a ({signal_7625, signal_4358}), .b ({signal_7610, signal_4362}), .c ({signal_7849, signal_4587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4352 ( .a ({signal_7613, signal_4361}), .b ({signal_7610, signal_4362}), .c ({signal_7850, signal_4588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4353 ( .a ({signal_7607, signal_4363}), .b ({signal_7598, signal_4366}), .c ({signal_7851, signal_4589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4354 ( .a ({signal_7607, signal_4363}), .b ({signal_7562, signal_4368}), .c ({signal_7852, signal_4590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4355 ( .a ({signal_7607, signal_4363}), .b ({signal_7838, signal_4369}), .c ({signal_7853, signal_4591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4356 ( .a ({signal_7598, signal_4366}), .b ({signal_7562, signal_4368}), .c ({signal_7854, signal_4592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4357 ( .a ({signal_7595, signal_4367}), .b ({signal_7838, signal_4369}), .c ({signal_7855, signal_4593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4358 ( .a ({signal_7604, signal_4364}), .b ({signal_7601, signal_4365}), .c ({signal_7856, signal_4594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4359 ( .a ({signal_7604, signal_4364}), .b ({signal_7562, signal_4368}), .c ({signal_7857, signal_4595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4360 ( .a ({signal_7601, signal_4365}), .b ({signal_7562, signal_4368}), .c ({signal_7858, signal_4596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4361 ( .a ({signal_7598, signal_4366}), .b ({signal_7823, signal_4370}), .c ({signal_7859, signal_4597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4362 ( .a ({signal_7838, signal_4369}), .b ({signal_7823, signal_4370}), .c ({signal_7860, signal_4598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4363 ( .a ({signal_7796, signal_4371}), .b ({signal_7721, signal_4374}), .c ({signal_7861, signal_4599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4364 ( .a ({signal_7796, signal_4371}), .b ({signal_7655, signal_4376}), .c ({signal_7862, signal_4600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4365 ( .a ({signal_7796, signal_4371}), .b ({signal_7622, signal_4377}), .c ({signal_7863, signal_4601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4366 ( .a ({signal_7721, signal_4374}), .b ({signal_7655, signal_4376}), .c ({signal_7864, signal_4602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4367 ( .a ({signal_7688, signal_4375}), .b ({signal_7622, signal_4377}), .c ({signal_7865, signal_4603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4368 ( .a ({signal_7763, signal_4372}), .b ({signal_7742, signal_4373}), .c ({signal_7866, signal_4604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4369 ( .a ({signal_7763, signal_4372}), .b ({signal_7655, signal_4376}), .c ({signal_7867, signal_4605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4370 ( .a ({signal_7742, signal_4373}), .b ({signal_7655, signal_4376}), .c ({signal_7868, signal_4606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4371 ( .a ({signal_7721, signal_4374}), .b ({signal_7529, signal_4378}), .c ({signal_7869, signal_4607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4372 ( .a ({signal_7622, signal_4377}), .b ({signal_7529, signal_4378}), .c ({signal_7870, signal_4608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4373 ( .a ({signal_7661, signal_4347}), .b ({signal_7649, signal_4350}), .c ({signal_7871, signal_4609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4374 ( .a ({signal_7661, signal_4347}), .b ({signal_7643, signal_4352}), .c ({signal_7872, signal_4610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4375 ( .a ({signal_7661, signal_4347}), .b ({signal_7640, signal_4353}), .c ({signal_7873, signal_4611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4376 ( .a ({signal_7649, signal_4350}), .b ({signal_7643, signal_4352}), .c ({signal_7874, signal_4612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4377 ( .a ({signal_7646, signal_4351}), .b ({signal_7640, signal_4353}), .c ({signal_7875, signal_4613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4378 ( .a ({signal_7658, signal_4348}), .b ({signal_7652, signal_4349}), .c ({signal_7876, signal_4614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4379 ( .a ({signal_7658, signal_4348}), .b ({signal_7643, signal_4352}), .c ({signal_7877, signal_4615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4380 ( .a ({signal_7652, signal_4349}), .b ({signal_7643, signal_4352}), .c ({signal_7878, signal_4616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4381 ( .a ({signal_7649, signal_4350}), .b ({signal_7637, signal_4354}), .c ({signal_7879, signal_4617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4382 ( .a ({signal_7640, signal_4353}), .b ({signal_7637, signal_4354}), .c ({signal_7880, signal_4618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4383 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7911, signal_4619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4384 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7912, signal_4620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4385 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7913, signal_4621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4386 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_7914, signal_4622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4387 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_7915, signal_4623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4388 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_7916, signal_4624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4389 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_7917, signal_4625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4390 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_7918, signal_4626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4391 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_7919, signal_4627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4392 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_7920, signal_4628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4393 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_7921, signal_4629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4394 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_7922, signal_4630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4395 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7923, signal_4631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4396 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_7924, signal_4632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4397 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7925, signal_4633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4398 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_7926, signal_4634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4399 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_7927, signal_4635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4400 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_7928, signal_4636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4401 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_7929, signal_4637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4402 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7930, signal_4638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4403 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7931, signal_4639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4404 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7932, signal_4640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4405 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7933, signal_4641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4406 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_7934, signal_4642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4407 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_7935, signal_4643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4408 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_7936, signal_4644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4409 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_7937, signal_4645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4410 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_7938, signal_4646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4411 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_7939, signal_4647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4412 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_7940, signal_4648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4413 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7941, signal_4649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4414 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7942, signal_4650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4415 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7943, signal_4651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4416 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_7944, signal_4652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4417 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_7945, signal_4653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4418 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_7946, signal_4654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4419 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_7947, signal_4655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4420 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_7948, signal_4656}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4421 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_7949, signal_4657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4422 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_7950, signal_4658}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4423 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7951, signal_4659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4424 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7952, signal_4660}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4425 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7953, signal_4661}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4426 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_7954, signal_4662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4427 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_7955, signal_4663}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4428 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_7956, signal_4664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4429 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_7957, signal_4665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4430 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_7958, signal_4666}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4431 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_7959, signal_4667}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4432 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_7960, signal_4668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4433 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7961, signal_4669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4434 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7962, signal_4670}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4435 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7963, signal_4671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4436 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_7964, signal_4672}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4437 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_7965, signal_4673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4438 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_7966, signal_4674}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4439 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_7967, signal_4675}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4440 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_7968, signal_4676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4441 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_7969, signal_4677}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4442 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_7970, signal_4678}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4443 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7971, signal_4679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4444 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7972, signal_4680}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4445 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7973, signal_4681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4446 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_7974, signal_4682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4447 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_7975, signal_4683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4448 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_7976, signal_4684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4449 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_7977, signal_4685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4450 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_7978, signal_4686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4451 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_7979, signal_4687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4452 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_7980, signal_4688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4453 ( .a ({signal_7881, signal_4549}), .b ({signal_7885, signal_4553}), .c ({signal_8073, signal_4689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4454 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_7886, signal_4554}), .c ({signal_8074, signal_4690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4455 ( .a ({signal_7883, signal_4551}), .b ({signal_7884, signal_4552}), .c ({signal_8075, signal_4691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4456 ( .a ({signal_7885, signal_4553}), .b ({signal_7887, signal_4555}), .c ({signal_8076, signal_4692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4457 ( .a ({signal_7885, signal_4553}), .b ({signal_7888, signal_4556}), .c ({signal_8077, signal_4693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4458 ( .a ({signal_7886, signal_4554}), .b ({signal_7889, signal_4557}), .c ({signal_8078, signal_4694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4459 ( .a ({signal_7886, signal_4554}), .b ({signal_7890, signal_4558}), .c ({signal_8079, signal_4695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4460 ( .a ({signal_7881, signal_4549}), .b ({signal_7888, signal_4556}), .c ({signal_8080, signal_4696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4461 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7981, signal_4697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4462 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7982, signal_4698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4463 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7983, signal_4699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4464 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_7984, signal_4700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4465 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_7985, signal_4701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4466 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_7986, signal_4702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4467 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_7987, signal_4703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4468 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_7988, signal_4704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4469 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_7989, signal_4705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4470 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_7990, signal_4706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4471 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7991, signal_4707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4472 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7992, signal_4708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4473 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7993, signal_4709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4474 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_7994, signal_4710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4475 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_7995, signal_4711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4476 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_7996, signal_4712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4477 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_7997, signal_4713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4478 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_7998, signal_4714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4479 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_7999, signal_4715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4480 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_8000, signal_4716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4481 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8001, signal_4717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4482 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8002, signal_4718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4483 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8003, signal_4719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4484 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_8004, signal_4720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4485 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_8005, signal_4721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4486 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_8006, signal_4722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4487 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_8007, signal_4723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4488 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_8008, signal_4724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4489 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_8009, signal_4725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4490 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_8010, signal_4726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4491 ( .a ({signal_7891, signal_4559}), .b ({signal_7895, signal_4563}), .c ({signal_8081, signal_4727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4492 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_7896, signal_4564}), .c ({signal_8082, signal_4728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4493 ( .a ({signal_7893, signal_4561}), .b ({signal_7894, signal_4562}), .c ({signal_8083, signal_4729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4494 ( .a ({signal_7895, signal_4563}), .b ({signal_7897, signal_4565}), .c ({signal_8084, signal_4730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4495 ( .a ({signal_7895, signal_4563}), .b ({signal_7898, signal_4566}), .c ({signal_8085, signal_4731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4496 ( .a ({signal_7896, signal_4564}), .b ({signal_7899, signal_4567}), .c ({signal_8086, signal_4732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4497 ( .a ({signal_7896, signal_4564}), .b ({signal_7900, signal_4568}), .c ({signal_8087, signal_4733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4498 ( .a ({signal_7891, signal_4559}), .b ({signal_7898, signal_4566}), .c ({signal_8088, signal_4734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4499 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_8011, signal_4735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4500 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8012, signal_4736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4501 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_8013, signal_4737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4502 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8014, signal_4738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4503 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_8015, signal_4739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4504 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_8016, signal_4740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4505 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8017, signal_4741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4506 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8018, signal_4742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4507 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_8019, signal_4743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4508 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_8020, signal_4744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4509 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8021, signal_4745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4510 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8022, signal_4746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4511 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8023, signal_4747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4512 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_8024, signal_4748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4513 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_8025, signal_4749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4514 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_8026, signal_4750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4515 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_8027, signal_4751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4516 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_8028, signal_4752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4517 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_8029, signal_4753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4518 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_8030, signal_4754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4519 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8031, signal_4755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4520 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8032, signal_4756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4521 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8033, signal_4757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4522 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_8034, signal_4758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4523 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_8035, signal_4759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4524 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_8036, signal_4760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4525 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_8037, signal_4761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4526 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_8038, signal_4762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4527 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_8039, signal_4763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4528 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_8040, signal_4764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4529 ( .a ({signal_7901, signal_4569}), .b ({signal_7905, signal_4573}), .c ({signal_8089, signal_4765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4530 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_7906, signal_4574}), .c ({signal_8090, signal_4766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4531 ( .a ({signal_7903, signal_4571}), .b ({signal_7904, signal_4572}), .c ({signal_8091, signal_4767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4532 ( .a ({signal_7905, signal_4573}), .b ({signal_7907, signal_4575}), .c ({signal_8092, signal_4768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4533 ( .a ({signal_7905, signal_4573}), .b ({signal_7908, signal_4576}), .c ({signal_8093, signal_4769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4534 ( .a ({signal_7906, signal_4574}), .b ({signal_7909, signal_4577}), .c ({signal_8094, signal_4770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4535 ( .a ({signal_7906, signal_4574}), .b ({signal_7910, signal_4578}), .c ({signal_8095, signal_4771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4536 ( .a ({signal_7901, signal_4569}), .b ({signal_7908, signal_4576}), .c ({signal_8096, signal_4772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4537 ( .a ({signal_7841, signal_4579}), .b ({signal_7845, signal_4583}), .c ({signal_8041, signal_4773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4538 ( .a ({signal_7610, signal_4362}), .b ({signal_7846, signal_4584}), .c ({signal_8042, signal_4774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4539 ( .a ({signal_7843, signal_4581}), .b ({signal_7844, signal_4582}), .c ({signal_8043, signal_4775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4540 ( .a ({signal_7845, signal_4583}), .b ({signal_7847, signal_4585}), .c ({signal_8044, signal_4776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4541 ( .a ({signal_7845, signal_4583}), .b ({signal_7848, signal_4586}), .c ({signal_8045, signal_4777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4542 ( .a ({signal_7846, signal_4584}), .b ({signal_7849, signal_4587}), .c ({signal_8046, signal_4778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4543 ( .a ({signal_7846, signal_4584}), .b ({signal_7850, signal_4588}), .c ({signal_8047, signal_4779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4544 ( .a ({signal_7841, signal_4579}), .b ({signal_7848, signal_4586}), .c ({signal_8048, signal_4780}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4545 ( .a ({signal_7851, signal_4589}), .b ({signal_7855, signal_4593}), .c ({signal_8049, signal_4781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4546 ( .a ({signal_7823, signal_4370}), .b ({signal_7856, signal_4594}), .c ({signal_8050, signal_4782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4547 ( .a ({signal_7853, signal_4591}), .b ({signal_7854, signal_4592}), .c ({signal_8051, signal_4783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4548 ( .a ({signal_7855, signal_4593}), .b ({signal_7857, signal_4595}), .c ({signal_8052, signal_4784}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4549 ( .a ({signal_7855, signal_4593}), .b ({signal_7858, signal_4596}), .c ({signal_8053, signal_4785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4550 ( .a ({signal_7856, signal_4594}), .b ({signal_7859, signal_4597}), .c ({signal_8054, signal_4786}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4551 ( .a ({signal_7856, signal_4594}), .b ({signal_7860, signal_4598}), .c ({signal_8055, signal_4787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4552 ( .a ({signal_7851, signal_4589}), .b ({signal_7858, signal_4596}), .c ({signal_8056, signal_4788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4553 ( .a ({signal_7861, signal_4599}), .b ({signal_7865, signal_4603}), .c ({signal_8057, signal_4789}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4554 ( .a ({signal_7529, signal_4378}), .b ({signal_7866, signal_4604}), .c ({signal_8058, signal_4790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4555 ( .a ({signal_7863, signal_4601}), .b ({signal_7864, signal_4602}), .c ({signal_8059, signal_4791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4556 ( .a ({signal_7865, signal_4603}), .b ({signal_7867, signal_4605}), .c ({signal_8060, signal_4792}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4557 ( .a ({signal_7865, signal_4603}), .b ({signal_7868, signal_4606}), .c ({signal_8061, signal_4793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4558 ( .a ({signal_7866, signal_4604}), .b ({signal_7869, signal_4607}), .c ({signal_8062, signal_4794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4559 ( .a ({signal_7866, signal_4604}), .b ({signal_7870, signal_4608}), .c ({signal_8063, signal_4795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4560 ( .a ({signal_7861, signal_4599}), .b ({signal_7868, signal_4606}), .c ({signal_8064, signal_4796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4561 ( .a ({signal_7871, signal_4609}), .b ({signal_7875, signal_4613}), .c ({signal_8065, signal_4797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4562 ( .a ({signal_7637, signal_4354}), .b ({signal_7876, signal_4614}), .c ({signal_8066, signal_4798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4563 ( .a ({signal_7873, signal_4611}), .b ({signal_7874, signal_4612}), .c ({signal_8067, signal_4799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4564 ( .a ({signal_7875, signal_4613}), .b ({signal_7877, signal_4615}), .c ({signal_8068, signal_4800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4565 ( .a ({signal_7875, signal_4613}), .b ({signal_7878, signal_4616}), .c ({signal_8069, signal_4801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4566 ( .a ({signal_7876, signal_4614}), .b ({signal_7879, signal_4617}), .c ({signal_8070, signal_4802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4567 ( .a ({signal_7876, signal_4614}), .b ({signal_7880, signal_4618}), .c ({signal_8071, signal_4803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4568 ( .a ({signal_7871, signal_4609}), .b ({signal_7878, signal_4616}), .c ({signal_8072, signal_4804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4611 ( .a ({signal_7911, signal_4619}), .b ({signal_7915, signal_4623}), .c ({signal_8121, signal_4847}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4612 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_7916, signal_4624}), .c ({signal_8122, signal_4848}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4613 ( .a ({signal_7913, signal_4621}), .b ({signal_7914, signal_4622}), .c ({signal_8123, signal_4849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4614 ( .a ({signal_7915, signal_4623}), .b ({signal_7917, signal_4625}), .c ({signal_8124, signal_4850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4615 ( .a ({signal_7915, signal_4623}), .b ({signal_7918, signal_4626}), .c ({signal_8125, signal_4851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4616 ( .a ({signal_7916, signal_4624}), .b ({signal_7919, signal_4627}), .c ({signal_8126, signal_4852}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4617 ( .a ({signal_7916, signal_4624}), .b ({signal_7920, signal_4628}), .c ({signal_8127, signal_4853}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4618 ( .a ({signal_7911, signal_4619}), .b ({signal_7918, signal_4626}), .c ({signal_8128, signal_4854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4619 ( .a ({signal_7921, signal_4629}), .b ({signal_7925, signal_4633}), .c ({signal_8129, signal_4855}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4620 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_7926, signal_4634}), .c ({signal_8130, signal_4856}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4621 ( .a ({signal_7923, signal_4631}), .b ({signal_7924, signal_4632}), .c ({signal_8131, signal_4857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4622 ( .a ({signal_7925, signal_4633}), .b ({signal_7927, signal_4635}), .c ({signal_8132, signal_4858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4623 ( .a ({signal_7925, signal_4633}), .b ({signal_7928, signal_4636}), .c ({signal_8133, signal_4859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4624 ( .a ({signal_7926, signal_4634}), .b ({signal_7929, signal_4637}), .c ({signal_8134, signal_4860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4625 ( .a ({signal_7926, signal_4634}), .b ({signal_7930, signal_4638}), .c ({signal_8135, signal_4861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4626 ( .a ({signal_7921, signal_4629}), .b ({signal_7928, signal_4636}), .c ({signal_8136, signal_4862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4627 ( .a ({signal_7931, signal_4639}), .b ({signal_7935, signal_4643}), .c ({signal_8137, signal_4863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4628 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_7936, signal_4644}), .c ({signal_8138, signal_4864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4629 ( .a ({signal_7933, signal_4641}), .b ({signal_7934, signal_4642}), .c ({signal_8139, signal_4865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4630 ( .a ({signal_7935, signal_4643}), .b ({signal_7937, signal_4645}), .c ({signal_8140, signal_4866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4631 ( .a ({signal_7935, signal_4643}), .b ({signal_7938, signal_4646}), .c ({signal_8141, signal_4867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4632 ( .a ({signal_7936, signal_4644}), .b ({signal_7939, signal_4647}), .c ({signal_8142, signal_4868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4633 ( .a ({signal_7936, signal_4644}), .b ({signal_7940, signal_4648}), .c ({signal_8143, signal_4869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4634 ( .a ({signal_7931, signal_4639}), .b ({signal_7938, signal_4646}), .c ({signal_8144, signal_4870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4635 ( .a ({signal_7941, signal_4649}), .b ({signal_7945, signal_4653}), .c ({signal_8145, signal_4871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4636 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_7946, signal_4654}), .c ({signal_8146, signal_4872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4637 ( .a ({signal_7943, signal_4651}), .b ({signal_7944, signal_4652}), .c ({signal_8147, signal_4873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4638 ( .a ({signal_7945, signal_4653}), .b ({signal_7947, signal_4655}), .c ({signal_8148, signal_4874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4639 ( .a ({signal_7945, signal_4653}), .b ({signal_7948, signal_4656}), .c ({signal_8149, signal_4875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4640 ( .a ({signal_7946, signal_4654}), .b ({signal_7949, signal_4657}), .c ({signal_8150, signal_4876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4641 ( .a ({signal_7946, signal_4654}), .b ({signal_7950, signal_4658}), .c ({signal_8151, signal_4877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4642 ( .a ({signal_7941, signal_4649}), .b ({signal_7948, signal_4656}), .c ({signal_8152, signal_4878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4643 ( .a ({signal_7951, signal_4659}), .b ({signal_7955, signal_4663}), .c ({signal_8153, signal_4879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4644 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_7956, signal_4664}), .c ({signal_8154, signal_4880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4645 ( .a ({signal_7953, signal_4661}), .b ({signal_7954, signal_4662}), .c ({signal_8155, signal_4881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4646 ( .a ({signal_7955, signal_4663}), .b ({signal_7957, signal_4665}), .c ({signal_8156, signal_4882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4647 ( .a ({signal_7955, signal_4663}), .b ({signal_7958, signal_4666}), .c ({signal_8157, signal_4883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4648 ( .a ({signal_7956, signal_4664}), .b ({signal_7959, signal_4667}), .c ({signal_8158, signal_4884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4649 ( .a ({signal_7956, signal_4664}), .b ({signal_7960, signal_4668}), .c ({signal_8159, signal_4885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4650 ( .a ({signal_7951, signal_4659}), .b ({signal_7958, signal_4666}), .c ({signal_8160, signal_4886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4651 ( .a ({signal_7961, signal_4669}), .b ({signal_7965, signal_4673}), .c ({signal_8161, signal_4887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4652 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_7966, signal_4674}), .c ({signal_8162, signal_4888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4653 ( .a ({signal_7963, signal_4671}), .b ({signal_7964, signal_4672}), .c ({signal_8163, signal_4889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4654 ( .a ({signal_7965, signal_4673}), .b ({signal_7967, signal_4675}), .c ({signal_8164, signal_4890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4655 ( .a ({signal_7965, signal_4673}), .b ({signal_7968, signal_4676}), .c ({signal_8165, signal_4891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4656 ( .a ({signal_7966, signal_4674}), .b ({signal_7969, signal_4677}), .c ({signal_8166, signal_4892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4657 ( .a ({signal_7966, signal_4674}), .b ({signal_7970, signal_4678}), .c ({signal_8167, signal_4893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4658 ( .a ({signal_7961, signal_4669}), .b ({signal_7968, signal_4676}), .c ({signal_8168, signal_4894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4659 ( .a ({signal_7971, signal_4679}), .b ({signal_7975, signal_4683}), .c ({signal_8169, signal_4895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4660 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_7976, signal_4684}), .c ({signal_8170, signal_4896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4661 ( .a ({signal_7973, signal_4681}), .b ({signal_7974, signal_4682}), .c ({signal_8171, signal_4897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4662 ( .a ({signal_7975, signal_4683}), .b ({signal_7977, signal_4685}), .c ({signal_8172, signal_4898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4663 ( .a ({signal_7975, signal_4683}), .b ({signal_7978, signal_4686}), .c ({signal_8173, signal_4899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4664 ( .a ({signal_7976, signal_4684}), .b ({signal_7979, signal_4687}), .c ({signal_8174, signal_4900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4665 ( .a ({signal_7976, signal_4684}), .b ({signal_7980, signal_4688}), .c ({signal_8175, signal_4901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4666 ( .a ({signal_7971, signal_4679}), .b ({signal_7978, signal_4686}), .c ({signal_8176, signal_4902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4667 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_8073, signal_4689}), .c ({signal_8271, signal_4903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4668 ( .a ({signal_7886, signal_4554}), .b ({signal_8073, signal_4689}), .c ({signal_8272, signal_4904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4669 ( .a ({signal_7887, signal_4555}), .b ({signal_8073, signal_4689}), .c ({signal_8273, signal_4905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4670 ( .a ({signal_8074, signal_4690}), .b ({signal_8077, signal_4693}), .c ({signal_8274, signal_4906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4671 ( .a ({signal_7881, signal_4549}), .b ({signal_8078, signal_4694}), .c ({signal_8275, signal_4907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4672 ( .a ({signal_7882, signal_4550}), .b ({signal_8079, signal_4695}), .c ({signal_8276, signal_4908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4673 ( .a ({signal_7883, signal_4551}), .b ({signal_8077, signal_4693}), .c ({signal_8277, signal_4909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4674 ( .a ({signal_7981, signal_4697}), .b ({signal_7985, signal_4701}), .c ({signal_8177, signal_4910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4675 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_7986, signal_4702}), .c ({signal_8178, signal_4911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4676 ( .a ({signal_7983, signal_4699}), .b ({signal_7984, signal_4700}), .c ({signal_8179, signal_4912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4677 ( .a ({signal_7985, signal_4701}), .b ({signal_7987, signal_4703}), .c ({signal_8180, signal_4913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4678 ( .a ({signal_7985, signal_4701}), .b ({signal_7988, signal_4704}), .c ({signal_8181, signal_4914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4679 ( .a ({signal_7986, signal_4702}), .b ({signal_7989, signal_4705}), .c ({signal_8182, signal_4915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4680 ( .a ({signal_7986, signal_4702}), .b ({signal_7990, signal_4706}), .c ({signal_8183, signal_4916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4681 ( .a ({signal_7981, signal_4697}), .b ({signal_7988, signal_4704}), .c ({signal_8184, signal_4917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4682 ( .a ({signal_7991, signal_4707}), .b ({signal_7995, signal_4711}), .c ({signal_8185, signal_4918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4683 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_7996, signal_4712}), .c ({signal_8186, signal_4919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4684 ( .a ({signal_7993, signal_4709}), .b ({signal_7994, signal_4710}), .c ({signal_8187, signal_4920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4685 ( .a ({signal_7995, signal_4711}), .b ({signal_7997, signal_4713}), .c ({signal_8188, signal_4921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4686 ( .a ({signal_7995, signal_4711}), .b ({signal_7998, signal_4714}), .c ({signal_8189, signal_4922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4687 ( .a ({signal_7996, signal_4712}), .b ({signal_7999, signal_4715}), .c ({signal_8190, signal_4923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4688 ( .a ({signal_7996, signal_4712}), .b ({signal_8000, signal_4716}), .c ({signal_8191, signal_4924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4689 ( .a ({signal_7991, signal_4707}), .b ({signal_7998, signal_4714}), .c ({signal_8192, signal_4925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4690 ( .a ({signal_8001, signal_4717}), .b ({signal_8005, signal_4721}), .c ({signal_8193, signal_4926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4691 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8006, signal_4722}), .c ({signal_8194, signal_4927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4692 ( .a ({signal_8003, signal_4719}), .b ({signal_8004, signal_4720}), .c ({signal_8195, signal_4928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4693 ( .a ({signal_8005, signal_4721}), .b ({signal_8007, signal_4723}), .c ({signal_8196, signal_4929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4694 ( .a ({signal_8005, signal_4721}), .b ({signal_8008, signal_4724}), .c ({signal_8197, signal_4930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4695 ( .a ({signal_8006, signal_4722}), .b ({signal_8009, signal_4725}), .c ({signal_8198, signal_4931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4696 ( .a ({signal_8006, signal_4722}), .b ({signal_8010, signal_4726}), .c ({signal_8199, signal_4932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4697 ( .a ({signal_8001, signal_4717}), .b ({signal_8008, signal_4724}), .c ({signal_8200, signal_4933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4698 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_8081, signal_4727}), .c ({signal_8278, signal_4934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4699 ( .a ({signal_7896, signal_4564}), .b ({signal_8081, signal_4727}), .c ({signal_8279, signal_4935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4700 ( .a ({signal_7897, signal_4565}), .b ({signal_8081, signal_4727}), .c ({signal_8280, signal_4936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4701 ( .a ({signal_8082, signal_4728}), .b ({signal_8085, signal_4731}), .c ({signal_8281, signal_4937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4702 ( .a ({signal_7891, signal_4559}), .b ({signal_8086, signal_4732}), .c ({signal_8282, signal_4938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4703 ( .a ({signal_7892, signal_4560}), .b ({signal_8087, signal_4733}), .c ({signal_8283, signal_4939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4704 ( .a ({signal_7893, signal_4561}), .b ({signal_8085, signal_4731}), .c ({signal_8284, signal_4940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4705 ( .a ({signal_8011, signal_4735}), .b ({signal_8015, signal_4739}), .c ({signal_8201, signal_4941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4706 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8016, signal_4740}), .c ({signal_8202, signal_4942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4707 ( .a ({signal_8013, signal_4737}), .b ({signal_8014, signal_4738}), .c ({signal_8203, signal_4943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4708 ( .a ({signal_8015, signal_4739}), .b ({signal_8017, signal_4741}), .c ({signal_8204, signal_4944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4709 ( .a ({signal_8015, signal_4739}), .b ({signal_8018, signal_4742}), .c ({signal_8205, signal_4945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4710 ( .a ({signal_8016, signal_4740}), .b ({signal_8019, signal_4743}), .c ({signal_8206, signal_4946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4711 ( .a ({signal_8016, signal_4740}), .b ({signal_8020, signal_4744}), .c ({signal_8207, signal_4947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4712 ( .a ({signal_8011, signal_4735}), .b ({signal_8018, signal_4742}), .c ({signal_8208, signal_4948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4713 ( .a ({signal_8021, signal_4745}), .b ({signal_8025, signal_4749}), .c ({signal_8209, signal_4949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4714 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8026, signal_4750}), .c ({signal_8210, signal_4950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4715 ( .a ({signal_8023, signal_4747}), .b ({signal_8024, signal_4748}), .c ({signal_8211, signal_4951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4716 ( .a ({signal_8025, signal_4749}), .b ({signal_8027, signal_4751}), .c ({signal_8212, signal_4952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4717 ( .a ({signal_8025, signal_4749}), .b ({signal_8028, signal_4752}), .c ({signal_8213, signal_4953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4718 ( .a ({signal_8026, signal_4750}), .b ({signal_8029, signal_4753}), .c ({signal_8214, signal_4954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4719 ( .a ({signal_8026, signal_4750}), .b ({signal_8030, signal_4754}), .c ({signal_8215, signal_4955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4720 ( .a ({signal_8021, signal_4745}), .b ({signal_8028, signal_4752}), .c ({signal_8216, signal_4956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4721 ( .a ({signal_8031, signal_4755}), .b ({signal_8035, signal_4759}), .c ({signal_8217, signal_4957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4722 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8036, signal_4760}), .c ({signal_8218, signal_4958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4723 ( .a ({signal_8033, signal_4757}), .b ({signal_8034, signal_4758}), .c ({signal_8219, signal_4959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4724 ( .a ({signal_8035, signal_4759}), .b ({signal_8037, signal_4761}), .c ({signal_8220, signal_4960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4725 ( .a ({signal_8035, signal_4759}), .b ({signal_8038, signal_4762}), .c ({signal_8221, signal_4961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4726 ( .a ({signal_8036, signal_4760}), .b ({signal_8039, signal_4763}), .c ({signal_8222, signal_4962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4727 ( .a ({signal_8036, signal_4760}), .b ({signal_8040, signal_4764}), .c ({signal_8223, signal_4963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4728 ( .a ({signal_8031, signal_4755}), .b ({signal_8038, signal_4762}), .c ({signal_8224, signal_4964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4729 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_8089, signal_4765}), .c ({signal_8285, signal_4965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4730 ( .a ({signal_7906, signal_4574}), .b ({signal_8089, signal_4765}), .c ({signal_8286, signal_4966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4731 ( .a ({signal_7907, signal_4575}), .b ({signal_8089, signal_4765}), .c ({signal_8287, signal_4967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4732 ( .a ({signal_8090, signal_4766}), .b ({signal_8093, signal_4769}), .c ({signal_8288, signal_4968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4733 ( .a ({signal_7901, signal_4569}), .b ({signal_8094, signal_4770}), .c ({signal_8289, signal_4969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4734 ( .a ({signal_7902, signal_4570}), .b ({signal_8095, signal_4771}), .c ({signal_8290, signal_4970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4735 ( .a ({signal_7903, signal_4571}), .b ({signal_8093, signal_4769}), .c ({signal_8291, signal_4971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4736 ( .a ({signal_7610, signal_4362}), .b ({signal_8041, signal_4773}), .c ({signal_8225, signal_4972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4737 ( .a ({signal_7846, signal_4584}), .b ({signal_8041, signal_4773}), .c ({signal_8226, signal_4973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4738 ( .a ({signal_7847, signal_4585}), .b ({signal_8041, signal_4773}), .c ({signal_8227, signal_4974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4739 ( .a ({signal_8042, signal_4774}), .b ({signal_8045, signal_4777}), .c ({signal_8228, signal_4975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4740 ( .a ({signal_7841, signal_4579}), .b ({signal_8046, signal_4778}), .c ({signal_8229, signal_4976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4741 ( .a ({signal_7842, signal_4580}), .b ({signal_8047, signal_4779}), .c ({signal_8230, signal_4977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4742 ( .a ({signal_7843, signal_4581}), .b ({signal_8045, signal_4777}), .c ({signal_8231, signal_4978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4743 ( .a ({signal_7823, signal_4370}), .b ({signal_8049, signal_4781}), .c ({signal_8232, signal_4979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4744 ( .a ({signal_7856, signal_4594}), .b ({signal_8049, signal_4781}), .c ({signal_8233, signal_4980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4745 ( .a ({signal_7857, signal_4595}), .b ({signal_8049, signal_4781}), .c ({signal_8234, signal_4981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4746 ( .a ({signal_8050, signal_4782}), .b ({signal_8053, signal_4785}), .c ({signal_8235, signal_4982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4747 ( .a ({signal_7851, signal_4589}), .b ({signal_8054, signal_4786}), .c ({signal_8236, signal_4983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4748 ( .a ({signal_7852, signal_4590}), .b ({signal_8055, signal_4787}), .c ({signal_8237, signal_4984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4749 ( .a ({signal_7853, signal_4591}), .b ({signal_8053, signal_4785}), .c ({signal_8238, signal_4985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4750 ( .a ({signal_7529, signal_4378}), .b ({signal_8057, signal_4789}), .c ({signal_8239, signal_4986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4751 ( .a ({signal_7866, signal_4604}), .b ({signal_8057, signal_4789}), .c ({signal_8240, signal_4987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4752 ( .a ({signal_7867, signal_4605}), .b ({signal_8057, signal_4789}), .c ({signal_8241, signal_4988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4753 ( .a ({signal_8058, signal_4790}), .b ({signal_8061, signal_4793}), .c ({signal_8242, signal_4989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4754 ( .a ({signal_7861, signal_4599}), .b ({signal_8062, signal_4794}), .c ({signal_8243, signal_4990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4755 ( .a ({signal_7862, signal_4600}), .b ({signal_8063, signal_4795}), .c ({signal_8244, signal_4991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4756 ( .a ({signal_7863, signal_4601}), .b ({signal_8061, signal_4793}), .c ({signal_8245, signal_4992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4757 ( .a ({signal_7637, signal_4354}), .b ({signal_8065, signal_4797}), .c ({signal_8246, signal_4993}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4758 ( .a ({signal_7876, signal_4614}), .b ({signal_8065, signal_4797}), .c ({signal_8247, signal_4994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4759 ( .a ({signal_7877, signal_4615}), .b ({signal_8065, signal_4797}), .c ({signal_8248, signal_4995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4760 ( .a ({signal_8066, signal_4798}), .b ({signal_8069, signal_4801}), .c ({signal_8249, signal_4996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4761 ( .a ({signal_7871, signal_4609}), .b ({signal_8070, signal_4802}), .c ({signal_8250, signal_4997}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4762 ( .a ({signal_7872, signal_4610}), .b ({signal_8071, signal_4803}), .c ({signal_8251, signal_4998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4763 ( .a ({signal_7873, signal_4611}), .b ({signal_8069, signal_4801}), .c ({signal_8252, signal_4999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4863 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_8121, signal_4847}), .c ({signal_8382, signal_5099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4864 ( .a ({signal_7916, signal_4624}), .b ({signal_8121, signal_4847}), .c ({signal_8383, signal_5100}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4865 ( .a ({signal_7917, signal_4625}), .b ({signal_8121, signal_4847}), .c ({signal_8384, signal_5101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4866 ( .a ({signal_8122, signal_4848}), .b ({signal_8125, signal_4851}), .c ({signal_8385, signal_5102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4867 ( .a ({signal_7911, signal_4619}), .b ({signal_8126, signal_4852}), .c ({signal_8386, signal_5103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4868 ( .a ({signal_7912, signal_4620}), .b ({signal_8127, signal_4853}), .c ({signal_8387, signal_5104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4869 ( .a ({signal_7913, signal_4621}), .b ({signal_8125, signal_4851}), .c ({signal_8388, signal_5105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4870 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_8129, signal_4855}), .c ({signal_8389, signal_5106}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4871 ( .a ({signal_7926, signal_4634}), .b ({signal_8129, signal_4855}), .c ({signal_8390, signal_5107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4872 ( .a ({signal_7927, signal_4635}), .b ({signal_8129, signal_4855}), .c ({signal_8391, signal_5108}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4873 ( .a ({signal_8130, signal_4856}), .b ({signal_8133, signal_4859}), .c ({signal_8392, signal_5109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4874 ( .a ({signal_7921, signal_4629}), .b ({signal_8134, signal_4860}), .c ({signal_8393, signal_5110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4875 ( .a ({signal_7922, signal_4630}), .b ({signal_8135, signal_4861}), .c ({signal_8394, signal_5111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4876 ( .a ({signal_7923, signal_4631}), .b ({signal_8133, signal_4859}), .c ({signal_8395, signal_5112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4877 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_8137, signal_4863}), .c ({signal_8396, signal_5113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4878 ( .a ({signal_7936, signal_4644}), .b ({signal_8137, signal_4863}), .c ({signal_8397, signal_5114}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4879 ( .a ({signal_7937, signal_4645}), .b ({signal_8137, signal_4863}), .c ({signal_8398, signal_5115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4880 ( .a ({signal_8138, signal_4864}), .b ({signal_8141, signal_4867}), .c ({signal_8399, signal_5116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4881 ( .a ({signal_7931, signal_4639}), .b ({signal_8142, signal_4868}), .c ({signal_8400, signal_5117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4882 ( .a ({signal_7932, signal_4640}), .b ({signal_8143, signal_4869}), .c ({signal_8401, signal_5118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4883 ( .a ({signal_7933, signal_4641}), .b ({signal_8141, signal_4867}), .c ({signal_8402, signal_5119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4884 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_8145, signal_4871}), .c ({signal_8403, signal_5120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4885 ( .a ({signal_7946, signal_4654}), .b ({signal_8145, signal_4871}), .c ({signal_8404, signal_5121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4886 ( .a ({signal_7947, signal_4655}), .b ({signal_8145, signal_4871}), .c ({signal_8405, signal_5122}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4887 ( .a ({signal_8146, signal_4872}), .b ({signal_8149, signal_4875}), .c ({signal_8406, signal_5123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4888 ( .a ({signal_7941, signal_4649}), .b ({signal_8150, signal_4876}), .c ({signal_8407, signal_5124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4889 ( .a ({signal_7942, signal_4650}), .b ({signal_8151, signal_4877}), .c ({signal_8408, signal_5125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4890 ( .a ({signal_7943, signal_4651}), .b ({signal_8149, signal_4875}), .c ({signal_8409, signal_5126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4891 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_8153, signal_4879}), .c ({signal_8410, signal_5127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4892 ( .a ({signal_7956, signal_4664}), .b ({signal_8153, signal_4879}), .c ({signal_8411, signal_5128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4893 ( .a ({signal_7957, signal_4665}), .b ({signal_8153, signal_4879}), .c ({signal_8412, signal_5129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4894 ( .a ({signal_8154, signal_4880}), .b ({signal_8157, signal_4883}), .c ({signal_8413, signal_5130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4895 ( .a ({signal_7951, signal_4659}), .b ({signal_8158, signal_4884}), .c ({signal_8414, signal_5131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4896 ( .a ({signal_7952, signal_4660}), .b ({signal_8159, signal_4885}), .c ({signal_8415, signal_5132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4897 ( .a ({signal_7953, signal_4661}), .b ({signal_8157, signal_4883}), .c ({signal_8416, signal_5133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4898 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_8161, signal_4887}), .c ({signal_8417, signal_5134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4899 ( .a ({signal_7966, signal_4674}), .b ({signal_8161, signal_4887}), .c ({signal_8418, signal_5135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4900 ( .a ({signal_7967, signal_4675}), .b ({signal_8161, signal_4887}), .c ({signal_8419, signal_5136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4901 ( .a ({signal_8162, signal_4888}), .b ({signal_8165, signal_4891}), .c ({signal_8420, signal_5137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4902 ( .a ({signal_7961, signal_4669}), .b ({signal_8166, signal_4892}), .c ({signal_8421, signal_5138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4903 ( .a ({signal_7962, signal_4670}), .b ({signal_8167, signal_4893}), .c ({signal_8422, signal_5139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4904 ( .a ({signal_7963, signal_4671}), .b ({signal_8165, signal_4891}), .c ({signal_8423, signal_5140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4905 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_8169, signal_4895}), .c ({signal_8424, signal_5141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4906 ( .a ({signal_7976, signal_4684}), .b ({signal_8169, signal_4895}), .c ({signal_8425, signal_5142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4907 ( .a ({signal_7977, signal_4685}), .b ({signal_8169, signal_4895}), .c ({signal_8426, signal_5143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4908 ( .a ({signal_8170, signal_4896}), .b ({signal_8173, signal_4899}), .c ({signal_8427, signal_5144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4909 ( .a ({signal_7971, signal_4679}), .b ({signal_8174, signal_4900}), .c ({signal_8428, signal_5145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4910 ( .a ({signal_7972, signal_4680}), .b ({signal_8175, signal_4901}), .c ({signal_8429, signal_5146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4911 ( .a ({signal_7973, signal_4681}), .b ({signal_8173, signal_4899}), .c ({signal_8430, signal_5147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4912 ( .a ({signal_7882, signal_4550}), .b ({signal_8272, signal_4904}), .c ({signal_8506, signal_5148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4913 ( .a ({signal_8274, signal_4906}), .b ({signal_8275, signal_4907}), .c ({signal_8507, signal_5149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4918 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_8177, signal_4910}), .c ({signal_8431, signal_5154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4919 ( .a ({signal_7986, signal_4702}), .b ({signal_8177, signal_4910}), .c ({signal_8432, signal_5155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4920 ( .a ({signal_7987, signal_4703}), .b ({signal_8177, signal_4910}), .c ({signal_8433, signal_5156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4921 ( .a ({signal_8178, signal_4911}), .b ({signal_8181, signal_4914}), .c ({signal_8434, signal_5157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4922 ( .a ({signal_7981, signal_4697}), .b ({signal_8182, signal_4915}), .c ({signal_8435, signal_5158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4923 ( .a ({signal_7982, signal_4698}), .b ({signal_8183, signal_4916}), .c ({signal_8436, signal_5159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4924 ( .a ({signal_7983, signal_4699}), .b ({signal_8181, signal_4914}), .c ({signal_8437, signal_5160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4925 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_8185, signal_4918}), .c ({signal_8438, signal_5161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4926 ( .a ({signal_7996, signal_4712}), .b ({signal_8185, signal_4918}), .c ({signal_8439, signal_5162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4927 ( .a ({signal_7997, signal_4713}), .b ({signal_8185, signal_4918}), .c ({signal_8440, signal_5163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4928 ( .a ({signal_8186, signal_4919}), .b ({signal_8189, signal_4922}), .c ({signal_8441, signal_5164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4929 ( .a ({signal_7991, signal_4707}), .b ({signal_8190, signal_4923}), .c ({signal_8442, signal_5165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4930 ( .a ({signal_7992, signal_4708}), .b ({signal_8191, signal_4924}), .c ({signal_8443, signal_5166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4931 ( .a ({signal_7993, signal_4709}), .b ({signal_8189, signal_4922}), .c ({signal_8444, signal_5167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4932 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8193, signal_4926}), .c ({signal_8445, signal_5168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4933 ( .a ({signal_8006, signal_4722}), .b ({signal_8193, signal_4926}), .c ({signal_8446, signal_5169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4934 ( .a ({signal_8007, signal_4723}), .b ({signal_8193, signal_4926}), .c ({signal_8447, signal_5170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4935 ( .a ({signal_8194, signal_4927}), .b ({signal_8197, signal_4930}), .c ({signal_8448, signal_5171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4936 ( .a ({signal_8001, signal_4717}), .b ({signal_8198, signal_4931}), .c ({signal_8449, signal_5172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4937 ( .a ({signal_8002, signal_4718}), .b ({signal_8199, signal_4932}), .c ({signal_8450, signal_5173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4938 ( .a ({signal_8003, signal_4719}), .b ({signal_8197, signal_4930}), .c ({signal_8451, signal_5174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4939 ( .a ({signal_7892, signal_4560}), .b ({signal_8279, signal_4935}), .c ({signal_8512, signal_5175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4940 ( .a ({signal_8281, signal_4937}), .b ({signal_8282, signal_4938}), .c ({signal_8513, signal_5176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4945 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8201, signal_4941}), .c ({signal_8452, signal_5181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4946 ( .a ({signal_8016, signal_4740}), .b ({signal_8201, signal_4941}), .c ({signal_8453, signal_5182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4947 ( .a ({signal_8017, signal_4741}), .b ({signal_8201, signal_4941}), .c ({signal_8454, signal_5183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4948 ( .a ({signal_8202, signal_4942}), .b ({signal_8205, signal_4945}), .c ({signal_8455, signal_5184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4949 ( .a ({signal_8011, signal_4735}), .b ({signal_8206, signal_4946}), .c ({signal_8456, signal_5185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4950 ( .a ({signal_8012, signal_4736}), .b ({signal_8207, signal_4947}), .c ({signal_8457, signal_5186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4951 ( .a ({signal_8013, signal_4737}), .b ({signal_8205, signal_4945}), .c ({signal_8458, signal_5187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4952 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8209, signal_4949}), .c ({signal_8459, signal_5188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4953 ( .a ({signal_8026, signal_4750}), .b ({signal_8209, signal_4949}), .c ({signal_8460, signal_5189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4954 ( .a ({signal_8027, signal_4751}), .b ({signal_8209, signal_4949}), .c ({signal_8461, signal_5190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4955 ( .a ({signal_8210, signal_4950}), .b ({signal_8213, signal_4953}), .c ({signal_8462, signal_5191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4956 ( .a ({signal_8021, signal_4745}), .b ({signal_8214, signal_4954}), .c ({signal_8463, signal_5192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4957 ( .a ({signal_8022, signal_4746}), .b ({signal_8215, signal_4955}), .c ({signal_8464, signal_5193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4958 ( .a ({signal_8023, signal_4747}), .b ({signal_8213, signal_4953}), .c ({signal_8465, signal_5194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4959 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8217, signal_4957}), .c ({signal_8466, signal_5195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4960 ( .a ({signal_8036, signal_4760}), .b ({signal_8217, signal_4957}), .c ({signal_8467, signal_5196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4961 ( .a ({signal_8037, signal_4761}), .b ({signal_8217, signal_4957}), .c ({signal_8468, signal_5197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4962 ( .a ({signal_8218, signal_4958}), .b ({signal_8221, signal_4961}), .c ({signal_8469, signal_5198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4963 ( .a ({signal_8031, signal_4755}), .b ({signal_8222, signal_4962}), .c ({signal_8470, signal_5199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4964 ( .a ({signal_8032, signal_4756}), .b ({signal_8223, signal_4963}), .c ({signal_8471, signal_5200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4965 ( .a ({signal_8033, signal_4757}), .b ({signal_8221, signal_4961}), .c ({signal_8472, signal_5201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4966 ( .a ({signal_7902, signal_4570}), .b ({signal_8286, signal_4966}), .c ({signal_8518, signal_5202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4967 ( .a ({signal_8288, signal_4968}), .b ({signal_8289, signal_4969}), .c ({signal_8519, signal_5203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4972 ( .a ({signal_7842, signal_4580}), .b ({signal_8226, signal_4973}), .c ({signal_8473, signal_5208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4973 ( .a ({signal_8228, signal_4975}), .b ({signal_8229, signal_4976}), .c ({signal_8474, signal_5209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4978 ( .a ({signal_7852, signal_4590}), .b ({signal_8233, signal_4980}), .c ({signal_8479, signal_5214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4979 ( .a ({signal_8235, signal_4982}), .b ({signal_8236, signal_4983}), .c ({signal_8480, signal_5215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4984 ( .a ({signal_7862, signal_4600}), .b ({signal_8240, signal_4987}), .c ({signal_8485, signal_5220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4985 ( .a ({signal_8242, signal_4989}), .b ({signal_8243, signal_4990}), .c ({signal_8486, signal_5221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4990 ( .a ({signal_7872, signal_4610}), .b ({signal_8247, signal_4994}), .c ({signal_8491, signal_5226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4991 ( .a ({signal_8249, signal_4996}), .b ({signal_8250, signal_4997}), .c ({signal_8492, signal_5227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5035 ( .a ({signal_7912, signal_4620}), .b ({signal_8383, signal_5100}), .c ({signal_8563, signal_5271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5036 ( .a ({signal_8385, signal_5102}), .b ({signal_8386, signal_5103}), .c ({signal_8564, signal_5272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5041 ( .a ({signal_7922, signal_4630}), .b ({signal_8390, signal_5107}), .c ({signal_8569, signal_5277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5042 ( .a ({signal_8392, signal_5109}), .b ({signal_8393, signal_5110}), .c ({signal_8570, signal_5278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5047 ( .a ({signal_7932, signal_4640}), .b ({signal_8397, signal_5114}), .c ({signal_8575, signal_5283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5048 ( .a ({signal_8399, signal_5116}), .b ({signal_8400, signal_5117}), .c ({signal_8576, signal_5284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5053 ( .a ({signal_7942, signal_4650}), .b ({signal_8404, signal_5121}), .c ({signal_8581, signal_5289}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5054 ( .a ({signal_8406, signal_5123}), .b ({signal_8407, signal_5124}), .c ({signal_8582, signal_5290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5059 ( .a ({signal_7952, signal_4660}), .b ({signal_8411, signal_5128}), .c ({signal_8587, signal_5295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5060 ( .a ({signal_8413, signal_5130}), .b ({signal_8414, signal_5131}), .c ({signal_8588, signal_5296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5065 ( .a ({signal_7962, signal_4670}), .b ({signal_8418, signal_5135}), .c ({signal_8593, signal_5301}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5066 ( .a ({signal_8420, signal_5137}), .b ({signal_8421, signal_5138}), .c ({signal_8594, signal_5302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5071 ( .a ({signal_7972, signal_4680}), .b ({signal_8425, signal_5142}), .c ({signal_8599, signal_5307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5072 ( .a ({signal_8427, signal_5144}), .b ({signal_8428, signal_5145}), .c ({signal_8600, signal_5308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5082 ( .a ({signal_7982, signal_4698}), .b ({signal_8432, signal_5155}), .c ({signal_8605, signal_5318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5083 ( .a ({signal_8434, signal_5157}), .b ({signal_8435, signal_5158}), .c ({signal_8606, signal_5319}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5088 ( .a ({signal_7992, signal_4708}), .b ({signal_8439, signal_5162}), .c ({signal_8611, signal_5324}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5089 ( .a ({signal_8441, signal_5164}), .b ({signal_8442, signal_5165}), .c ({signal_8612, signal_5325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5094 ( .a ({signal_8002, signal_4718}), .b ({signal_8446, signal_5169}), .c ({signal_8617, signal_5330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5095 ( .a ({signal_8448, signal_5171}), .b ({signal_8449, signal_5172}), .c ({signal_8618, signal_5331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5105 ( .a ({signal_8012, signal_4736}), .b ({signal_8453, signal_5182}), .c ({signal_8623, signal_5341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5106 ( .a ({signal_8455, signal_5184}), .b ({signal_8456, signal_5185}), .c ({signal_8624, signal_5342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5111 ( .a ({signal_8022, signal_4746}), .b ({signal_8460, signal_5189}), .c ({signal_8629, signal_5347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5112 ( .a ({signal_8462, signal_5191}), .b ({signal_8463, signal_5192}), .c ({signal_8630, signal_5348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5117 ( .a ({signal_8032, signal_4756}), .b ({signal_8467, signal_5196}), .c ({signal_8635, signal_5353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5118 ( .a ({signal_8469, signal_5198}), .b ({signal_8470, signal_5199}), .c ({signal_8636, signal_5354}) ) ;

    /* cells in depth 1 */
    buf_clk cell_7581 ( .C (clk), .D (signal_4905), .Q (signal_12469) ) ;
    buf_clk cell_7583 ( .C (clk), .D (signal_8273), .Q (signal_12471) ) ;
    buf_clk cell_7585 ( .C (clk), .D (signal_4909), .Q (signal_12473) ) ;
    buf_clk cell_7587 ( .C (clk), .D (signal_8277), .Q (signal_12475) ) ;
    buf_clk cell_7589 ( .C (clk), .D (signal_4936), .Q (signal_12477) ) ;
    buf_clk cell_7591 ( .C (clk), .D (signal_8280), .Q (signal_12479) ) ;
    buf_clk cell_7593 ( .C (clk), .D (signal_4940), .Q (signal_12481) ) ;
    buf_clk cell_7595 ( .C (clk), .D (signal_8284), .Q (signal_12483) ) ;
    buf_clk cell_7597 ( .C (clk), .D (signal_4967), .Q (signal_12485) ) ;
    buf_clk cell_7599 ( .C (clk), .D (signal_8287), .Q (signal_12487) ) ;
    buf_clk cell_7601 ( .C (clk), .D (signal_4971), .Q (signal_12489) ) ;
    buf_clk cell_7603 ( .C (clk), .D (signal_8291), .Q (signal_12491) ) ;
    buf_clk cell_7605 ( .C (clk), .D (signal_4974), .Q (signal_12493) ) ;
    buf_clk cell_7607 ( .C (clk), .D (signal_8227), .Q (signal_12495) ) ;
    buf_clk cell_7609 ( .C (clk), .D (signal_4978), .Q (signal_12497) ) ;
    buf_clk cell_7611 ( .C (clk), .D (signal_8231), .Q (signal_12499) ) ;
    buf_clk cell_7613 ( .C (clk), .D (signal_4981), .Q (signal_12501) ) ;
    buf_clk cell_7615 ( .C (clk), .D (signal_8234), .Q (signal_12503) ) ;
    buf_clk cell_7617 ( .C (clk), .D (signal_4985), .Q (signal_12505) ) ;
    buf_clk cell_7619 ( .C (clk), .D (signal_8238), .Q (signal_12507) ) ;
    buf_clk cell_7621 ( .C (clk), .D (signal_4988), .Q (signal_12509) ) ;
    buf_clk cell_7623 ( .C (clk), .D (signal_8241), .Q (signal_12511) ) ;
    buf_clk cell_7625 ( .C (clk), .D (signal_4992), .Q (signal_12513) ) ;
    buf_clk cell_7627 ( .C (clk), .D (signal_8245), .Q (signal_12515) ) ;
    buf_clk cell_7629 ( .C (clk), .D (signal_4995), .Q (signal_12517) ) ;
    buf_clk cell_7631 ( .C (clk), .D (signal_8248), .Q (signal_12519) ) ;
    buf_clk cell_7633 ( .C (clk), .D (signal_4999), .Q (signal_12521) ) ;
    buf_clk cell_7635 ( .C (clk), .D (signal_8252), .Q (signal_12523) ) ;
    buf_clk cell_7637 ( .C (clk), .D (signal_5101), .Q (signal_12525) ) ;
    buf_clk cell_7639 ( .C (clk), .D (signal_8384), .Q (signal_12527) ) ;
    buf_clk cell_7641 ( .C (clk), .D (signal_5105), .Q (signal_12529) ) ;
    buf_clk cell_7643 ( .C (clk), .D (signal_8388), .Q (signal_12531) ) ;
    buf_clk cell_7645 ( .C (clk), .D (signal_5108), .Q (signal_12533) ) ;
    buf_clk cell_7647 ( .C (clk), .D (signal_8391), .Q (signal_12535) ) ;
    buf_clk cell_7649 ( .C (clk), .D (signal_5112), .Q (signal_12537) ) ;
    buf_clk cell_7651 ( .C (clk), .D (signal_8395), .Q (signal_12539) ) ;
    buf_clk cell_7653 ( .C (clk), .D (signal_5115), .Q (signal_12541) ) ;
    buf_clk cell_7655 ( .C (clk), .D (signal_8398), .Q (signal_12543) ) ;
    buf_clk cell_7657 ( .C (clk), .D (signal_5119), .Q (signal_12545) ) ;
    buf_clk cell_7659 ( .C (clk), .D (signal_8402), .Q (signal_12547) ) ;
    buf_clk cell_7661 ( .C (clk), .D (signal_5122), .Q (signal_12549) ) ;
    buf_clk cell_7663 ( .C (clk), .D (signal_8405), .Q (signal_12551) ) ;
    buf_clk cell_7665 ( .C (clk), .D (signal_5126), .Q (signal_12553) ) ;
    buf_clk cell_7667 ( .C (clk), .D (signal_8409), .Q (signal_12555) ) ;
    buf_clk cell_7669 ( .C (clk), .D (signal_5129), .Q (signal_12557) ) ;
    buf_clk cell_7671 ( .C (clk), .D (signal_8412), .Q (signal_12559) ) ;
    buf_clk cell_7673 ( .C (clk), .D (signal_5133), .Q (signal_12561) ) ;
    buf_clk cell_7675 ( .C (clk), .D (signal_8416), .Q (signal_12563) ) ;
    buf_clk cell_7677 ( .C (clk), .D (signal_5136), .Q (signal_12565) ) ;
    buf_clk cell_7679 ( .C (clk), .D (signal_8419), .Q (signal_12567) ) ;
    buf_clk cell_7681 ( .C (clk), .D (signal_5140), .Q (signal_12569) ) ;
    buf_clk cell_7683 ( .C (clk), .D (signal_8423), .Q (signal_12571) ) ;
    buf_clk cell_7685 ( .C (clk), .D (signal_5143), .Q (signal_12573) ) ;
    buf_clk cell_7687 ( .C (clk), .D (signal_8426), .Q (signal_12575) ) ;
    buf_clk cell_7689 ( .C (clk), .D (signal_5147), .Q (signal_12577) ) ;
    buf_clk cell_7691 ( .C (clk), .D (signal_8430), .Q (signal_12579) ) ;
    buf_clk cell_7693 ( .C (clk), .D (signal_5148), .Q (signal_12581) ) ;
    buf_clk cell_7695 ( .C (clk), .D (signal_8506), .Q (signal_12583) ) ;
    buf_clk cell_7697 ( .C (clk), .D (signal_5156), .Q (signal_12585) ) ;
    buf_clk cell_7699 ( .C (clk), .D (signal_8433), .Q (signal_12587) ) ;
    buf_clk cell_7701 ( .C (clk), .D (signal_5160), .Q (signal_12589) ) ;
    buf_clk cell_7703 ( .C (clk), .D (signal_8437), .Q (signal_12591) ) ;
    buf_clk cell_7705 ( .C (clk), .D (signal_5163), .Q (signal_12593) ) ;
    buf_clk cell_7707 ( .C (clk), .D (signal_8440), .Q (signal_12595) ) ;
    buf_clk cell_7709 ( .C (clk), .D (signal_5167), .Q (signal_12597) ) ;
    buf_clk cell_7711 ( .C (clk), .D (signal_8444), .Q (signal_12599) ) ;
    buf_clk cell_7713 ( .C (clk), .D (signal_5170), .Q (signal_12601) ) ;
    buf_clk cell_7715 ( .C (clk), .D (signal_8447), .Q (signal_12603) ) ;
    buf_clk cell_7717 ( .C (clk), .D (signal_5174), .Q (signal_12605) ) ;
    buf_clk cell_7719 ( .C (clk), .D (signal_8451), .Q (signal_12607) ) ;
    buf_clk cell_7721 ( .C (clk), .D (signal_5175), .Q (signal_12609) ) ;
    buf_clk cell_7723 ( .C (clk), .D (signal_8512), .Q (signal_12611) ) ;
    buf_clk cell_7725 ( .C (clk), .D (signal_5183), .Q (signal_12613) ) ;
    buf_clk cell_7727 ( .C (clk), .D (signal_8454), .Q (signal_12615) ) ;
    buf_clk cell_7729 ( .C (clk), .D (signal_5187), .Q (signal_12617) ) ;
    buf_clk cell_7731 ( .C (clk), .D (signal_8458), .Q (signal_12619) ) ;
    buf_clk cell_7733 ( .C (clk), .D (signal_5190), .Q (signal_12621) ) ;
    buf_clk cell_7735 ( .C (clk), .D (signal_8461), .Q (signal_12623) ) ;
    buf_clk cell_7737 ( .C (clk), .D (signal_5194), .Q (signal_12625) ) ;
    buf_clk cell_7739 ( .C (clk), .D (signal_8465), .Q (signal_12627) ) ;
    buf_clk cell_7741 ( .C (clk), .D (signal_5197), .Q (signal_12629) ) ;
    buf_clk cell_7743 ( .C (clk), .D (signal_8468), .Q (signal_12631) ) ;
    buf_clk cell_7745 ( .C (clk), .D (signal_5201), .Q (signal_12633) ) ;
    buf_clk cell_7747 ( .C (clk), .D (signal_8472), .Q (signal_12635) ) ;
    buf_clk cell_7749 ( .C (clk), .D (signal_5202), .Q (signal_12637) ) ;
    buf_clk cell_7751 ( .C (clk), .D (signal_8518), .Q (signal_12639) ) ;
    buf_clk cell_7753 ( .C (clk), .D (signal_5208), .Q (signal_12641) ) ;
    buf_clk cell_7755 ( .C (clk), .D (signal_8473), .Q (signal_12643) ) ;
    buf_clk cell_7757 ( .C (clk), .D (signal_5214), .Q (signal_12645) ) ;
    buf_clk cell_7759 ( .C (clk), .D (signal_8479), .Q (signal_12647) ) ;
    buf_clk cell_7761 ( .C (clk), .D (signal_5220), .Q (signal_12649) ) ;
    buf_clk cell_7763 ( .C (clk), .D (signal_8485), .Q (signal_12651) ) ;
    buf_clk cell_7765 ( .C (clk), .D (signal_5226), .Q (signal_12653) ) ;
    buf_clk cell_7767 ( .C (clk), .D (signal_8491), .Q (signal_12655) ) ;
    buf_clk cell_7769 ( .C (clk), .D (signal_5271), .Q (signal_12657) ) ;
    buf_clk cell_7771 ( .C (clk), .D (signal_8563), .Q (signal_12659) ) ;
    buf_clk cell_7773 ( .C (clk), .D (signal_5277), .Q (signal_12661) ) ;
    buf_clk cell_7775 ( .C (clk), .D (signal_8569), .Q (signal_12663) ) ;
    buf_clk cell_7777 ( .C (clk), .D (signal_5283), .Q (signal_12665) ) ;
    buf_clk cell_7779 ( .C (clk), .D (signal_8575), .Q (signal_12667) ) ;
    buf_clk cell_7781 ( .C (clk), .D (signal_5289), .Q (signal_12669) ) ;
    buf_clk cell_7783 ( .C (clk), .D (signal_8581), .Q (signal_12671) ) ;
    buf_clk cell_7785 ( .C (clk), .D (signal_5295), .Q (signal_12673) ) ;
    buf_clk cell_7787 ( .C (clk), .D (signal_8587), .Q (signal_12675) ) ;
    buf_clk cell_7789 ( .C (clk), .D (signal_5301), .Q (signal_12677) ) ;
    buf_clk cell_7791 ( .C (clk), .D (signal_8593), .Q (signal_12679) ) ;
    buf_clk cell_7793 ( .C (clk), .D (signal_5307), .Q (signal_12681) ) ;
    buf_clk cell_7795 ( .C (clk), .D (signal_8599), .Q (signal_12683) ) ;
    buf_clk cell_7797 ( .C (clk), .D (signal_5318), .Q (signal_12685) ) ;
    buf_clk cell_7799 ( .C (clk), .D (signal_8605), .Q (signal_12687) ) ;
    buf_clk cell_7801 ( .C (clk), .D (signal_5324), .Q (signal_12689) ) ;
    buf_clk cell_7803 ( .C (clk), .D (signal_8611), .Q (signal_12691) ) ;
    buf_clk cell_7805 ( .C (clk), .D (signal_5330), .Q (signal_12693) ) ;
    buf_clk cell_7807 ( .C (clk), .D (signal_8617), .Q (signal_12695) ) ;
    buf_clk cell_7809 ( .C (clk), .D (signal_5341), .Q (signal_12697) ) ;
    buf_clk cell_7811 ( .C (clk), .D (signal_8623), .Q (signal_12699) ) ;
    buf_clk cell_7813 ( .C (clk), .D (signal_5347), .Q (signal_12701) ) ;
    buf_clk cell_7815 ( .C (clk), .D (signal_8629), .Q (signal_12703) ) ;
    buf_clk cell_7817 ( .C (clk), .D (signal_5353), .Q (signal_12705) ) ;
    buf_clk cell_7819 ( .C (clk), .D (signal_8635), .Q (signal_12707) ) ;
    buf_clk cell_7821 ( .C (clk), .D (signal_5149), .Q (signal_12709) ) ;
    buf_clk cell_7823 ( .C (clk), .D (signal_8507), .Q (signal_12711) ) ;
    buf_clk cell_7825 ( .C (clk), .D (signal_5176), .Q (signal_12713) ) ;
    buf_clk cell_7827 ( .C (clk), .D (signal_8513), .Q (signal_12715) ) ;
    buf_clk cell_7829 ( .C (clk), .D (signal_5203), .Q (signal_12717) ) ;
    buf_clk cell_7831 ( .C (clk), .D (signal_8519), .Q (signal_12719) ) ;
    buf_clk cell_7833 ( .C (clk), .D (signal_5209), .Q (signal_12721) ) ;
    buf_clk cell_7835 ( .C (clk), .D (signal_8474), .Q (signal_12723) ) ;
    buf_clk cell_7837 ( .C (clk), .D (signal_5215), .Q (signal_12725) ) ;
    buf_clk cell_7839 ( .C (clk), .D (signal_8480), .Q (signal_12727) ) ;
    buf_clk cell_7841 ( .C (clk), .D (signal_5221), .Q (signal_12729) ) ;
    buf_clk cell_7843 ( .C (clk), .D (signal_8486), .Q (signal_12731) ) ;
    buf_clk cell_7845 ( .C (clk), .D (signal_5227), .Q (signal_12733) ) ;
    buf_clk cell_7847 ( .C (clk), .D (signal_8492), .Q (signal_12735) ) ;
    buf_clk cell_7849 ( .C (clk), .D (signal_5272), .Q (signal_12737) ) ;
    buf_clk cell_7851 ( .C (clk), .D (signal_8564), .Q (signal_12739) ) ;
    buf_clk cell_7853 ( .C (clk), .D (signal_5278), .Q (signal_12741) ) ;
    buf_clk cell_7855 ( .C (clk), .D (signal_8570), .Q (signal_12743) ) ;
    buf_clk cell_7857 ( .C (clk), .D (signal_5284), .Q (signal_12745) ) ;
    buf_clk cell_7859 ( .C (clk), .D (signal_8576), .Q (signal_12747) ) ;
    buf_clk cell_7861 ( .C (clk), .D (signal_5290), .Q (signal_12749) ) ;
    buf_clk cell_7863 ( .C (clk), .D (signal_8582), .Q (signal_12751) ) ;
    buf_clk cell_7865 ( .C (clk), .D (signal_5296), .Q (signal_12753) ) ;
    buf_clk cell_7867 ( .C (clk), .D (signal_8588), .Q (signal_12755) ) ;
    buf_clk cell_7869 ( .C (clk), .D (signal_5302), .Q (signal_12757) ) ;
    buf_clk cell_7871 ( .C (clk), .D (signal_8594), .Q (signal_12759) ) ;
    buf_clk cell_7873 ( .C (clk), .D (signal_5308), .Q (signal_12761) ) ;
    buf_clk cell_7875 ( .C (clk), .D (signal_8600), .Q (signal_12763) ) ;
    buf_clk cell_7877 ( .C (clk), .D (signal_5319), .Q (signal_12765) ) ;
    buf_clk cell_7879 ( .C (clk), .D (signal_8606), .Q (signal_12767) ) ;
    buf_clk cell_7881 ( .C (clk), .D (signal_5325), .Q (signal_12769) ) ;
    buf_clk cell_7883 ( .C (clk), .D (signal_8612), .Q (signal_12771) ) ;
    buf_clk cell_7885 ( .C (clk), .D (signal_5331), .Q (signal_12773) ) ;
    buf_clk cell_7887 ( .C (clk), .D (signal_8618), .Q (signal_12775) ) ;
    buf_clk cell_7889 ( .C (clk), .D (signal_5342), .Q (signal_12777) ) ;
    buf_clk cell_7891 ( .C (clk), .D (signal_8624), .Q (signal_12779) ) ;
    buf_clk cell_7893 ( .C (clk), .D (signal_5348), .Q (signal_12781) ) ;
    buf_clk cell_7895 ( .C (clk), .D (signal_8630), .Q (signal_12783) ) ;
    buf_clk cell_7897 ( .C (clk), .D (signal_5354), .Q (signal_12785) ) ;
    buf_clk cell_7899 ( .C (clk), .D (signal_8636), .Q (signal_12787) ) ;
    buf_clk cell_8541 ( .C (clk), .D (signal_402), .Q (signal_13429) ) ;
    buf_clk cell_8549 ( .C (clk), .D (signal_396), .Q (signal_13437) ) ;
    buf_clk cell_8557 ( .C (clk), .D (signal_397), .Q (signal_13445) ) ;
    buf_clk cell_8565 ( .C (clk), .D (signal_398), .Q (signal_13453) ) ;
    buf_clk cell_8573 ( .C (clk), .D (signal_399), .Q (signal_13461) ) ;
    buf_clk cell_8581 ( .C (clk), .D (signal_400), .Q (signal_13469) ) ;
    buf_clk cell_8589 ( .C (clk), .D (signal_401), .Q (signal_13477) ) ;
    buf_clk cell_8597 ( .C (clk), .D (reset), .Q (signal_13485) ) ;
    buf_clk cell_8605 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_13493) ) ;
    buf_clk cell_8613 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_13501) ) ;
    buf_clk cell_8621 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_13509) ) ;
    buf_clk cell_8629 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_13517) ) ;
    buf_clk cell_8637 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_13525) ) ;
    buf_clk cell_8645 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_13533) ) ;
    buf_clk cell_8653 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_13541) ) ;
    buf_clk cell_8661 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_13549) ) ;
    buf_clk cell_8669 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_13557) ) ;
    buf_clk cell_8677 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_13565) ) ;
    buf_clk cell_8685 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_13573) ) ;
    buf_clk cell_8693 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_13581) ) ;
    buf_clk cell_8701 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_13589) ) ;
    buf_clk cell_8709 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_13597) ) ;
    buf_clk cell_8717 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_13605) ) ;
    buf_clk cell_8725 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_13613) ) ;
    buf_clk cell_8733 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_13621) ) ;
    buf_clk cell_8741 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_13629) ) ;
    buf_clk cell_8749 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_13637) ) ;
    buf_clk cell_8757 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_13645) ) ;
    buf_clk cell_8765 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_13653) ) ;
    buf_clk cell_8773 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_13661) ) ;
    buf_clk cell_8781 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_13669) ) ;
    buf_clk cell_8789 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_13677) ) ;
    buf_clk cell_8797 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_13685) ) ;
    buf_clk cell_8805 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_13693) ) ;
    buf_clk cell_8813 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_13701) ) ;
    buf_clk cell_8821 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_13709) ) ;
    buf_clk cell_8829 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_13717) ) ;
    buf_clk cell_8837 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_13725) ) ;
    buf_clk cell_8845 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_13733) ) ;
    buf_clk cell_8853 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_13741) ) ;
    buf_clk cell_8861 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_13749) ) ;
    buf_clk cell_8869 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_13757) ) ;
    buf_clk cell_8877 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_13765) ) ;
    buf_clk cell_8885 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_13773) ) ;
    buf_clk cell_8893 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_13781) ) ;
    buf_clk cell_8901 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_13789) ) ;
    buf_clk cell_8909 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_13797) ) ;
    buf_clk cell_8917 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_13805) ) ;
    buf_clk cell_8925 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_13813) ) ;
    buf_clk cell_8933 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_13821) ) ;
    buf_clk cell_8941 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_13829) ) ;
    buf_clk cell_8949 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_13837) ) ;
    buf_clk cell_8957 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_13845) ) ;
    buf_clk cell_8965 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_13853) ) ;
    buf_clk cell_8973 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_13861) ) ;
    buf_clk cell_8981 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_13869) ) ;
    buf_clk cell_8989 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_13877) ) ;
    buf_clk cell_8997 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_13885) ) ;
    buf_clk cell_9005 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_13893) ) ;
    buf_clk cell_9013 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_13901) ) ;
    buf_clk cell_9021 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_13909) ) ;
    buf_clk cell_9029 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_13917) ) ;
    buf_clk cell_9037 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_13925) ) ;
    buf_clk cell_9045 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_13933) ) ;
    buf_clk cell_9053 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_13941) ) ;
    buf_clk cell_9061 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_13949) ) ;
    buf_clk cell_9069 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_13957) ) ;
    buf_clk cell_9077 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_13965) ) ;
    buf_clk cell_9085 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_13973) ) ;
    buf_clk cell_9093 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_13981) ) ;
    buf_clk cell_9101 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_13989) ) ;
    buf_clk cell_9109 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_13997) ) ;
    buf_clk cell_9117 ( .C (clk), .D (plaintext_s0[32]), .Q (signal_14005) ) ;
    buf_clk cell_9125 ( .C (clk), .D (plaintext_s1[32]), .Q (signal_14013) ) ;
    buf_clk cell_9133 ( .C (clk), .D (plaintext_s0[33]), .Q (signal_14021) ) ;
    buf_clk cell_9141 ( .C (clk), .D (plaintext_s1[33]), .Q (signal_14029) ) ;
    buf_clk cell_9149 ( .C (clk), .D (plaintext_s0[34]), .Q (signal_14037) ) ;
    buf_clk cell_9157 ( .C (clk), .D (plaintext_s1[34]), .Q (signal_14045) ) ;
    buf_clk cell_9165 ( .C (clk), .D (plaintext_s0[35]), .Q (signal_14053) ) ;
    buf_clk cell_9173 ( .C (clk), .D (plaintext_s1[35]), .Q (signal_14061) ) ;
    buf_clk cell_9181 ( .C (clk), .D (plaintext_s0[36]), .Q (signal_14069) ) ;
    buf_clk cell_9189 ( .C (clk), .D (plaintext_s1[36]), .Q (signal_14077) ) ;
    buf_clk cell_9197 ( .C (clk), .D (plaintext_s0[37]), .Q (signal_14085) ) ;
    buf_clk cell_9205 ( .C (clk), .D (plaintext_s1[37]), .Q (signal_14093) ) ;
    buf_clk cell_9213 ( .C (clk), .D (plaintext_s0[38]), .Q (signal_14101) ) ;
    buf_clk cell_9221 ( .C (clk), .D (plaintext_s1[38]), .Q (signal_14109) ) ;
    buf_clk cell_9229 ( .C (clk), .D (plaintext_s0[39]), .Q (signal_14117) ) ;
    buf_clk cell_9237 ( .C (clk), .D (plaintext_s1[39]), .Q (signal_14125) ) ;
    buf_clk cell_9245 ( .C (clk), .D (plaintext_s0[40]), .Q (signal_14133) ) ;
    buf_clk cell_9253 ( .C (clk), .D (plaintext_s1[40]), .Q (signal_14141) ) ;
    buf_clk cell_9261 ( .C (clk), .D (plaintext_s0[41]), .Q (signal_14149) ) ;
    buf_clk cell_9269 ( .C (clk), .D (plaintext_s1[41]), .Q (signal_14157) ) ;
    buf_clk cell_9277 ( .C (clk), .D (plaintext_s0[42]), .Q (signal_14165) ) ;
    buf_clk cell_9285 ( .C (clk), .D (plaintext_s1[42]), .Q (signal_14173) ) ;
    buf_clk cell_9293 ( .C (clk), .D (plaintext_s0[43]), .Q (signal_14181) ) ;
    buf_clk cell_9301 ( .C (clk), .D (plaintext_s1[43]), .Q (signal_14189) ) ;
    buf_clk cell_9309 ( .C (clk), .D (plaintext_s0[44]), .Q (signal_14197) ) ;
    buf_clk cell_9317 ( .C (clk), .D (plaintext_s1[44]), .Q (signal_14205) ) ;
    buf_clk cell_9325 ( .C (clk), .D (plaintext_s0[45]), .Q (signal_14213) ) ;
    buf_clk cell_9333 ( .C (clk), .D (plaintext_s1[45]), .Q (signal_14221) ) ;
    buf_clk cell_9341 ( .C (clk), .D (plaintext_s0[46]), .Q (signal_14229) ) ;
    buf_clk cell_9349 ( .C (clk), .D (plaintext_s1[46]), .Q (signal_14237) ) ;
    buf_clk cell_9357 ( .C (clk), .D (plaintext_s0[47]), .Q (signal_14245) ) ;
    buf_clk cell_9365 ( .C (clk), .D (plaintext_s1[47]), .Q (signal_14253) ) ;
    buf_clk cell_9373 ( .C (clk), .D (plaintext_s0[48]), .Q (signal_14261) ) ;
    buf_clk cell_9381 ( .C (clk), .D (plaintext_s1[48]), .Q (signal_14269) ) ;
    buf_clk cell_9389 ( .C (clk), .D (plaintext_s0[49]), .Q (signal_14277) ) ;
    buf_clk cell_9397 ( .C (clk), .D (plaintext_s1[49]), .Q (signal_14285) ) ;
    buf_clk cell_9405 ( .C (clk), .D (plaintext_s0[50]), .Q (signal_14293) ) ;
    buf_clk cell_9413 ( .C (clk), .D (plaintext_s1[50]), .Q (signal_14301) ) ;
    buf_clk cell_9421 ( .C (clk), .D (plaintext_s0[51]), .Q (signal_14309) ) ;
    buf_clk cell_9429 ( .C (clk), .D (plaintext_s1[51]), .Q (signal_14317) ) ;
    buf_clk cell_9437 ( .C (clk), .D (plaintext_s0[52]), .Q (signal_14325) ) ;
    buf_clk cell_9445 ( .C (clk), .D (plaintext_s1[52]), .Q (signal_14333) ) ;
    buf_clk cell_9453 ( .C (clk), .D (plaintext_s0[53]), .Q (signal_14341) ) ;
    buf_clk cell_9461 ( .C (clk), .D (plaintext_s1[53]), .Q (signal_14349) ) ;
    buf_clk cell_9469 ( .C (clk), .D (plaintext_s0[54]), .Q (signal_14357) ) ;
    buf_clk cell_9477 ( .C (clk), .D (plaintext_s1[54]), .Q (signal_14365) ) ;
    buf_clk cell_9485 ( .C (clk), .D (plaintext_s0[55]), .Q (signal_14373) ) ;
    buf_clk cell_9493 ( .C (clk), .D (plaintext_s1[55]), .Q (signal_14381) ) ;
    buf_clk cell_9501 ( .C (clk), .D (plaintext_s0[56]), .Q (signal_14389) ) ;
    buf_clk cell_9509 ( .C (clk), .D (plaintext_s1[56]), .Q (signal_14397) ) ;
    buf_clk cell_9517 ( .C (clk), .D (plaintext_s0[57]), .Q (signal_14405) ) ;
    buf_clk cell_9525 ( .C (clk), .D (plaintext_s1[57]), .Q (signal_14413) ) ;
    buf_clk cell_9533 ( .C (clk), .D (plaintext_s0[58]), .Q (signal_14421) ) ;
    buf_clk cell_9541 ( .C (clk), .D (plaintext_s1[58]), .Q (signal_14429) ) ;
    buf_clk cell_9549 ( .C (clk), .D (plaintext_s0[59]), .Q (signal_14437) ) ;
    buf_clk cell_9557 ( .C (clk), .D (plaintext_s1[59]), .Q (signal_14445) ) ;
    buf_clk cell_9565 ( .C (clk), .D (plaintext_s0[60]), .Q (signal_14453) ) ;
    buf_clk cell_9573 ( .C (clk), .D (plaintext_s1[60]), .Q (signal_14461) ) ;
    buf_clk cell_9581 ( .C (clk), .D (plaintext_s0[61]), .Q (signal_14469) ) ;
    buf_clk cell_9589 ( .C (clk), .D (plaintext_s1[61]), .Q (signal_14477) ) ;
    buf_clk cell_9597 ( .C (clk), .D (plaintext_s0[62]), .Q (signal_14485) ) ;
    buf_clk cell_9605 ( .C (clk), .D (plaintext_s1[62]), .Q (signal_14493) ) ;
    buf_clk cell_9613 ( .C (clk), .D (plaintext_s0[63]), .Q (signal_14501) ) ;
    buf_clk cell_9621 ( .C (clk), .D (plaintext_s1[63]), .Q (signal_14509) ) ;
    buf_clk cell_9629 ( .C (clk), .D (plaintext_s0[64]), .Q (signal_14517) ) ;
    buf_clk cell_9637 ( .C (clk), .D (plaintext_s1[64]), .Q (signal_14525) ) ;
    buf_clk cell_9645 ( .C (clk), .D (plaintext_s0[65]), .Q (signal_14533) ) ;
    buf_clk cell_9653 ( .C (clk), .D (plaintext_s1[65]), .Q (signal_14541) ) ;
    buf_clk cell_9661 ( .C (clk), .D (plaintext_s0[66]), .Q (signal_14549) ) ;
    buf_clk cell_9669 ( .C (clk), .D (plaintext_s1[66]), .Q (signal_14557) ) ;
    buf_clk cell_9677 ( .C (clk), .D (plaintext_s0[67]), .Q (signal_14565) ) ;
    buf_clk cell_9685 ( .C (clk), .D (plaintext_s1[67]), .Q (signal_14573) ) ;
    buf_clk cell_9693 ( .C (clk), .D (plaintext_s0[68]), .Q (signal_14581) ) ;
    buf_clk cell_9701 ( .C (clk), .D (plaintext_s1[68]), .Q (signal_14589) ) ;
    buf_clk cell_9709 ( .C (clk), .D (plaintext_s0[69]), .Q (signal_14597) ) ;
    buf_clk cell_9717 ( .C (clk), .D (plaintext_s1[69]), .Q (signal_14605) ) ;
    buf_clk cell_9725 ( .C (clk), .D (plaintext_s0[70]), .Q (signal_14613) ) ;
    buf_clk cell_9733 ( .C (clk), .D (plaintext_s1[70]), .Q (signal_14621) ) ;
    buf_clk cell_9741 ( .C (clk), .D (plaintext_s0[71]), .Q (signal_14629) ) ;
    buf_clk cell_9749 ( .C (clk), .D (plaintext_s1[71]), .Q (signal_14637) ) ;
    buf_clk cell_9757 ( .C (clk), .D (plaintext_s0[72]), .Q (signal_14645) ) ;
    buf_clk cell_9765 ( .C (clk), .D (plaintext_s1[72]), .Q (signal_14653) ) ;
    buf_clk cell_9773 ( .C (clk), .D (plaintext_s0[73]), .Q (signal_14661) ) ;
    buf_clk cell_9781 ( .C (clk), .D (plaintext_s1[73]), .Q (signal_14669) ) ;
    buf_clk cell_9789 ( .C (clk), .D (plaintext_s0[74]), .Q (signal_14677) ) ;
    buf_clk cell_9797 ( .C (clk), .D (plaintext_s1[74]), .Q (signal_14685) ) ;
    buf_clk cell_9805 ( .C (clk), .D (plaintext_s0[75]), .Q (signal_14693) ) ;
    buf_clk cell_9813 ( .C (clk), .D (plaintext_s1[75]), .Q (signal_14701) ) ;
    buf_clk cell_9821 ( .C (clk), .D (plaintext_s0[76]), .Q (signal_14709) ) ;
    buf_clk cell_9829 ( .C (clk), .D (plaintext_s1[76]), .Q (signal_14717) ) ;
    buf_clk cell_9837 ( .C (clk), .D (plaintext_s0[77]), .Q (signal_14725) ) ;
    buf_clk cell_9845 ( .C (clk), .D (plaintext_s1[77]), .Q (signal_14733) ) ;
    buf_clk cell_9853 ( .C (clk), .D (plaintext_s0[78]), .Q (signal_14741) ) ;
    buf_clk cell_9861 ( .C (clk), .D (plaintext_s1[78]), .Q (signal_14749) ) ;
    buf_clk cell_9869 ( .C (clk), .D (plaintext_s0[79]), .Q (signal_14757) ) ;
    buf_clk cell_9877 ( .C (clk), .D (plaintext_s1[79]), .Q (signal_14765) ) ;
    buf_clk cell_9885 ( .C (clk), .D (plaintext_s0[80]), .Q (signal_14773) ) ;
    buf_clk cell_9893 ( .C (clk), .D (plaintext_s1[80]), .Q (signal_14781) ) ;
    buf_clk cell_9901 ( .C (clk), .D (plaintext_s0[81]), .Q (signal_14789) ) ;
    buf_clk cell_9909 ( .C (clk), .D (plaintext_s1[81]), .Q (signal_14797) ) ;
    buf_clk cell_9917 ( .C (clk), .D (plaintext_s0[82]), .Q (signal_14805) ) ;
    buf_clk cell_9925 ( .C (clk), .D (plaintext_s1[82]), .Q (signal_14813) ) ;
    buf_clk cell_9933 ( .C (clk), .D (plaintext_s0[83]), .Q (signal_14821) ) ;
    buf_clk cell_9941 ( .C (clk), .D (plaintext_s1[83]), .Q (signal_14829) ) ;
    buf_clk cell_9949 ( .C (clk), .D (plaintext_s0[84]), .Q (signal_14837) ) ;
    buf_clk cell_9957 ( .C (clk), .D (plaintext_s1[84]), .Q (signal_14845) ) ;
    buf_clk cell_9965 ( .C (clk), .D (plaintext_s0[85]), .Q (signal_14853) ) ;
    buf_clk cell_9973 ( .C (clk), .D (plaintext_s1[85]), .Q (signal_14861) ) ;
    buf_clk cell_9981 ( .C (clk), .D (plaintext_s0[86]), .Q (signal_14869) ) ;
    buf_clk cell_9989 ( .C (clk), .D (plaintext_s1[86]), .Q (signal_14877) ) ;
    buf_clk cell_9997 ( .C (clk), .D (plaintext_s0[87]), .Q (signal_14885) ) ;
    buf_clk cell_10005 ( .C (clk), .D (plaintext_s1[87]), .Q (signal_14893) ) ;
    buf_clk cell_10013 ( .C (clk), .D (plaintext_s0[88]), .Q (signal_14901) ) ;
    buf_clk cell_10021 ( .C (clk), .D (plaintext_s1[88]), .Q (signal_14909) ) ;
    buf_clk cell_10029 ( .C (clk), .D (plaintext_s0[89]), .Q (signal_14917) ) ;
    buf_clk cell_10037 ( .C (clk), .D (plaintext_s1[89]), .Q (signal_14925) ) ;
    buf_clk cell_10045 ( .C (clk), .D (plaintext_s0[90]), .Q (signal_14933) ) ;
    buf_clk cell_10053 ( .C (clk), .D (plaintext_s1[90]), .Q (signal_14941) ) ;
    buf_clk cell_10061 ( .C (clk), .D (plaintext_s0[91]), .Q (signal_14949) ) ;
    buf_clk cell_10069 ( .C (clk), .D (plaintext_s1[91]), .Q (signal_14957) ) ;
    buf_clk cell_10077 ( .C (clk), .D (plaintext_s0[92]), .Q (signal_14965) ) ;
    buf_clk cell_10085 ( .C (clk), .D (plaintext_s1[92]), .Q (signal_14973) ) ;
    buf_clk cell_10093 ( .C (clk), .D (plaintext_s0[93]), .Q (signal_14981) ) ;
    buf_clk cell_10101 ( .C (clk), .D (plaintext_s1[93]), .Q (signal_14989) ) ;
    buf_clk cell_10109 ( .C (clk), .D (plaintext_s0[94]), .Q (signal_14997) ) ;
    buf_clk cell_10117 ( .C (clk), .D (plaintext_s1[94]), .Q (signal_15005) ) ;
    buf_clk cell_10125 ( .C (clk), .D (plaintext_s0[95]), .Q (signal_15013) ) ;
    buf_clk cell_10133 ( .C (clk), .D (plaintext_s1[95]), .Q (signal_15021) ) ;
    buf_clk cell_10141 ( .C (clk), .D (plaintext_s0[96]), .Q (signal_15029) ) ;
    buf_clk cell_10149 ( .C (clk), .D (plaintext_s1[96]), .Q (signal_15037) ) ;
    buf_clk cell_10157 ( .C (clk), .D (plaintext_s0[97]), .Q (signal_15045) ) ;
    buf_clk cell_10165 ( .C (clk), .D (plaintext_s1[97]), .Q (signal_15053) ) ;
    buf_clk cell_10173 ( .C (clk), .D (plaintext_s0[98]), .Q (signal_15061) ) ;
    buf_clk cell_10181 ( .C (clk), .D (plaintext_s1[98]), .Q (signal_15069) ) ;
    buf_clk cell_10189 ( .C (clk), .D (plaintext_s0[99]), .Q (signal_15077) ) ;
    buf_clk cell_10197 ( .C (clk), .D (plaintext_s1[99]), .Q (signal_15085) ) ;
    buf_clk cell_10205 ( .C (clk), .D (plaintext_s0[100]), .Q (signal_15093) ) ;
    buf_clk cell_10213 ( .C (clk), .D (plaintext_s1[100]), .Q (signal_15101) ) ;
    buf_clk cell_10221 ( .C (clk), .D (plaintext_s0[101]), .Q (signal_15109) ) ;
    buf_clk cell_10229 ( .C (clk), .D (plaintext_s1[101]), .Q (signal_15117) ) ;
    buf_clk cell_10237 ( .C (clk), .D (plaintext_s0[102]), .Q (signal_15125) ) ;
    buf_clk cell_10245 ( .C (clk), .D (plaintext_s1[102]), .Q (signal_15133) ) ;
    buf_clk cell_10253 ( .C (clk), .D (plaintext_s0[103]), .Q (signal_15141) ) ;
    buf_clk cell_10261 ( .C (clk), .D (plaintext_s1[103]), .Q (signal_15149) ) ;
    buf_clk cell_10269 ( .C (clk), .D (plaintext_s0[104]), .Q (signal_15157) ) ;
    buf_clk cell_10277 ( .C (clk), .D (plaintext_s1[104]), .Q (signal_15165) ) ;
    buf_clk cell_10285 ( .C (clk), .D (plaintext_s0[105]), .Q (signal_15173) ) ;
    buf_clk cell_10293 ( .C (clk), .D (plaintext_s1[105]), .Q (signal_15181) ) ;
    buf_clk cell_10301 ( .C (clk), .D (plaintext_s0[106]), .Q (signal_15189) ) ;
    buf_clk cell_10309 ( .C (clk), .D (plaintext_s1[106]), .Q (signal_15197) ) ;
    buf_clk cell_10317 ( .C (clk), .D (plaintext_s0[107]), .Q (signal_15205) ) ;
    buf_clk cell_10325 ( .C (clk), .D (plaintext_s1[107]), .Q (signal_15213) ) ;
    buf_clk cell_10333 ( .C (clk), .D (plaintext_s0[108]), .Q (signal_15221) ) ;
    buf_clk cell_10341 ( .C (clk), .D (plaintext_s1[108]), .Q (signal_15229) ) ;
    buf_clk cell_10349 ( .C (clk), .D (plaintext_s0[109]), .Q (signal_15237) ) ;
    buf_clk cell_10357 ( .C (clk), .D (plaintext_s1[109]), .Q (signal_15245) ) ;
    buf_clk cell_10365 ( .C (clk), .D (plaintext_s0[110]), .Q (signal_15253) ) ;
    buf_clk cell_10373 ( .C (clk), .D (plaintext_s1[110]), .Q (signal_15261) ) ;
    buf_clk cell_10381 ( .C (clk), .D (plaintext_s0[111]), .Q (signal_15269) ) ;
    buf_clk cell_10389 ( .C (clk), .D (plaintext_s1[111]), .Q (signal_15277) ) ;
    buf_clk cell_10397 ( .C (clk), .D (plaintext_s0[112]), .Q (signal_15285) ) ;
    buf_clk cell_10405 ( .C (clk), .D (plaintext_s1[112]), .Q (signal_15293) ) ;
    buf_clk cell_10413 ( .C (clk), .D (plaintext_s0[113]), .Q (signal_15301) ) ;
    buf_clk cell_10421 ( .C (clk), .D (plaintext_s1[113]), .Q (signal_15309) ) ;
    buf_clk cell_10429 ( .C (clk), .D (plaintext_s0[114]), .Q (signal_15317) ) ;
    buf_clk cell_10437 ( .C (clk), .D (plaintext_s1[114]), .Q (signal_15325) ) ;
    buf_clk cell_10445 ( .C (clk), .D (plaintext_s0[115]), .Q (signal_15333) ) ;
    buf_clk cell_10453 ( .C (clk), .D (plaintext_s1[115]), .Q (signal_15341) ) ;
    buf_clk cell_10461 ( .C (clk), .D (plaintext_s0[116]), .Q (signal_15349) ) ;
    buf_clk cell_10469 ( .C (clk), .D (plaintext_s1[116]), .Q (signal_15357) ) ;
    buf_clk cell_10477 ( .C (clk), .D (plaintext_s0[117]), .Q (signal_15365) ) ;
    buf_clk cell_10485 ( .C (clk), .D (plaintext_s1[117]), .Q (signal_15373) ) ;
    buf_clk cell_10493 ( .C (clk), .D (plaintext_s0[118]), .Q (signal_15381) ) ;
    buf_clk cell_10501 ( .C (clk), .D (plaintext_s1[118]), .Q (signal_15389) ) ;
    buf_clk cell_10509 ( .C (clk), .D (plaintext_s0[119]), .Q (signal_15397) ) ;
    buf_clk cell_10517 ( .C (clk), .D (plaintext_s1[119]), .Q (signal_15405) ) ;
    buf_clk cell_10525 ( .C (clk), .D (plaintext_s0[120]), .Q (signal_15413) ) ;
    buf_clk cell_10533 ( .C (clk), .D (plaintext_s1[120]), .Q (signal_15421) ) ;
    buf_clk cell_10541 ( .C (clk), .D (plaintext_s0[121]), .Q (signal_15429) ) ;
    buf_clk cell_10549 ( .C (clk), .D (plaintext_s1[121]), .Q (signal_15437) ) ;
    buf_clk cell_10557 ( .C (clk), .D (plaintext_s0[122]), .Q (signal_15445) ) ;
    buf_clk cell_10565 ( .C (clk), .D (plaintext_s1[122]), .Q (signal_15453) ) ;
    buf_clk cell_10573 ( .C (clk), .D (plaintext_s0[123]), .Q (signal_15461) ) ;
    buf_clk cell_10581 ( .C (clk), .D (plaintext_s1[123]), .Q (signal_15469) ) ;
    buf_clk cell_10589 ( .C (clk), .D (plaintext_s0[124]), .Q (signal_15477) ) ;
    buf_clk cell_10597 ( .C (clk), .D (plaintext_s1[124]), .Q (signal_15485) ) ;
    buf_clk cell_10605 ( .C (clk), .D (plaintext_s0[125]), .Q (signal_15493) ) ;
    buf_clk cell_10613 ( .C (clk), .D (plaintext_s1[125]), .Q (signal_15501) ) ;
    buf_clk cell_10621 ( .C (clk), .D (plaintext_s0[126]), .Q (signal_15509) ) ;
    buf_clk cell_10629 ( .C (clk), .D (plaintext_s1[126]), .Q (signal_15517) ) ;
    buf_clk cell_10637 ( .C (clk), .D (plaintext_s0[127]), .Q (signal_15525) ) ;
    buf_clk cell_10645 ( .C (clk), .D (plaintext_s1[127]), .Q (signal_15533) ) ;
    buf_clk cell_10653 ( .C (clk), .D (key_s0[0]), .Q (signal_15541) ) ;
    buf_clk cell_10661 ( .C (clk), .D (key_s1[0]), .Q (signal_15549) ) ;
    buf_clk cell_10669 ( .C (clk), .D (key_s0[1]), .Q (signal_15557) ) ;
    buf_clk cell_10677 ( .C (clk), .D (key_s1[1]), .Q (signal_15565) ) ;
    buf_clk cell_10685 ( .C (clk), .D (key_s0[2]), .Q (signal_15573) ) ;
    buf_clk cell_10693 ( .C (clk), .D (key_s1[2]), .Q (signal_15581) ) ;
    buf_clk cell_10701 ( .C (clk), .D (key_s0[3]), .Q (signal_15589) ) ;
    buf_clk cell_10709 ( .C (clk), .D (key_s1[3]), .Q (signal_15597) ) ;
    buf_clk cell_10717 ( .C (clk), .D (key_s0[4]), .Q (signal_15605) ) ;
    buf_clk cell_10725 ( .C (clk), .D (key_s1[4]), .Q (signal_15613) ) ;
    buf_clk cell_10733 ( .C (clk), .D (key_s0[5]), .Q (signal_15621) ) ;
    buf_clk cell_10741 ( .C (clk), .D (key_s1[5]), .Q (signal_15629) ) ;
    buf_clk cell_10749 ( .C (clk), .D (key_s0[6]), .Q (signal_15637) ) ;
    buf_clk cell_10757 ( .C (clk), .D (key_s1[6]), .Q (signal_15645) ) ;
    buf_clk cell_10765 ( .C (clk), .D (key_s0[7]), .Q (signal_15653) ) ;
    buf_clk cell_10773 ( .C (clk), .D (key_s1[7]), .Q (signal_15661) ) ;
    buf_clk cell_10781 ( .C (clk), .D (key_s0[8]), .Q (signal_15669) ) ;
    buf_clk cell_10789 ( .C (clk), .D (key_s1[8]), .Q (signal_15677) ) ;
    buf_clk cell_10797 ( .C (clk), .D (key_s0[9]), .Q (signal_15685) ) ;
    buf_clk cell_10805 ( .C (clk), .D (key_s1[9]), .Q (signal_15693) ) ;
    buf_clk cell_10813 ( .C (clk), .D (key_s0[10]), .Q (signal_15701) ) ;
    buf_clk cell_10821 ( .C (clk), .D (key_s1[10]), .Q (signal_15709) ) ;
    buf_clk cell_10829 ( .C (clk), .D (key_s0[11]), .Q (signal_15717) ) ;
    buf_clk cell_10837 ( .C (clk), .D (key_s1[11]), .Q (signal_15725) ) ;
    buf_clk cell_10845 ( .C (clk), .D (key_s0[12]), .Q (signal_15733) ) ;
    buf_clk cell_10853 ( .C (clk), .D (key_s1[12]), .Q (signal_15741) ) ;
    buf_clk cell_10861 ( .C (clk), .D (key_s0[13]), .Q (signal_15749) ) ;
    buf_clk cell_10869 ( .C (clk), .D (key_s1[13]), .Q (signal_15757) ) ;
    buf_clk cell_10877 ( .C (clk), .D (key_s0[14]), .Q (signal_15765) ) ;
    buf_clk cell_10885 ( .C (clk), .D (key_s1[14]), .Q (signal_15773) ) ;
    buf_clk cell_10893 ( .C (clk), .D (key_s0[15]), .Q (signal_15781) ) ;
    buf_clk cell_10901 ( .C (clk), .D (key_s1[15]), .Q (signal_15789) ) ;
    buf_clk cell_10909 ( .C (clk), .D (key_s0[16]), .Q (signal_15797) ) ;
    buf_clk cell_10917 ( .C (clk), .D (key_s1[16]), .Q (signal_15805) ) ;
    buf_clk cell_10925 ( .C (clk), .D (key_s0[17]), .Q (signal_15813) ) ;
    buf_clk cell_10933 ( .C (clk), .D (key_s1[17]), .Q (signal_15821) ) ;
    buf_clk cell_10941 ( .C (clk), .D (key_s0[18]), .Q (signal_15829) ) ;
    buf_clk cell_10949 ( .C (clk), .D (key_s1[18]), .Q (signal_15837) ) ;
    buf_clk cell_10957 ( .C (clk), .D (key_s0[19]), .Q (signal_15845) ) ;
    buf_clk cell_10965 ( .C (clk), .D (key_s1[19]), .Q (signal_15853) ) ;
    buf_clk cell_10973 ( .C (clk), .D (key_s0[20]), .Q (signal_15861) ) ;
    buf_clk cell_10981 ( .C (clk), .D (key_s1[20]), .Q (signal_15869) ) ;
    buf_clk cell_10989 ( .C (clk), .D (key_s0[21]), .Q (signal_15877) ) ;
    buf_clk cell_10997 ( .C (clk), .D (key_s1[21]), .Q (signal_15885) ) ;
    buf_clk cell_11005 ( .C (clk), .D (key_s0[22]), .Q (signal_15893) ) ;
    buf_clk cell_11013 ( .C (clk), .D (key_s1[22]), .Q (signal_15901) ) ;
    buf_clk cell_11021 ( .C (clk), .D (key_s0[23]), .Q (signal_15909) ) ;
    buf_clk cell_11029 ( .C (clk), .D (key_s1[23]), .Q (signal_15917) ) ;
    buf_clk cell_11037 ( .C (clk), .D (key_s0[24]), .Q (signal_15925) ) ;
    buf_clk cell_11045 ( .C (clk), .D (key_s1[24]), .Q (signal_15933) ) ;
    buf_clk cell_11053 ( .C (clk), .D (key_s0[25]), .Q (signal_15941) ) ;
    buf_clk cell_11061 ( .C (clk), .D (key_s1[25]), .Q (signal_15949) ) ;
    buf_clk cell_11069 ( .C (clk), .D (key_s0[26]), .Q (signal_15957) ) ;
    buf_clk cell_11077 ( .C (clk), .D (key_s1[26]), .Q (signal_15965) ) ;
    buf_clk cell_11085 ( .C (clk), .D (key_s0[27]), .Q (signal_15973) ) ;
    buf_clk cell_11093 ( .C (clk), .D (key_s1[27]), .Q (signal_15981) ) ;
    buf_clk cell_11101 ( .C (clk), .D (key_s0[28]), .Q (signal_15989) ) ;
    buf_clk cell_11109 ( .C (clk), .D (key_s1[28]), .Q (signal_15997) ) ;
    buf_clk cell_11117 ( .C (clk), .D (key_s0[29]), .Q (signal_16005) ) ;
    buf_clk cell_11125 ( .C (clk), .D (key_s1[29]), .Q (signal_16013) ) ;
    buf_clk cell_11133 ( .C (clk), .D (key_s0[30]), .Q (signal_16021) ) ;
    buf_clk cell_11141 ( .C (clk), .D (key_s1[30]), .Q (signal_16029) ) ;
    buf_clk cell_11149 ( .C (clk), .D (key_s0[31]), .Q (signal_16037) ) ;
    buf_clk cell_11157 ( .C (clk), .D (key_s1[31]), .Q (signal_16045) ) ;
    buf_clk cell_11165 ( .C (clk), .D (key_s0[32]), .Q (signal_16053) ) ;
    buf_clk cell_11173 ( .C (clk), .D (key_s1[32]), .Q (signal_16061) ) ;
    buf_clk cell_11181 ( .C (clk), .D (key_s0[33]), .Q (signal_16069) ) ;
    buf_clk cell_11189 ( .C (clk), .D (key_s1[33]), .Q (signal_16077) ) ;
    buf_clk cell_11197 ( .C (clk), .D (key_s0[34]), .Q (signal_16085) ) ;
    buf_clk cell_11205 ( .C (clk), .D (key_s1[34]), .Q (signal_16093) ) ;
    buf_clk cell_11213 ( .C (clk), .D (key_s0[35]), .Q (signal_16101) ) ;
    buf_clk cell_11221 ( .C (clk), .D (key_s1[35]), .Q (signal_16109) ) ;
    buf_clk cell_11229 ( .C (clk), .D (key_s0[36]), .Q (signal_16117) ) ;
    buf_clk cell_11237 ( .C (clk), .D (key_s1[36]), .Q (signal_16125) ) ;
    buf_clk cell_11245 ( .C (clk), .D (key_s0[37]), .Q (signal_16133) ) ;
    buf_clk cell_11253 ( .C (clk), .D (key_s1[37]), .Q (signal_16141) ) ;
    buf_clk cell_11261 ( .C (clk), .D (key_s0[38]), .Q (signal_16149) ) ;
    buf_clk cell_11269 ( .C (clk), .D (key_s1[38]), .Q (signal_16157) ) ;
    buf_clk cell_11277 ( .C (clk), .D (key_s0[39]), .Q (signal_16165) ) ;
    buf_clk cell_11285 ( .C (clk), .D (key_s1[39]), .Q (signal_16173) ) ;
    buf_clk cell_11293 ( .C (clk), .D (key_s0[40]), .Q (signal_16181) ) ;
    buf_clk cell_11301 ( .C (clk), .D (key_s1[40]), .Q (signal_16189) ) ;
    buf_clk cell_11309 ( .C (clk), .D (key_s0[41]), .Q (signal_16197) ) ;
    buf_clk cell_11317 ( .C (clk), .D (key_s1[41]), .Q (signal_16205) ) ;
    buf_clk cell_11325 ( .C (clk), .D (key_s0[42]), .Q (signal_16213) ) ;
    buf_clk cell_11333 ( .C (clk), .D (key_s1[42]), .Q (signal_16221) ) ;
    buf_clk cell_11341 ( .C (clk), .D (key_s0[43]), .Q (signal_16229) ) ;
    buf_clk cell_11349 ( .C (clk), .D (key_s1[43]), .Q (signal_16237) ) ;
    buf_clk cell_11357 ( .C (clk), .D (key_s0[44]), .Q (signal_16245) ) ;
    buf_clk cell_11365 ( .C (clk), .D (key_s1[44]), .Q (signal_16253) ) ;
    buf_clk cell_11373 ( .C (clk), .D (key_s0[45]), .Q (signal_16261) ) ;
    buf_clk cell_11381 ( .C (clk), .D (key_s1[45]), .Q (signal_16269) ) ;
    buf_clk cell_11389 ( .C (clk), .D (key_s0[46]), .Q (signal_16277) ) ;
    buf_clk cell_11397 ( .C (clk), .D (key_s1[46]), .Q (signal_16285) ) ;
    buf_clk cell_11405 ( .C (clk), .D (key_s0[47]), .Q (signal_16293) ) ;
    buf_clk cell_11413 ( .C (clk), .D (key_s1[47]), .Q (signal_16301) ) ;
    buf_clk cell_11421 ( .C (clk), .D (key_s0[48]), .Q (signal_16309) ) ;
    buf_clk cell_11429 ( .C (clk), .D (key_s1[48]), .Q (signal_16317) ) ;
    buf_clk cell_11437 ( .C (clk), .D (key_s0[49]), .Q (signal_16325) ) ;
    buf_clk cell_11445 ( .C (clk), .D (key_s1[49]), .Q (signal_16333) ) ;
    buf_clk cell_11453 ( .C (clk), .D (key_s0[50]), .Q (signal_16341) ) ;
    buf_clk cell_11461 ( .C (clk), .D (key_s1[50]), .Q (signal_16349) ) ;
    buf_clk cell_11469 ( .C (clk), .D (key_s0[51]), .Q (signal_16357) ) ;
    buf_clk cell_11477 ( .C (clk), .D (key_s1[51]), .Q (signal_16365) ) ;
    buf_clk cell_11485 ( .C (clk), .D (key_s0[52]), .Q (signal_16373) ) ;
    buf_clk cell_11493 ( .C (clk), .D (key_s1[52]), .Q (signal_16381) ) ;
    buf_clk cell_11501 ( .C (clk), .D (key_s0[53]), .Q (signal_16389) ) ;
    buf_clk cell_11509 ( .C (clk), .D (key_s1[53]), .Q (signal_16397) ) ;
    buf_clk cell_11517 ( .C (clk), .D (key_s0[54]), .Q (signal_16405) ) ;
    buf_clk cell_11525 ( .C (clk), .D (key_s1[54]), .Q (signal_16413) ) ;
    buf_clk cell_11533 ( .C (clk), .D (key_s0[55]), .Q (signal_16421) ) ;
    buf_clk cell_11541 ( .C (clk), .D (key_s1[55]), .Q (signal_16429) ) ;
    buf_clk cell_11549 ( .C (clk), .D (key_s0[56]), .Q (signal_16437) ) ;
    buf_clk cell_11557 ( .C (clk), .D (key_s1[56]), .Q (signal_16445) ) ;
    buf_clk cell_11565 ( .C (clk), .D (key_s0[57]), .Q (signal_16453) ) ;
    buf_clk cell_11573 ( .C (clk), .D (key_s1[57]), .Q (signal_16461) ) ;
    buf_clk cell_11581 ( .C (clk), .D (key_s0[58]), .Q (signal_16469) ) ;
    buf_clk cell_11589 ( .C (clk), .D (key_s1[58]), .Q (signal_16477) ) ;
    buf_clk cell_11597 ( .C (clk), .D (key_s0[59]), .Q (signal_16485) ) ;
    buf_clk cell_11605 ( .C (clk), .D (key_s1[59]), .Q (signal_16493) ) ;
    buf_clk cell_11613 ( .C (clk), .D (key_s0[60]), .Q (signal_16501) ) ;
    buf_clk cell_11621 ( .C (clk), .D (key_s1[60]), .Q (signal_16509) ) ;
    buf_clk cell_11629 ( .C (clk), .D (key_s0[61]), .Q (signal_16517) ) ;
    buf_clk cell_11637 ( .C (clk), .D (key_s1[61]), .Q (signal_16525) ) ;
    buf_clk cell_11645 ( .C (clk), .D (key_s0[62]), .Q (signal_16533) ) ;
    buf_clk cell_11653 ( .C (clk), .D (key_s1[62]), .Q (signal_16541) ) ;
    buf_clk cell_11661 ( .C (clk), .D (key_s0[63]), .Q (signal_16549) ) ;
    buf_clk cell_11669 ( .C (clk), .D (key_s1[63]), .Q (signal_16557) ) ;
    buf_clk cell_11677 ( .C (clk), .D (key_s0[64]), .Q (signal_16565) ) ;
    buf_clk cell_11685 ( .C (clk), .D (key_s1[64]), .Q (signal_16573) ) ;
    buf_clk cell_11693 ( .C (clk), .D (key_s0[65]), .Q (signal_16581) ) ;
    buf_clk cell_11701 ( .C (clk), .D (key_s1[65]), .Q (signal_16589) ) ;
    buf_clk cell_11709 ( .C (clk), .D (key_s0[66]), .Q (signal_16597) ) ;
    buf_clk cell_11717 ( .C (clk), .D (key_s1[66]), .Q (signal_16605) ) ;
    buf_clk cell_11725 ( .C (clk), .D (key_s0[67]), .Q (signal_16613) ) ;
    buf_clk cell_11733 ( .C (clk), .D (key_s1[67]), .Q (signal_16621) ) ;
    buf_clk cell_11741 ( .C (clk), .D (key_s0[68]), .Q (signal_16629) ) ;
    buf_clk cell_11749 ( .C (clk), .D (key_s1[68]), .Q (signal_16637) ) ;
    buf_clk cell_11757 ( .C (clk), .D (key_s0[69]), .Q (signal_16645) ) ;
    buf_clk cell_11765 ( .C (clk), .D (key_s1[69]), .Q (signal_16653) ) ;
    buf_clk cell_11773 ( .C (clk), .D (key_s0[70]), .Q (signal_16661) ) ;
    buf_clk cell_11781 ( .C (clk), .D (key_s1[70]), .Q (signal_16669) ) ;
    buf_clk cell_11789 ( .C (clk), .D (key_s0[71]), .Q (signal_16677) ) ;
    buf_clk cell_11797 ( .C (clk), .D (key_s1[71]), .Q (signal_16685) ) ;
    buf_clk cell_11805 ( .C (clk), .D (key_s0[72]), .Q (signal_16693) ) ;
    buf_clk cell_11813 ( .C (clk), .D (key_s1[72]), .Q (signal_16701) ) ;
    buf_clk cell_11821 ( .C (clk), .D (key_s0[73]), .Q (signal_16709) ) ;
    buf_clk cell_11829 ( .C (clk), .D (key_s1[73]), .Q (signal_16717) ) ;
    buf_clk cell_11837 ( .C (clk), .D (key_s0[74]), .Q (signal_16725) ) ;
    buf_clk cell_11845 ( .C (clk), .D (key_s1[74]), .Q (signal_16733) ) ;
    buf_clk cell_11853 ( .C (clk), .D (key_s0[75]), .Q (signal_16741) ) ;
    buf_clk cell_11861 ( .C (clk), .D (key_s1[75]), .Q (signal_16749) ) ;
    buf_clk cell_11869 ( .C (clk), .D (key_s0[76]), .Q (signal_16757) ) ;
    buf_clk cell_11877 ( .C (clk), .D (key_s1[76]), .Q (signal_16765) ) ;
    buf_clk cell_11885 ( .C (clk), .D (key_s0[77]), .Q (signal_16773) ) ;
    buf_clk cell_11893 ( .C (clk), .D (key_s1[77]), .Q (signal_16781) ) ;
    buf_clk cell_11901 ( .C (clk), .D (key_s0[78]), .Q (signal_16789) ) ;
    buf_clk cell_11909 ( .C (clk), .D (key_s1[78]), .Q (signal_16797) ) ;
    buf_clk cell_11917 ( .C (clk), .D (key_s0[79]), .Q (signal_16805) ) ;
    buf_clk cell_11925 ( .C (clk), .D (key_s1[79]), .Q (signal_16813) ) ;
    buf_clk cell_11933 ( .C (clk), .D (key_s0[80]), .Q (signal_16821) ) ;
    buf_clk cell_11941 ( .C (clk), .D (key_s1[80]), .Q (signal_16829) ) ;
    buf_clk cell_11949 ( .C (clk), .D (key_s0[81]), .Q (signal_16837) ) ;
    buf_clk cell_11957 ( .C (clk), .D (key_s1[81]), .Q (signal_16845) ) ;
    buf_clk cell_11965 ( .C (clk), .D (key_s0[82]), .Q (signal_16853) ) ;
    buf_clk cell_11973 ( .C (clk), .D (key_s1[82]), .Q (signal_16861) ) ;
    buf_clk cell_11981 ( .C (clk), .D (key_s0[83]), .Q (signal_16869) ) ;
    buf_clk cell_11989 ( .C (clk), .D (key_s1[83]), .Q (signal_16877) ) ;
    buf_clk cell_11997 ( .C (clk), .D (key_s0[84]), .Q (signal_16885) ) ;
    buf_clk cell_12005 ( .C (clk), .D (key_s1[84]), .Q (signal_16893) ) ;
    buf_clk cell_12013 ( .C (clk), .D (key_s0[85]), .Q (signal_16901) ) ;
    buf_clk cell_12021 ( .C (clk), .D (key_s1[85]), .Q (signal_16909) ) ;
    buf_clk cell_12029 ( .C (clk), .D (key_s0[86]), .Q (signal_16917) ) ;
    buf_clk cell_12037 ( .C (clk), .D (key_s1[86]), .Q (signal_16925) ) ;
    buf_clk cell_12045 ( .C (clk), .D (key_s0[87]), .Q (signal_16933) ) ;
    buf_clk cell_12053 ( .C (clk), .D (key_s1[87]), .Q (signal_16941) ) ;
    buf_clk cell_12061 ( .C (clk), .D (key_s0[88]), .Q (signal_16949) ) ;
    buf_clk cell_12069 ( .C (clk), .D (key_s1[88]), .Q (signal_16957) ) ;
    buf_clk cell_12077 ( .C (clk), .D (key_s0[89]), .Q (signal_16965) ) ;
    buf_clk cell_12085 ( .C (clk), .D (key_s1[89]), .Q (signal_16973) ) ;
    buf_clk cell_12093 ( .C (clk), .D (key_s0[90]), .Q (signal_16981) ) ;
    buf_clk cell_12101 ( .C (clk), .D (key_s1[90]), .Q (signal_16989) ) ;
    buf_clk cell_12109 ( .C (clk), .D (key_s0[91]), .Q (signal_16997) ) ;
    buf_clk cell_12117 ( .C (clk), .D (key_s1[91]), .Q (signal_17005) ) ;
    buf_clk cell_12125 ( .C (clk), .D (key_s0[92]), .Q (signal_17013) ) ;
    buf_clk cell_12133 ( .C (clk), .D (key_s1[92]), .Q (signal_17021) ) ;
    buf_clk cell_12141 ( .C (clk), .D (key_s0[93]), .Q (signal_17029) ) ;
    buf_clk cell_12149 ( .C (clk), .D (key_s1[93]), .Q (signal_17037) ) ;
    buf_clk cell_12157 ( .C (clk), .D (key_s0[94]), .Q (signal_17045) ) ;
    buf_clk cell_12165 ( .C (clk), .D (key_s1[94]), .Q (signal_17053) ) ;
    buf_clk cell_12173 ( .C (clk), .D (key_s0[95]), .Q (signal_17061) ) ;
    buf_clk cell_12181 ( .C (clk), .D (key_s1[95]), .Q (signal_17069) ) ;
    buf_clk cell_12189 ( .C (clk), .D (key_s0[96]), .Q (signal_17077) ) ;
    buf_clk cell_12197 ( .C (clk), .D (key_s1[96]), .Q (signal_17085) ) ;
    buf_clk cell_12205 ( .C (clk), .D (key_s0[97]), .Q (signal_17093) ) ;
    buf_clk cell_12213 ( .C (clk), .D (key_s1[97]), .Q (signal_17101) ) ;
    buf_clk cell_12221 ( .C (clk), .D (key_s0[98]), .Q (signal_17109) ) ;
    buf_clk cell_12229 ( .C (clk), .D (key_s1[98]), .Q (signal_17117) ) ;
    buf_clk cell_12237 ( .C (clk), .D (key_s0[99]), .Q (signal_17125) ) ;
    buf_clk cell_12245 ( .C (clk), .D (key_s1[99]), .Q (signal_17133) ) ;
    buf_clk cell_12253 ( .C (clk), .D (key_s0[100]), .Q (signal_17141) ) ;
    buf_clk cell_12261 ( .C (clk), .D (key_s1[100]), .Q (signal_17149) ) ;
    buf_clk cell_12269 ( .C (clk), .D (key_s0[101]), .Q (signal_17157) ) ;
    buf_clk cell_12277 ( .C (clk), .D (key_s1[101]), .Q (signal_17165) ) ;
    buf_clk cell_12285 ( .C (clk), .D (key_s0[102]), .Q (signal_17173) ) ;
    buf_clk cell_12293 ( .C (clk), .D (key_s1[102]), .Q (signal_17181) ) ;
    buf_clk cell_12301 ( .C (clk), .D (key_s0[103]), .Q (signal_17189) ) ;
    buf_clk cell_12309 ( .C (clk), .D (key_s1[103]), .Q (signal_17197) ) ;
    buf_clk cell_12317 ( .C (clk), .D (key_s0[104]), .Q (signal_17205) ) ;
    buf_clk cell_12325 ( .C (clk), .D (key_s1[104]), .Q (signal_17213) ) ;
    buf_clk cell_12333 ( .C (clk), .D (key_s0[105]), .Q (signal_17221) ) ;
    buf_clk cell_12341 ( .C (clk), .D (key_s1[105]), .Q (signal_17229) ) ;
    buf_clk cell_12349 ( .C (clk), .D (key_s0[106]), .Q (signal_17237) ) ;
    buf_clk cell_12357 ( .C (clk), .D (key_s1[106]), .Q (signal_17245) ) ;
    buf_clk cell_12365 ( .C (clk), .D (key_s0[107]), .Q (signal_17253) ) ;
    buf_clk cell_12373 ( .C (clk), .D (key_s1[107]), .Q (signal_17261) ) ;
    buf_clk cell_12381 ( .C (clk), .D (key_s0[108]), .Q (signal_17269) ) ;
    buf_clk cell_12389 ( .C (clk), .D (key_s1[108]), .Q (signal_17277) ) ;
    buf_clk cell_12397 ( .C (clk), .D (key_s0[109]), .Q (signal_17285) ) ;
    buf_clk cell_12405 ( .C (clk), .D (key_s1[109]), .Q (signal_17293) ) ;
    buf_clk cell_12413 ( .C (clk), .D (key_s0[110]), .Q (signal_17301) ) ;
    buf_clk cell_12421 ( .C (clk), .D (key_s1[110]), .Q (signal_17309) ) ;
    buf_clk cell_12429 ( .C (clk), .D (key_s0[111]), .Q (signal_17317) ) ;
    buf_clk cell_12437 ( .C (clk), .D (key_s1[111]), .Q (signal_17325) ) ;
    buf_clk cell_12445 ( .C (clk), .D (key_s0[112]), .Q (signal_17333) ) ;
    buf_clk cell_12453 ( .C (clk), .D (key_s1[112]), .Q (signal_17341) ) ;
    buf_clk cell_12461 ( .C (clk), .D (key_s0[113]), .Q (signal_17349) ) ;
    buf_clk cell_12469 ( .C (clk), .D (key_s1[113]), .Q (signal_17357) ) ;
    buf_clk cell_12477 ( .C (clk), .D (key_s0[114]), .Q (signal_17365) ) ;
    buf_clk cell_12485 ( .C (clk), .D (key_s1[114]), .Q (signal_17373) ) ;
    buf_clk cell_12493 ( .C (clk), .D (key_s0[115]), .Q (signal_17381) ) ;
    buf_clk cell_12501 ( .C (clk), .D (key_s1[115]), .Q (signal_17389) ) ;
    buf_clk cell_12509 ( .C (clk), .D (key_s0[116]), .Q (signal_17397) ) ;
    buf_clk cell_12517 ( .C (clk), .D (key_s1[116]), .Q (signal_17405) ) ;
    buf_clk cell_12525 ( .C (clk), .D (key_s0[117]), .Q (signal_17413) ) ;
    buf_clk cell_12533 ( .C (clk), .D (key_s1[117]), .Q (signal_17421) ) ;
    buf_clk cell_12541 ( .C (clk), .D (key_s0[118]), .Q (signal_17429) ) ;
    buf_clk cell_12549 ( .C (clk), .D (key_s1[118]), .Q (signal_17437) ) ;
    buf_clk cell_12557 ( .C (clk), .D (key_s0[119]), .Q (signal_17445) ) ;
    buf_clk cell_12565 ( .C (clk), .D (key_s1[119]), .Q (signal_17453) ) ;
    buf_clk cell_12573 ( .C (clk), .D (key_s0[120]), .Q (signal_17461) ) ;
    buf_clk cell_12581 ( .C (clk), .D (key_s1[120]), .Q (signal_17469) ) ;
    buf_clk cell_12589 ( .C (clk), .D (key_s0[121]), .Q (signal_17477) ) ;
    buf_clk cell_12597 ( .C (clk), .D (key_s1[121]), .Q (signal_17485) ) ;
    buf_clk cell_12605 ( .C (clk), .D (key_s0[122]), .Q (signal_17493) ) ;
    buf_clk cell_12613 ( .C (clk), .D (key_s1[122]), .Q (signal_17501) ) ;
    buf_clk cell_12621 ( .C (clk), .D (key_s0[123]), .Q (signal_17509) ) ;
    buf_clk cell_12629 ( .C (clk), .D (key_s1[123]), .Q (signal_17517) ) ;
    buf_clk cell_12637 ( .C (clk), .D (key_s0[124]), .Q (signal_17525) ) ;
    buf_clk cell_12645 ( .C (clk), .D (key_s1[124]), .Q (signal_17533) ) ;
    buf_clk cell_12653 ( .C (clk), .D (key_s0[125]), .Q (signal_17541) ) ;
    buf_clk cell_12661 ( .C (clk), .D (key_s1[125]), .Q (signal_17549) ) ;
    buf_clk cell_12669 ( .C (clk), .D (key_s0[126]), .Q (signal_17557) ) ;
    buf_clk cell_12677 ( .C (clk), .D (key_s1[126]), .Q (signal_17565) ) ;
    buf_clk cell_12685 ( .C (clk), .D (key_s0[127]), .Q (signal_17573) ) ;
    buf_clk cell_12693 ( .C (clk), .D (key_s1[127]), .Q (signal_17581) ) ;
    buf_clk cell_12701 ( .C (clk), .D (signal_4347), .Q (signal_17589) ) ;
    buf_clk cell_12709 ( .C (clk), .D (signal_7661), .Q (signal_17597) ) ;
    buf_clk cell_12717 ( .C (clk), .D (signal_4315), .Q (signal_17605) ) ;
    buf_clk cell_12725 ( .C (clk), .D (signal_7503), .Q (signal_17613) ) ;
    buf_clk cell_12733 ( .C (clk), .D (signal_4283), .Q (signal_17621) ) ;
    buf_clk cell_12741 ( .C (clk), .D (signal_7527), .Q (signal_17629) ) ;
    buf_clk cell_12749 ( .C (clk), .D (signal_4348), .Q (signal_17637) ) ;
    buf_clk cell_12757 ( .C (clk), .D (signal_7658), .Q (signal_17645) ) ;
    buf_clk cell_12765 ( .C (clk), .D (signal_4316), .Q (signal_17653) ) ;
    buf_clk cell_12773 ( .C (clk), .D (signal_7500), .Q (signal_17661) ) ;
    buf_clk cell_12781 ( .C (clk), .D (signal_4284), .Q (signal_17669) ) ;
    buf_clk cell_12789 ( .C (clk), .D (signal_7524), .Q (signal_17677) ) ;
    buf_clk cell_12797 ( .C (clk), .D (signal_4349), .Q (signal_17685) ) ;
    buf_clk cell_12805 ( .C (clk), .D (signal_7652), .Q (signal_17693) ) ;
    buf_clk cell_12813 ( .C (clk), .D (signal_4317), .Q (signal_17701) ) ;
    buf_clk cell_12821 ( .C (clk), .D (signal_7497), .Q (signal_17709) ) ;
    buf_clk cell_12829 ( .C (clk), .D (signal_4285), .Q (signal_17717) ) ;
    buf_clk cell_12837 ( .C (clk), .D (signal_7521), .Q (signal_17725) ) ;
    buf_clk cell_12845 ( .C (clk), .D (signal_4350), .Q (signal_17733) ) ;
    buf_clk cell_12853 ( .C (clk), .D (signal_7649), .Q (signal_17741) ) ;
    buf_clk cell_12861 ( .C (clk), .D (signal_4318), .Q (signal_17749) ) ;
    buf_clk cell_12869 ( .C (clk), .D (signal_7494), .Q (signal_17757) ) ;
    buf_clk cell_12877 ( .C (clk), .D (signal_4286), .Q (signal_17765) ) ;
    buf_clk cell_12885 ( .C (clk), .D (signal_7518), .Q (signal_17773) ) ;
    buf_clk cell_12893 ( .C (clk), .D (signal_4351), .Q (signal_17781) ) ;
    buf_clk cell_12901 ( .C (clk), .D (signal_7646), .Q (signal_17789) ) ;
    buf_clk cell_12909 ( .C (clk), .D (signal_4319), .Q (signal_17797) ) ;
    buf_clk cell_12917 ( .C (clk), .D (signal_7491), .Q (signal_17805) ) ;
    buf_clk cell_12925 ( .C (clk), .D (signal_4287), .Q (signal_17813) ) ;
    buf_clk cell_12933 ( .C (clk), .D (signal_7515), .Q (signal_17821) ) ;
    buf_clk cell_12941 ( .C (clk), .D (signal_4352), .Q (signal_17829) ) ;
    buf_clk cell_12949 ( .C (clk), .D (signal_7643), .Q (signal_17837) ) ;
    buf_clk cell_12957 ( .C (clk), .D (signal_4320), .Q (signal_17845) ) ;
    buf_clk cell_12965 ( .C (clk), .D (signal_7488), .Q (signal_17853) ) ;
    buf_clk cell_12973 ( .C (clk), .D (signal_4288), .Q (signal_17861) ) ;
    buf_clk cell_12981 ( .C (clk), .D (signal_7512), .Q (signal_17869) ) ;
    buf_clk cell_12989 ( .C (clk), .D (signal_4353), .Q (signal_17877) ) ;
    buf_clk cell_12997 ( .C (clk), .D (signal_7640), .Q (signal_17885) ) ;
    buf_clk cell_13005 ( .C (clk), .D (signal_4321), .Q (signal_17893) ) ;
    buf_clk cell_13013 ( .C (clk), .D (signal_7485), .Q (signal_17901) ) ;
    buf_clk cell_13021 ( .C (clk), .D (signal_4289), .Q (signal_17909) ) ;
    buf_clk cell_13029 ( .C (clk), .D (signal_7509), .Q (signal_17917) ) ;
    buf_clk cell_13037 ( .C (clk), .D (signal_4354), .Q (signal_17925) ) ;
    buf_clk cell_13045 ( .C (clk), .D (signal_7637), .Q (signal_17933) ) ;
    buf_clk cell_13053 ( .C (clk), .D (signal_4322), .Q (signal_17941) ) ;
    buf_clk cell_13061 ( .C (clk), .D (signal_7482), .Q (signal_17949) ) ;
    buf_clk cell_13069 ( .C (clk), .D (signal_4290), .Q (signal_17957) ) ;
    buf_clk cell_13077 ( .C (clk), .D (signal_7506), .Q (signal_17965) ) ;
    buf_clk cell_13085 ( .C (clk), .D (signal_4251), .Q (signal_17973) ) ;
    buf_clk cell_13093 ( .C (clk), .D (signal_7479), .Q (signal_17981) ) ;
    buf_clk cell_13101 ( .C (clk), .D (signal_4252), .Q (signal_17989) ) ;
    buf_clk cell_13109 ( .C (clk), .D (signal_7476), .Q (signal_17997) ) ;
    buf_clk cell_13117 ( .C (clk), .D (signal_4253), .Q (signal_18005) ) ;
    buf_clk cell_13125 ( .C (clk), .D (signal_7473), .Q (signal_18013) ) ;
    buf_clk cell_13133 ( .C (clk), .D (signal_4254), .Q (signal_18021) ) ;
    buf_clk cell_13141 ( .C (clk), .D (signal_7470), .Q (signal_18029) ) ;
    buf_clk cell_13149 ( .C (clk), .D (signal_4255), .Q (signal_18037) ) ;
    buf_clk cell_13157 ( .C (clk), .D (signal_7467), .Q (signal_18045) ) ;
    buf_clk cell_13165 ( .C (clk), .D (signal_4256), .Q (signal_18053) ) ;
    buf_clk cell_13173 ( .C (clk), .D (signal_7464), .Q (signal_18061) ) ;
    buf_clk cell_13181 ( .C (clk), .D (signal_4257), .Q (signal_18069) ) ;
    buf_clk cell_13189 ( .C (clk), .D (signal_7461), .Q (signal_18077) ) ;
    buf_clk cell_13197 ( .C (clk), .D (signal_4258), .Q (signal_18085) ) ;
    buf_clk cell_13205 ( .C (clk), .D (signal_7458), .Q (signal_18093) ) ;
    buf_clk cell_13213 ( .C (clk), .D (signal_393), .Q (signal_18101) ) ;
    buf_clk cell_13221 ( .C (clk), .D (signal_394), .Q (signal_18109) ) ;
    buf_clk cell_13229 ( .C (clk), .D (signal_4379), .Q (signal_18117) ) ;
    buf_clk cell_13237 ( .C (clk), .D (signal_4380), .Q (signal_18125) ) ;
    buf_clk cell_13245 ( .C (clk), .D (signal_4381), .Q (signal_18133) ) ;
    buf_clk cell_13253 ( .C (clk), .D (signal_4382), .Q (signal_18141) ) ;
    buf_clk cell_13261 ( .C (clk), .D (signal_4383), .Q (signal_18149) ) ;
    buf_clk cell_13269 ( .C (clk), .D (signal_4384), .Q (signal_18157) ) ;
    buf_clk cell_13277 ( .C (clk), .D (signal_4903), .Q (signal_18165) ) ;
    buf_clk cell_13283 ( .C (clk), .D (signal_8271), .Q (signal_18171) ) ;
    buf_clk cell_13289 ( .C (clk), .D (ciphertext_s0[56]), .Q (signal_18177) ) ;
    buf_clk cell_13295 ( .C (clk), .D (ciphertext_s1[56]), .Q (signal_18183) ) ;
    buf_clk cell_13301 ( .C (clk), .D (signal_4690), .Q (signal_18189) ) ;
    buf_clk cell_13307 ( .C (clk), .D (signal_8074), .Q (signal_18195) ) ;
    buf_clk cell_13313 ( .C (clk), .D (signal_4906), .Q (signal_18201) ) ;
    buf_clk cell_13319 ( .C (clk), .D (signal_8274), .Q (signal_18207) ) ;
    buf_clk cell_13325 ( .C (clk), .D (signal_4908), .Q (signal_18213) ) ;
    buf_clk cell_13331 ( .C (clk), .D (signal_8276), .Q (signal_18219) ) ;
    buf_clk cell_13337 ( .C (clk), .D (signal_4694), .Q (signal_18225) ) ;
    buf_clk cell_13343 ( .C (clk), .D (signal_8078), .Q (signal_18231) ) ;
    buf_clk cell_13349 ( .C (clk), .D (signal_4695), .Q (signal_18237) ) ;
    buf_clk cell_13355 ( .C (clk), .D (signal_8079), .Q (signal_18243) ) ;
    buf_clk cell_13361 ( .C (clk), .D (signal_4907), .Q (signal_18249) ) ;
    buf_clk cell_13367 ( .C (clk), .D (signal_8275), .Q (signal_18255) ) ;
    buf_clk cell_13373 ( .C (clk), .D (signal_4934), .Q (signal_18261) ) ;
    buf_clk cell_13379 ( .C (clk), .D (signal_8278), .Q (signal_18267) ) ;
    buf_clk cell_13385 ( .C (clk), .D (ciphertext_s0[88]), .Q (signal_18273) ) ;
    buf_clk cell_13391 ( .C (clk), .D (ciphertext_s1[88]), .Q (signal_18279) ) ;
    buf_clk cell_13397 ( .C (clk), .D (signal_4728), .Q (signal_18285) ) ;
    buf_clk cell_13403 ( .C (clk), .D (signal_8082), .Q (signal_18291) ) ;
    buf_clk cell_13409 ( .C (clk), .D (signal_4937), .Q (signal_18297) ) ;
    buf_clk cell_13415 ( .C (clk), .D (signal_8281), .Q (signal_18303) ) ;
    buf_clk cell_13421 ( .C (clk), .D (signal_4939), .Q (signal_18309) ) ;
    buf_clk cell_13427 ( .C (clk), .D (signal_8283), .Q (signal_18315) ) ;
    buf_clk cell_13433 ( .C (clk), .D (signal_4732), .Q (signal_18321) ) ;
    buf_clk cell_13439 ( .C (clk), .D (signal_8086), .Q (signal_18327) ) ;
    buf_clk cell_13445 ( .C (clk), .D (signal_4733), .Q (signal_18333) ) ;
    buf_clk cell_13451 ( .C (clk), .D (signal_8087), .Q (signal_18339) ) ;
    buf_clk cell_13457 ( .C (clk), .D (signal_4938), .Q (signal_18345) ) ;
    buf_clk cell_13463 ( .C (clk), .D (signal_8282), .Q (signal_18351) ) ;
    buf_clk cell_13469 ( .C (clk), .D (signal_4965), .Q (signal_18357) ) ;
    buf_clk cell_13475 ( .C (clk), .D (signal_8285), .Q (signal_18363) ) ;
    buf_clk cell_13481 ( .C (clk), .D (ciphertext_s0[120]), .Q (signal_18369) ) ;
    buf_clk cell_13487 ( .C (clk), .D (ciphertext_s1[120]), .Q (signal_18375) ) ;
    buf_clk cell_13493 ( .C (clk), .D (signal_4766), .Q (signal_18381) ) ;
    buf_clk cell_13499 ( .C (clk), .D (signal_8090), .Q (signal_18387) ) ;
    buf_clk cell_13505 ( .C (clk), .D (signal_4968), .Q (signal_18393) ) ;
    buf_clk cell_13511 ( .C (clk), .D (signal_8288), .Q (signal_18399) ) ;
    buf_clk cell_13517 ( .C (clk), .D (signal_4970), .Q (signal_18405) ) ;
    buf_clk cell_13523 ( .C (clk), .D (signal_8290), .Q (signal_18411) ) ;
    buf_clk cell_13529 ( .C (clk), .D (signal_4770), .Q (signal_18417) ) ;
    buf_clk cell_13535 ( .C (clk), .D (signal_8094), .Q (signal_18423) ) ;
    buf_clk cell_13541 ( .C (clk), .D (signal_4771), .Q (signal_18429) ) ;
    buf_clk cell_13547 ( .C (clk), .D (signal_8095), .Q (signal_18435) ) ;
    buf_clk cell_13553 ( .C (clk), .D (signal_4969), .Q (signal_18441) ) ;
    buf_clk cell_13559 ( .C (clk), .D (signal_8289), .Q (signal_18447) ) ;
    buf_clk cell_13565 ( .C (clk), .D (signal_4972), .Q (signal_18453) ) ;
    buf_clk cell_13571 ( .C (clk), .D (signal_8225), .Q (signal_18459) ) ;
    buf_clk cell_13577 ( .C (clk), .D (signal_4362), .Q (signal_18465) ) ;
    buf_clk cell_13583 ( .C (clk), .D (signal_7610), .Q (signal_18471) ) ;
    buf_clk cell_13589 ( .C (clk), .D (signal_4774), .Q (signal_18477) ) ;
    buf_clk cell_13595 ( .C (clk), .D (signal_8042), .Q (signal_18483) ) ;
    buf_clk cell_13601 ( .C (clk), .D (signal_4975), .Q (signal_18489) ) ;
    buf_clk cell_13607 ( .C (clk), .D (signal_8228), .Q (signal_18495) ) ;
    buf_clk cell_13613 ( .C (clk), .D (signal_4977), .Q (signal_18501) ) ;
    buf_clk cell_13619 ( .C (clk), .D (signal_8230), .Q (signal_18507) ) ;
    buf_clk cell_13625 ( .C (clk), .D (signal_4778), .Q (signal_18513) ) ;
    buf_clk cell_13631 ( .C (clk), .D (signal_8046), .Q (signal_18519) ) ;
    buf_clk cell_13637 ( .C (clk), .D (signal_4779), .Q (signal_18525) ) ;
    buf_clk cell_13643 ( .C (clk), .D (signal_8047), .Q (signal_18531) ) ;
    buf_clk cell_13649 ( .C (clk), .D (signal_4976), .Q (signal_18537) ) ;
    buf_clk cell_13655 ( .C (clk), .D (signal_8229), .Q (signal_18543) ) ;
    buf_clk cell_13661 ( .C (clk), .D (signal_4979), .Q (signal_18549) ) ;
    buf_clk cell_13667 ( .C (clk), .D (signal_8232), .Q (signal_18555) ) ;
    buf_clk cell_13673 ( .C (clk), .D (signal_4370), .Q (signal_18561) ) ;
    buf_clk cell_13679 ( .C (clk), .D (signal_7823), .Q (signal_18567) ) ;
    buf_clk cell_13685 ( .C (clk), .D (signal_4782), .Q (signal_18573) ) ;
    buf_clk cell_13691 ( .C (clk), .D (signal_8050), .Q (signal_18579) ) ;
    buf_clk cell_13697 ( .C (clk), .D (signal_4982), .Q (signal_18585) ) ;
    buf_clk cell_13703 ( .C (clk), .D (signal_8235), .Q (signal_18591) ) ;
    buf_clk cell_13709 ( .C (clk), .D (signal_4984), .Q (signal_18597) ) ;
    buf_clk cell_13715 ( .C (clk), .D (signal_8237), .Q (signal_18603) ) ;
    buf_clk cell_13721 ( .C (clk), .D (signal_4786), .Q (signal_18609) ) ;
    buf_clk cell_13727 ( .C (clk), .D (signal_8054), .Q (signal_18615) ) ;
    buf_clk cell_13733 ( .C (clk), .D (signal_4787), .Q (signal_18621) ) ;
    buf_clk cell_13739 ( .C (clk), .D (signal_8055), .Q (signal_18627) ) ;
    buf_clk cell_13745 ( .C (clk), .D (signal_4983), .Q (signal_18633) ) ;
    buf_clk cell_13751 ( .C (clk), .D (signal_8236), .Q (signal_18639) ) ;
    buf_clk cell_13757 ( .C (clk), .D (signal_4986), .Q (signal_18645) ) ;
    buf_clk cell_13763 ( .C (clk), .D (signal_8239), .Q (signal_18651) ) ;
    buf_clk cell_13769 ( .C (clk), .D (signal_4378), .Q (signal_18657) ) ;
    buf_clk cell_13775 ( .C (clk), .D (signal_7529), .Q (signal_18663) ) ;
    buf_clk cell_13781 ( .C (clk), .D (signal_4790), .Q (signal_18669) ) ;
    buf_clk cell_13787 ( .C (clk), .D (signal_8058), .Q (signal_18675) ) ;
    buf_clk cell_13793 ( .C (clk), .D (signal_4989), .Q (signal_18681) ) ;
    buf_clk cell_13799 ( .C (clk), .D (signal_8242), .Q (signal_18687) ) ;
    buf_clk cell_13805 ( .C (clk), .D (signal_4991), .Q (signal_18693) ) ;
    buf_clk cell_13811 ( .C (clk), .D (signal_8244), .Q (signal_18699) ) ;
    buf_clk cell_13817 ( .C (clk), .D (signal_4794), .Q (signal_18705) ) ;
    buf_clk cell_13823 ( .C (clk), .D (signal_8062), .Q (signal_18711) ) ;
    buf_clk cell_13829 ( .C (clk), .D (signal_4795), .Q (signal_18717) ) ;
    buf_clk cell_13835 ( .C (clk), .D (signal_8063), .Q (signal_18723) ) ;
    buf_clk cell_13841 ( .C (clk), .D (signal_4990), .Q (signal_18729) ) ;
    buf_clk cell_13847 ( .C (clk), .D (signal_8243), .Q (signal_18735) ) ;
    buf_clk cell_13853 ( .C (clk), .D (signal_4993), .Q (signal_18741) ) ;
    buf_clk cell_13859 ( .C (clk), .D (signal_8246), .Q (signal_18747) ) ;
    buf_clk cell_13865 ( .C (clk), .D (signal_4798), .Q (signal_18753) ) ;
    buf_clk cell_13871 ( .C (clk), .D (signal_8066), .Q (signal_18759) ) ;
    buf_clk cell_13877 ( .C (clk), .D (signal_4996), .Q (signal_18765) ) ;
    buf_clk cell_13883 ( .C (clk), .D (signal_8249), .Q (signal_18771) ) ;
    buf_clk cell_13889 ( .C (clk), .D (signal_4998), .Q (signal_18777) ) ;
    buf_clk cell_13895 ( .C (clk), .D (signal_8251), .Q (signal_18783) ) ;
    buf_clk cell_13901 ( .C (clk), .D (signal_4802), .Q (signal_18789) ) ;
    buf_clk cell_13907 ( .C (clk), .D (signal_8070), .Q (signal_18795) ) ;
    buf_clk cell_13913 ( .C (clk), .D (signal_4803), .Q (signal_18801) ) ;
    buf_clk cell_13919 ( .C (clk), .D (signal_8071), .Q (signal_18807) ) ;
    buf_clk cell_13925 ( .C (clk), .D (signal_4997), .Q (signal_18813) ) ;
    buf_clk cell_13931 ( .C (clk), .D (signal_8250), .Q (signal_18819) ) ;
    buf_clk cell_13937 ( .C (clk), .D (signal_5099), .Q (signal_18825) ) ;
    buf_clk cell_13943 ( .C (clk), .D (signal_8382), .Q (signal_18831) ) ;
    buf_clk cell_13949 ( .C (clk), .D (ciphertext_s0[0]), .Q (signal_18837) ) ;
    buf_clk cell_13955 ( .C (clk), .D (ciphertext_s1[0]), .Q (signal_18843) ) ;
    buf_clk cell_13961 ( .C (clk), .D (signal_4848), .Q (signal_18849) ) ;
    buf_clk cell_13967 ( .C (clk), .D (signal_8122), .Q (signal_18855) ) ;
    buf_clk cell_13973 ( .C (clk), .D (signal_5102), .Q (signal_18861) ) ;
    buf_clk cell_13979 ( .C (clk), .D (signal_8385), .Q (signal_18867) ) ;
    buf_clk cell_13985 ( .C (clk), .D (signal_5104), .Q (signal_18873) ) ;
    buf_clk cell_13991 ( .C (clk), .D (signal_8387), .Q (signal_18879) ) ;
    buf_clk cell_13997 ( .C (clk), .D (signal_4852), .Q (signal_18885) ) ;
    buf_clk cell_14003 ( .C (clk), .D (signal_8126), .Q (signal_18891) ) ;
    buf_clk cell_14009 ( .C (clk), .D (signal_4853), .Q (signal_18897) ) ;
    buf_clk cell_14015 ( .C (clk), .D (signal_8127), .Q (signal_18903) ) ;
    buf_clk cell_14021 ( .C (clk), .D (signal_5103), .Q (signal_18909) ) ;
    buf_clk cell_14027 ( .C (clk), .D (signal_8386), .Q (signal_18915) ) ;
    buf_clk cell_14033 ( .C (clk), .D (signal_5106), .Q (signal_18921) ) ;
    buf_clk cell_14039 ( .C (clk), .D (signal_8389), .Q (signal_18927) ) ;
    buf_clk cell_14045 ( .C (clk), .D (ciphertext_s0[8]), .Q (signal_18933) ) ;
    buf_clk cell_14051 ( .C (clk), .D (ciphertext_s1[8]), .Q (signal_18939) ) ;
    buf_clk cell_14057 ( .C (clk), .D (signal_4856), .Q (signal_18945) ) ;
    buf_clk cell_14063 ( .C (clk), .D (signal_8130), .Q (signal_18951) ) ;
    buf_clk cell_14069 ( .C (clk), .D (signal_5109), .Q (signal_18957) ) ;
    buf_clk cell_14075 ( .C (clk), .D (signal_8392), .Q (signal_18963) ) ;
    buf_clk cell_14081 ( .C (clk), .D (signal_5111), .Q (signal_18969) ) ;
    buf_clk cell_14087 ( .C (clk), .D (signal_8394), .Q (signal_18975) ) ;
    buf_clk cell_14093 ( .C (clk), .D (signal_4860), .Q (signal_18981) ) ;
    buf_clk cell_14099 ( .C (clk), .D (signal_8134), .Q (signal_18987) ) ;
    buf_clk cell_14105 ( .C (clk), .D (signal_4861), .Q (signal_18993) ) ;
    buf_clk cell_14111 ( .C (clk), .D (signal_8135), .Q (signal_18999) ) ;
    buf_clk cell_14117 ( .C (clk), .D (signal_5110), .Q (signal_19005) ) ;
    buf_clk cell_14123 ( .C (clk), .D (signal_8393), .Q (signal_19011) ) ;
    buf_clk cell_14129 ( .C (clk), .D (signal_5113), .Q (signal_19017) ) ;
    buf_clk cell_14135 ( .C (clk), .D (signal_8396), .Q (signal_19023) ) ;
    buf_clk cell_14141 ( .C (clk), .D (ciphertext_s0[16]), .Q (signal_19029) ) ;
    buf_clk cell_14147 ( .C (clk), .D (ciphertext_s1[16]), .Q (signal_19035) ) ;
    buf_clk cell_14153 ( .C (clk), .D (signal_4864), .Q (signal_19041) ) ;
    buf_clk cell_14159 ( .C (clk), .D (signal_8138), .Q (signal_19047) ) ;
    buf_clk cell_14165 ( .C (clk), .D (signal_5116), .Q (signal_19053) ) ;
    buf_clk cell_14171 ( .C (clk), .D (signal_8399), .Q (signal_19059) ) ;
    buf_clk cell_14177 ( .C (clk), .D (signal_5118), .Q (signal_19065) ) ;
    buf_clk cell_14183 ( .C (clk), .D (signal_8401), .Q (signal_19071) ) ;
    buf_clk cell_14189 ( .C (clk), .D (signal_4868), .Q (signal_19077) ) ;
    buf_clk cell_14195 ( .C (clk), .D (signal_8142), .Q (signal_19083) ) ;
    buf_clk cell_14201 ( .C (clk), .D (signal_4869), .Q (signal_19089) ) ;
    buf_clk cell_14207 ( .C (clk), .D (signal_8143), .Q (signal_19095) ) ;
    buf_clk cell_14213 ( .C (clk), .D (signal_5117), .Q (signal_19101) ) ;
    buf_clk cell_14219 ( .C (clk), .D (signal_8400), .Q (signal_19107) ) ;
    buf_clk cell_14225 ( .C (clk), .D (signal_5120), .Q (signal_19113) ) ;
    buf_clk cell_14231 ( .C (clk), .D (signal_8403), .Q (signal_19119) ) ;
    buf_clk cell_14237 ( .C (clk), .D (ciphertext_s0[24]), .Q (signal_19125) ) ;
    buf_clk cell_14243 ( .C (clk), .D (ciphertext_s1[24]), .Q (signal_19131) ) ;
    buf_clk cell_14249 ( .C (clk), .D (signal_4872), .Q (signal_19137) ) ;
    buf_clk cell_14255 ( .C (clk), .D (signal_8146), .Q (signal_19143) ) ;
    buf_clk cell_14261 ( .C (clk), .D (signal_5123), .Q (signal_19149) ) ;
    buf_clk cell_14267 ( .C (clk), .D (signal_8406), .Q (signal_19155) ) ;
    buf_clk cell_14273 ( .C (clk), .D (signal_5125), .Q (signal_19161) ) ;
    buf_clk cell_14279 ( .C (clk), .D (signal_8408), .Q (signal_19167) ) ;
    buf_clk cell_14285 ( .C (clk), .D (signal_4876), .Q (signal_19173) ) ;
    buf_clk cell_14291 ( .C (clk), .D (signal_8150), .Q (signal_19179) ) ;
    buf_clk cell_14297 ( .C (clk), .D (signal_4877), .Q (signal_19185) ) ;
    buf_clk cell_14303 ( .C (clk), .D (signal_8151), .Q (signal_19191) ) ;
    buf_clk cell_14309 ( .C (clk), .D (signal_5124), .Q (signal_19197) ) ;
    buf_clk cell_14315 ( .C (clk), .D (signal_8407), .Q (signal_19203) ) ;
    buf_clk cell_14321 ( .C (clk), .D (signal_5127), .Q (signal_19209) ) ;
    buf_clk cell_14327 ( .C (clk), .D (signal_8410), .Q (signal_19215) ) ;
    buf_clk cell_14333 ( .C (clk), .D (ciphertext_s0[32]), .Q (signal_19221) ) ;
    buf_clk cell_14339 ( .C (clk), .D (ciphertext_s1[32]), .Q (signal_19227) ) ;
    buf_clk cell_14345 ( .C (clk), .D (signal_4880), .Q (signal_19233) ) ;
    buf_clk cell_14351 ( .C (clk), .D (signal_8154), .Q (signal_19239) ) ;
    buf_clk cell_14357 ( .C (clk), .D (signal_5130), .Q (signal_19245) ) ;
    buf_clk cell_14363 ( .C (clk), .D (signal_8413), .Q (signal_19251) ) ;
    buf_clk cell_14369 ( .C (clk), .D (signal_5132), .Q (signal_19257) ) ;
    buf_clk cell_14375 ( .C (clk), .D (signal_8415), .Q (signal_19263) ) ;
    buf_clk cell_14381 ( .C (clk), .D (signal_4884), .Q (signal_19269) ) ;
    buf_clk cell_14387 ( .C (clk), .D (signal_8158), .Q (signal_19275) ) ;
    buf_clk cell_14393 ( .C (clk), .D (signal_4885), .Q (signal_19281) ) ;
    buf_clk cell_14399 ( .C (clk), .D (signal_8159), .Q (signal_19287) ) ;
    buf_clk cell_14405 ( .C (clk), .D (signal_5131), .Q (signal_19293) ) ;
    buf_clk cell_14411 ( .C (clk), .D (signal_8414), .Q (signal_19299) ) ;
    buf_clk cell_14417 ( .C (clk), .D (signal_5134), .Q (signal_19305) ) ;
    buf_clk cell_14423 ( .C (clk), .D (signal_8417), .Q (signal_19311) ) ;
    buf_clk cell_14429 ( .C (clk), .D (ciphertext_s0[40]), .Q (signal_19317) ) ;
    buf_clk cell_14435 ( .C (clk), .D (ciphertext_s1[40]), .Q (signal_19323) ) ;
    buf_clk cell_14441 ( .C (clk), .D (signal_4888), .Q (signal_19329) ) ;
    buf_clk cell_14447 ( .C (clk), .D (signal_8162), .Q (signal_19335) ) ;
    buf_clk cell_14453 ( .C (clk), .D (signal_5137), .Q (signal_19341) ) ;
    buf_clk cell_14459 ( .C (clk), .D (signal_8420), .Q (signal_19347) ) ;
    buf_clk cell_14465 ( .C (clk), .D (signal_5139), .Q (signal_19353) ) ;
    buf_clk cell_14471 ( .C (clk), .D (signal_8422), .Q (signal_19359) ) ;
    buf_clk cell_14477 ( .C (clk), .D (signal_4892), .Q (signal_19365) ) ;
    buf_clk cell_14483 ( .C (clk), .D (signal_8166), .Q (signal_19371) ) ;
    buf_clk cell_14489 ( .C (clk), .D (signal_4893), .Q (signal_19377) ) ;
    buf_clk cell_14495 ( .C (clk), .D (signal_8167), .Q (signal_19383) ) ;
    buf_clk cell_14501 ( .C (clk), .D (signal_5138), .Q (signal_19389) ) ;
    buf_clk cell_14507 ( .C (clk), .D (signal_8421), .Q (signal_19395) ) ;
    buf_clk cell_14513 ( .C (clk), .D (signal_5141), .Q (signal_19401) ) ;
    buf_clk cell_14519 ( .C (clk), .D (signal_8424), .Q (signal_19407) ) ;
    buf_clk cell_14525 ( .C (clk), .D (ciphertext_s0[48]), .Q (signal_19413) ) ;
    buf_clk cell_14531 ( .C (clk), .D (ciphertext_s1[48]), .Q (signal_19419) ) ;
    buf_clk cell_14537 ( .C (clk), .D (signal_4896), .Q (signal_19425) ) ;
    buf_clk cell_14543 ( .C (clk), .D (signal_8170), .Q (signal_19431) ) ;
    buf_clk cell_14549 ( .C (clk), .D (signal_5144), .Q (signal_19437) ) ;
    buf_clk cell_14555 ( .C (clk), .D (signal_8427), .Q (signal_19443) ) ;
    buf_clk cell_14561 ( .C (clk), .D (signal_5146), .Q (signal_19449) ) ;
    buf_clk cell_14567 ( .C (clk), .D (signal_8429), .Q (signal_19455) ) ;
    buf_clk cell_14573 ( .C (clk), .D (signal_4900), .Q (signal_19461) ) ;
    buf_clk cell_14579 ( .C (clk), .D (signal_8174), .Q (signal_19467) ) ;
    buf_clk cell_14585 ( .C (clk), .D (signal_4901), .Q (signal_19473) ) ;
    buf_clk cell_14591 ( .C (clk), .D (signal_8175), .Q (signal_19479) ) ;
    buf_clk cell_14597 ( .C (clk), .D (signal_5145), .Q (signal_19485) ) ;
    buf_clk cell_14603 ( .C (clk), .D (signal_8428), .Q (signal_19491) ) ;
    buf_clk cell_14609 ( .C (clk), .D (signal_4689), .Q (signal_19497) ) ;
    buf_clk cell_14615 ( .C (clk), .D (signal_8073), .Q (signal_19503) ) ;
    buf_clk cell_14621 ( .C (clk), .D (signal_4693), .Q (signal_19509) ) ;
    buf_clk cell_14627 ( .C (clk), .D (signal_8077), .Q (signal_19515) ) ;
    buf_clk cell_14633 ( .C (clk), .D (signal_4692), .Q (signal_19521) ) ;
    buf_clk cell_14639 ( .C (clk), .D (signal_8076), .Q (signal_19527) ) ;
    buf_clk cell_14645 ( .C (clk), .D (signal_4904), .Q (signal_19533) ) ;
    buf_clk cell_14651 ( .C (clk), .D (signal_8272), .Q (signal_19539) ) ;
    buf_clk cell_14657 ( .C (clk), .D (signal_4691), .Q (signal_19545) ) ;
    buf_clk cell_14663 ( .C (clk), .D (signal_8075), .Q (signal_19551) ) ;
    buf_clk cell_14669 ( .C (clk), .D (signal_4551), .Q (signal_19557) ) ;
    buf_clk cell_14675 ( .C (clk), .D (signal_7883), .Q (signal_19563) ) ;
    buf_clk cell_14681 ( .C (clk), .D (signal_4549), .Q (signal_19569) ) ;
    buf_clk cell_14687 ( .C (clk), .D (signal_7881), .Q (signal_19575) ) ;
    buf_clk cell_14693 ( .C (clk), .D (signal_4550), .Q (signal_19581) ) ;
    buf_clk cell_14699 ( .C (clk), .D (signal_7882), .Q (signal_19587) ) ;
    buf_clk cell_14705 ( .C (clk), .D (signal_5154), .Q (signal_19593) ) ;
    buf_clk cell_14711 ( .C (clk), .D (signal_8431), .Q (signal_19599) ) ;
    buf_clk cell_14717 ( .C (clk), .D (ciphertext_s0[64]), .Q (signal_19605) ) ;
    buf_clk cell_14723 ( .C (clk), .D (ciphertext_s1[64]), .Q (signal_19611) ) ;
    buf_clk cell_14729 ( .C (clk), .D (signal_4911), .Q (signal_19617) ) ;
    buf_clk cell_14735 ( .C (clk), .D (signal_8178), .Q (signal_19623) ) ;
    buf_clk cell_14741 ( .C (clk), .D (signal_5157), .Q (signal_19629) ) ;
    buf_clk cell_14747 ( .C (clk), .D (signal_8434), .Q (signal_19635) ) ;
    buf_clk cell_14753 ( .C (clk), .D (signal_5159), .Q (signal_19641) ) ;
    buf_clk cell_14759 ( .C (clk), .D (signal_8436), .Q (signal_19647) ) ;
    buf_clk cell_14765 ( .C (clk), .D (signal_4915), .Q (signal_19653) ) ;
    buf_clk cell_14771 ( .C (clk), .D (signal_8182), .Q (signal_19659) ) ;
    buf_clk cell_14777 ( .C (clk), .D (signal_4916), .Q (signal_19665) ) ;
    buf_clk cell_14783 ( .C (clk), .D (signal_8183), .Q (signal_19671) ) ;
    buf_clk cell_14789 ( .C (clk), .D (signal_5158), .Q (signal_19677) ) ;
    buf_clk cell_14795 ( .C (clk), .D (signal_8435), .Q (signal_19683) ) ;
    buf_clk cell_14801 ( .C (clk), .D (signal_5161), .Q (signal_19689) ) ;
    buf_clk cell_14807 ( .C (clk), .D (signal_8438), .Q (signal_19695) ) ;
    buf_clk cell_14813 ( .C (clk), .D (ciphertext_s0[72]), .Q (signal_19701) ) ;
    buf_clk cell_14819 ( .C (clk), .D (ciphertext_s1[72]), .Q (signal_19707) ) ;
    buf_clk cell_14825 ( .C (clk), .D (signal_4919), .Q (signal_19713) ) ;
    buf_clk cell_14831 ( .C (clk), .D (signal_8186), .Q (signal_19719) ) ;
    buf_clk cell_14837 ( .C (clk), .D (signal_5164), .Q (signal_19725) ) ;
    buf_clk cell_14843 ( .C (clk), .D (signal_8441), .Q (signal_19731) ) ;
    buf_clk cell_14849 ( .C (clk), .D (signal_5166), .Q (signal_19737) ) ;
    buf_clk cell_14855 ( .C (clk), .D (signal_8443), .Q (signal_19743) ) ;
    buf_clk cell_14861 ( .C (clk), .D (signal_4923), .Q (signal_19749) ) ;
    buf_clk cell_14867 ( .C (clk), .D (signal_8190), .Q (signal_19755) ) ;
    buf_clk cell_14873 ( .C (clk), .D (signal_4924), .Q (signal_19761) ) ;
    buf_clk cell_14879 ( .C (clk), .D (signal_8191), .Q (signal_19767) ) ;
    buf_clk cell_14885 ( .C (clk), .D (signal_5165), .Q (signal_19773) ) ;
    buf_clk cell_14891 ( .C (clk), .D (signal_8442), .Q (signal_19779) ) ;
    buf_clk cell_14897 ( .C (clk), .D (signal_5168), .Q (signal_19785) ) ;
    buf_clk cell_14903 ( .C (clk), .D (signal_8445), .Q (signal_19791) ) ;
    buf_clk cell_14909 ( .C (clk), .D (ciphertext_s0[80]), .Q (signal_19797) ) ;
    buf_clk cell_14915 ( .C (clk), .D (ciphertext_s1[80]), .Q (signal_19803) ) ;
    buf_clk cell_14921 ( .C (clk), .D (signal_4927), .Q (signal_19809) ) ;
    buf_clk cell_14927 ( .C (clk), .D (signal_8194), .Q (signal_19815) ) ;
    buf_clk cell_14933 ( .C (clk), .D (signal_5171), .Q (signal_19821) ) ;
    buf_clk cell_14939 ( .C (clk), .D (signal_8448), .Q (signal_19827) ) ;
    buf_clk cell_14945 ( .C (clk), .D (signal_5173), .Q (signal_19833) ) ;
    buf_clk cell_14951 ( .C (clk), .D (signal_8450), .Q (signal_19839) ) ;
    buf_clk cell_14957 ( .C (clk), .D (signal_4931), .Q (signal_19845) ) ;
    buf_clk cell_14963 ( .C (clk), .D (signal_8198), .Q (signal_19851) ) ;
    buf_clk cell_14969 ( .C (clk), .D (signal_4932), .Q (signal_19857) ) ;
    buf_clk cell_14975 ( .C (clk), .D (signal_8199), .Q (signal_19863) ) ;
    buf_clk cell_14981 ( .C (clk), .D (signal_5172), .Q (signal_19869) ) ;
    buf_clk cell_14987 ( .C (clk), .D (signal_8449), .Q (signal_19875) ) ;
    buf_clk cell_14993 ( .C (clk), .D (signal_4727), .Q (signal_19881) ) ;
    buf_clk cell_14999 ( .C (clk), .D (signal_8081), .Q (signal_19887) ) ;
    buf_clk cell_15005 ( .C (clk), .D (signal_4731), .Q (signal_19893) ) ;
    buf_clk cell_15011 ( .C (clk), .D (signal_8085), .Q (signal_19899) ) ;
    buf_clk cell_15017 ( .C (clk), .D (signal_4730), .Q (signal_19905) ) ;
    buf_clk cell_15023 ( .C (clk), .D (signal_8084), .Q (signal_19911) ) ;
    buf_clk cell_15029 ( .C (clk), .D (signal_4935), .Q (signal_19917) ) ;
    buf_clk cell_15035 ( .C (clk), .D (signal_8279), .Q (signal_19923) ) ;
    buf_clk cell_15041 ( .C (clk), .D (signal_4729), .Q (signal_19929) ) ;
    buf_clk cell_15047 ( .C (clk), .D (signal_8083), .Q (signal_19935) ) ;
    buf_clk cell_15053 ( .C (clk), .D (signal_4561), .Q (signal_19941) ) ;
    buf_clk cell_15059 ( .C (clk), .D (signal_7893), .Q (signal_19947) ) ;
    buf_clk cell_15065 ( .C (clk), .D (signal_4559), .Q (signal_19953) ) ;
    buf_clk cell_15071 ( .C (clk), .D (signal_7891), .Q (signal_19959) ) ;
    buf_clk cell_15077 ( .C (clk), .D (signal_4560), .Q (signal_19965) ) ;
    buf_clk cell_15083 ( .C (clk), .D (signal_7892), .Q (signal_19971) ) ;
    buf_clk cell_15089 ( .C (clk), .D (signal_5181), .Q (signal_19977) ) ;
    buf_clk cell_15095 ( .C (clk), .D (signal_8452), .Q (signal_19983) ) ;
    buf_clk cell_15101 ( .C (clk), .D (ciphertext_s0[96]), .Q (signal_19989) ) ;
    buf_clk cell_15107 ( .C (clk), .D (ciphertext_s1[96]), .Q (signal_19995) ) ;
    buf_clk cell_15113 ( .C (clk), .D (signal_4942), .Q (signal_20001) ) ;
    buf_clk cell_15119 ( .C (clk), .D (signal_8202), .Q (signal_20007) ) ;
    buf_clk cell_15125 ( .C (clk), .D (signal_5184), .Q (signal_20013) ) ;
    buf_clk cell_15131 ( .C (clk), .D (signal_8455), .Q (signal_20019) ) ;
    buf_clk cell_15137 ( .C (clk), .D (signal_5186), .Q (signal_20025) ) ;
    buf_clk cell_15143 ( .C (clk), .D (signal_8457), .Q (signal_20031) ) ;
    buf_clk cell_15149 ( .C (clk), .D (signal_4946), .Q (signal_20037) ) ;
    buf_clk cell_15155 ( .C (clk), .D (signal_8206), .Q (signal_20043) ) ;
    buf_clk cell_15161 ( .C (clk), .D (signal_4947), .Q (signal_20049) ) ;
    buf_clk cell_15167 ( .C (clk), .D (signal_8207), .Q (signal_20055) ) ;
    buf_clk cell_15173 ( .C (clk), .D (signal_5185), .Q (signal_20061) ) ;
    buf_clk cell_15179 ( .C (clk), .D (signal_8456), .Q (signal_20067) ) ;
    buf_clk cell_15185 ( .C (clk), .D (signal_5188), .Q (signal_20073) ) ;
    buf_clk cell_15191 ( .C (clk), .D (signal_8459), .Q (signal_20079) ) ;
    buf_clk cell_15197 ( .C (clk), .D (ciphertext_s0[104]), .Q (signal_20085) ) ;
    buf_clk cell_15203 ( .C (clk), .D (ciphertext_s1[104]), .Q (signal_20091) ) ;
    buf_clk cell_15209 ( .C (clk), .D (signal_4950), .Q (signal_20097) ) ;
    buf_clk cell_15215 ( .C (clk), .D (signal_8210), .Q (signal_20103) ) ;
    buf_clk cell_15221 ( .C (clk), .D (signal_5191), .Q (signal_20109) ) ;
    buf_clk cell_15227 ( .C (clk), .D (signal_8462), .Q (signal_20115) ) ;
    buf_clk cell_15233 ( .C (clk), .D (signal_5193), .Q (signal_20121) ) ;
    buf_clk cell_15239 ( .C (clk), .D (signal_8464), .Q (signal_20127) ) ;
    buf_clk cell_15245 ( .C (clk), .D (signal_4954), .Q (signal_20133) ) ;
    buf_clk cell_15251 ( .C (clk), .D (signal_8214), .Q (signal_20139) ) ;
    buf_clk cell_15257 ( .C (clk), .D (signal_4955), .Q (signal_20145) ) ;
    buf_clk cell_15263 ( .C (clk), .D (signal_8215), .Q (signal_20151) ) ;
    buf_clk cell_15269 ( .C (clk), .D (signal_5192), .Q (signal_20157) ) ;
    buf_clk cell_15275 ( .C (clk), .D (signal_8463), .Q (signal_20163) ) ;
    buf_clk cell_15281 ( .C (clk), .D (signal_5195), .Q (signal_20169) ) ;
    buf_clk cell_15287 ( .C (clk), .D (signal_8466), .Q (signal_20175) ) ;
    buf_clk cell_15293 ( .C (clk), .D (ciphertext_s0[112]), .Q (signal_20181) ) ;
    buf_clk cell_15299 ( .C (clk), .D (ciphertext_s1[112]), .Q (signal_20187) ) ;
    buf_clk cell_15305 ( .C (clk), .D (signal_4958), .Q (signal_20193) ) ;
    buf_clk cell_15311 ( .C (clk), .D (signal_8218), .Q (signal_20199) ) ;
    buf_clk cell_15317 ( .C (clk), .D (signal_5198), .Q (signal_20205) ) ;
    buf_clk cell_15323 ( .C (clk), .D (signal_8469), .Q (signal_20211) ) ;
    buf_clk cell_15329 ( .C (clk), .D (signal_5200), .Q (signal_20217) ) ;
    buf_clk cell_15335 ( .C (clk), .D (signal_8471), .Q (signal_20223) ) ;
    buf_clk cell_15341 ( .C (clk), .D (signal_4962), .Q (signal_20229) ) ;
    buf_clk cell_15347 ( .C (clk), .D (signal_8222), .Q (signal_20235) ) ;
    buf_clk cell_15353 ( .C (clk), .D (signal_4963), .Q (signal_20241) ) ;
    buf_clk cell_15359 ( .C (clk), .D (signal_8223), .Q (signal_20247) ) ;
    buf_clk cell_15365 ( .C (clk), .D (signal_5199), .Q (signal_20253) ) ;
    buf_clk cell_15371 ( .C (clk), .D (signal_8470), .Q (signal_20259) ) ;
    buf_clk cell_15377 ( .C (clk), .D (signal_4765), .Q (signal_20265) ) ;
    buf_clk cell_15383 ( .C (clk), .D (signal_8089), .Q (signal_20271) ) ;
    buf_clk cell_15389 ( .C (clk), .D (signal_4769), .Q (signal_20277) ) ;
    buf_clk cell_15395 ( .C (clk), .D (signal_8093), .Q (signal_20283) ) ;
    buf_clk cell_15401 ( .C (clk), .D (signal_4768), .Q (signal_20289) ) ;
    buf_clk cell_15407 ( .C (clk), .D (signal_8092), .Q (signal_20295) ) ;
    buf_clk cell_15413 ( .C (clk), .D (signal_4966), .Q (signal_20301) ) ;
    buf_clk cell_15419 ( .C (clk), .D (signal_8286), .Q (signal_20307) ) ;
    buf_clk cell_15425 ( .C (clk), .D (signal_4767), .Q (signal_20313) ) ;
    buf_clk cell_15431 ( .C (clk), .D (signal_8091), .Q (signal_20319) ) ;
    buf_clk cell_15437 ( .C (clk), .D (signal_4571), .Q (signal_20325) ) ;
    buf_clk cell_15443 ( .C (clk), .D (signal_7903), .Q (signal_20331) ) ;
    buf_clk cell_15449 ( .C (clk), .D (signal_4569), .Q (signal_20337) ) ;
    buf_clk cell_15455 ( .C (clk), .D (signal_7901), .Q (signal_20343) ) ;
    buf_clk cell_15461 ( .C (clk), .D (signal_4570), .Q (signal_20349) ) ;
    buf_clk cell_15467 ( .C (clk), .D (signal_7902), .Q (signal_20355) ) ;
    buf_clk cell_15473 ( .C (clk), .D (signal_4773), .Q (signal_20361) ) ;
    buf_clk cell_15479 ( .C (clk), .D (signal_8041), .Q (signal_20367) ) ;
    buf_clk cell_15485 ( .C (clk), .D (signal_4777), .Q (signal_20373) ) ;
    buf_clk cell_15491 ( .C (clk), .D (signal_8045), .Q (signal_20379) ) ;
    buf_clk cell_15497 ( .C (clk), .D (signal_4776), .Q (signal_20385) ) ;
    buf_clk cell_15503 ( .C (clk), .D (signal_8044), .Q (signal_20391) ) ;
    buf_clk cell_15509 ( .C (clk), .D (signal_4973), .Q (signal_20397) ) ;
    buf_clk cell_15515 ( .C (clk), .D (signal_8226), .Q (signal_20403) ) ;
    buf_clk cell_15521 ( .C (clk), .D (signal_4775), .Q (signal_20409) ) ;
    buf_clk cell_15527 ( .C (clk), .D (signal_8043), .Q (signal_20415) ) ;
    buf_clk cell_15533 ( .C (clk), .D (signal_4581), .Q (signal_20421) ) ;
    buf_clk cell_15539 ( .C (clk), .D (signal_7843), .Q (signal_20427) ) ;
    buf_clk cell_15545 ( .C (clk), .D (signal_4579), .Q (signal_20433) ) ;
    buf_clk cell_15551 ( .C (clk), .D (signal_7841), .Q (signal_20439) ) ;
    buf_clk cell_15557 ( .C (clk), .D (signal_4580), .Q (signal_20445) ) ;
    buf_clk cell_15563 ( .C (clk), .D (signal_7842), .Q (signal_20451) ) ;
    buf_clk cell_15569 ( .C (clk), .D (signal_4781), .Q (signal_20457) ) ;
    buf_clk cell_15575 ( .C (clk), .D (signal_8049), .Q (signal_20463) ) ;
    buf_clk cell_15581 ( .C (clk), .D (signal_4785), .Q (signal_20469) ) ;
    buf_clk cell_15587 ( .C (clk), .D (signal_8053), .Q (signal_20475) ) ;
    buf_clk cell_15593 ( .C (clk), .D (signal_4784), .Q (signal_20481) ) ;
    buf_clk cell_15599 ( .C (clk), .D (signal_8052), .Q (signal_20487) ) ;
    buf_clk cell_15605 ( .C (clk), .D (signal_4980), .Q (signal_20493) ) ;
    buf_clk cell_15611 ( .C (clk), .D (signal_8233), .Q (signal_20499) ) ;
    buf_clk cell_15617 ( .C (clk), .D (signal_4783), .Q (signal_20505) ) ;
    buf_clk cell_15623 ( .C (clk), .D (signal_8051), .Q (signal_20511) ) ;
    buf_clk cell_15629 ( .C (clk), .D (signal_4591), .Q (signal_20517) ) ;
    buf_clk cell_15635 ( .C (clk), .D (signal_7853), .Q (signal_20523) ) ;
    buf_clk cell_15641 ( .C (clk), .D (signal_4589), .Q (signal_20529) ) ;
    buf_clk cell_15647 ( .C (clk), .D (signal_7851), .Q (signal_20535) ) ;
    buf_clk cell_15653 ( .C (clk), .D (signal_4590), .Q (signal_20541) ) ;
    buf_clk cell_15659 ( .C (clk), .D (signal_7852), .Q (signal_20547) ) ;
    buf_clk cell_15665 ( .C (clk), .D (signal_4789), .Q (signal_20553) ) ;
    buf_clk cell_15671 ( .C (clk), .D (signal_8057), .Q (signal_20559) ) ;
    buf_clk cell_15677 ( .C (clk), .D (signal_4793), .Q (signal_20565) ) ;
    buf_clk cell_15683 ( .C (clk), .D (signal_8061), .Q (signal_20571) ) ;
    buf_clk cell_15689 ( .C (clk), .D (signal_4792), .Q (signal_20577) ) ;
    buf_clk cell_15695 ( .C (clk), .D (signal_8060), .Q (signal_20583) ) ;
    buf_clk cell_15701 ( .C (clk), .D (signal_4987), .Q (signal_20589) ) ;
    buf_clk cell_15707 ( .C (clk), .D (signal_8240), .Q (signal_20595) ) ;
    buf_clk cell_15713 ( .C (clk), .D (signal_4791), .Q (signal_20601) ) ;
    buf_clk cell_15719 ( .C (clk), .D (signal_8059), .Q (signal_20607) ) ;
    buf_clk cell_15725 ( .C (clk), .D (signal_4601), .Q (signal_20613) ) ;
    buf_clk cell_15731 ( .C (clk), .D (signal_7863), .Q (signal_20619) ) ;
    buf_clk cell_15737 ( .C (clk), .D (signal_4599), .Q (signal_20625) ) ;
    buf_clk cell_15743 ( .C (clk), .D (signal_7861), .Q (signal_20631) ) ;
    buf_clk cell_15749 ( .C (clk), .D (signal_4600), .Q (signal_20637) ) ;
    buf_clk cell_15755 ( .C (clk), .D (signal_7862), .Q (signal_20643) ) ;
    buf_clk cell_15761 ( .C (clk), .D (signal_4797), .Q (signal_20649) ) ;
    buf_clk cell_15767 ( .C (clk), .D (signal_8065), .Q (signal_20655) ) ;
    buf_clk cell_15773 ( .C (clk), .D (signal_4801), .Q (signal_20661) ) ;
    buf_clk cell_15779 ( .C (clk), .D (signal_8069), .Q (signal_20667) ) ;
    buf_clk cell_15785 ( .C (clk), .D (signal_4800), .Q (signal_20673) ) ;
    buf_clk cell_15791 ( .C (clk), .D (signal_8068), .Q (signal_20679) ) ;
    buf_clk cell_15797 ( .C (clk), .D (signal_4994), .Q (signal_20685) ) ;
    buf_clk cell_15803 ( .C (clk), .D (signal_8247), .Q (signal_20691) ) ;
    buf_clk cell_15809 ( .C (clk), .D (signal_4799), .Q (signal_20697) ) ;
    buf_clk cell_15815 ( .C (clk), .D (signal_8067), .Q (signal_20703) ) ;
    buf_clk cell_15821 ( .C (clk), .D (signal_4611), .Q (signal_20709) ) ;
    buf_clk cell_15827 ( .C (clk), .D (signal_7873), .Q (signal_20715) ) ;
    buf_clk cell_15833 ( .C (clk), .D (signal_4609), .Q (signal_20721) ) ;
    buf_clk cell_15839 ( .C (clk), .D (signal_7871), .Q (signal_20727) ) ;
    buf_clk cell_15845 ( .C (clk), .D (signal_4610), .Q (signal_20733) ) ;
    buf_clk cell_15851 ( .C (clk), .D (signal_7872), .Q (signal_20739) ) ;
    buf_clk cell_15857 ( .C (clk), .D (signal_4847), .Q (signal_20745) ) ;
    buf_clk cell_15863 ( .C (clk), .D (signal_8121), .Q (signal_20751) ) ;
    buf_clk cell_15869 ( .C (clk), .D (signal_4851), .Q (signal_20757) ) ;
    buf_clk cell_15875 ( .C (clk), .D (signal_8125), .Q (signal_20763) ) ;
    buf_clk cell_15881 ( .C (clk), .D (signal_4850), .Q (signal_20769) ) ;
    buf_clk cell_15887 ( .C (clk), .D (signal_8124), .Q (signal_20775) ) ;
    buf_clk cell_15893 ( .C (clk), .D (signal_5100), .Q (signal_20781) ) ;
    buf_clk cell_15899 ( .C (clk), .D (signal_8383), .Q (signal_20787) ) ;
    buf_clk cell_15905 ( .C (clk), .D (signal_4849), .Q (signal_20793) ) ;
    buf_clk cell_15911 ( .C (clk), .D (signal_8123), .Q (signal_20799) ) ;
    buf_clk cell_15917 ( .C (clk), .D (signal_4621), .Q (signal_20805) ) ;
    buf_clk cell_15923 ( .C (clk), .D (signal_7913), .Q (signal_20811) ) ;
    buf_clk cell_15929 ( .C (clk), .D (signal_4619), .Q (signal_20817) ) ;
    buf_clk cell_15935 ( .C (clk), .D (signal_7911), .Q (signal_20823) ) ;
    buf_clk cell_15941 ( .C (clk), .D (signal_4620), .Q (signal_20829) ) ;
    buf_clk cell_15947 ( .C (clk), .D (signal_7912), .Q (signal_20835) ) ;
    buf_clk cell_15953 ( .C (clk), .D (signal_4855), .Q (signal_20841) ) ;
    buf_clk cell_15959 ( .C (clk), .D (signal_8129), .Q (signal_20847) ) ;
    buf_clk cell_15965 ( .C (clk), .D (signal_4859), .Q (signal_20853) ) ;
    buf_clk cell_15971 ( .C (clk), .D (signal_8133), .Q (signal_20859) ) ;
    buf_clk cell_15977 ( .C (clk), .D (signal_4858), .Q (signal_20865) ) ;
    buf_clk cell_15983 ( .C (clk), .D (signal_8132), .Q (signal_20871) ) ;
    buf_clk cell_15989 ( .C (clk), .D (signal_5107), .Q (signal_20877) ) ;
    buf_clk cell_15995 ( .C (clk), .D (signal_8390), .Q (signal_20883) ) ;
    buf_clk cell_16001 ( .C (clk), .D (signal_4857), .Q (signal_20889) ) ;
    buf_clk cell_16007 ( .C (clk), .D (signal_8131), .Q (signal_20895) ) ;
    buf_clk cell_16013 ( .C (clk), .D (signal_4631), .Q (signal_20901) ) ;
    buf_clk cell_16019 ( .C (clk), .D (signal_7923), .Q (signal_20907) ) ;
    buf_clk cell_16025 ( .C (clk), .D (signal_4629), .Q (signal_20913) ) ;
    buf_clk cell_16031 ( .C (clk), .D (signal_7921), .Q (signal_20919) ) ;
    buf_clk cell_16037 ( .C (clk), .D (signal_4630), .Q (signal_20925) ) ;
    buf_clk cell_16043 ( .C (clk), .D (signal_7922), .Q (signal_20931) ) ;
    buf_clk cell_16049 ( .C (clk), .D (signal_4863), .Q (signal_20937) ) ;
    buf_clk cell_16055 ( .C (clk), .D (signal_8137), .Q (signal_20943) ) ;
    buf_clk cell_16061 ( .C (clk), .D (signal_4867), .Q (signal_20949) ) ;
    buf_clk cell_16067 ( .C (clk), .D (signal_8141), .Q (signal_20955) ) ;
    buf_clk cell_16073 ( .C (clk), .D (signal_4866), .Q (signal_20961) ) ;
    buf_clk cell_16079 ( .C (clk), .D (signal_8140), .Q (signal_20967) ) ;
    buf_clk cell_16085 ( .C (clk), .D (signal_5114), .Q (signal_20973) ) ;
    buf_clk cell_16091 ( .C (clk), .D (signal_8397), .Q (signal_20979) ) ;
    buf_clk cell_16097 ( .C (clk), .D (signal_4865), .Q (signal_20985) ) ;
    buf_clk cell_16103 ( .C (clk), .D (signal_8139), .Q (signal_20991) ) ;
    buf_clk cell_16109 ( .C (clk), .D (signal_4641), .Q (signal_20997) ) ;
    buf_clk cell_16115 ( .C (clk), .D (signal_7933), .Q (signal_21003) ) ;
    buf_clk cell_16121 ( .C (clk), .D (signal_4639), .Q (signal_21009) ) ;
    buf_clk cell_16127 ( .C (clk), .D (signal_7931), .Q (signal_21015) ) ;
    buf_clk cell_16133 ( .C (clk), .D (signal_4640), .Q (signal_21021) ) ;
    buf_clk cell_16139 ( .C (clk), .D (signal_7932), .Q (signal_21027) ) ;
    buf_clk cell_16145 ( .C (clk), .D (signal_4871), .Q (signal_21033) ) ;
    buf_clk cell_16151 ( .C (clk), .D (signal_8145), .Q (signal_21039) ) ;
    buf_clk cell_16157 ( .C (clk), .D (signal_4875), .Q (signal_21045) ) ;
    buf_clk cell_16163 ( .C (clk), .D (signal_8149), .Q (signal_21051) ) ;
    buf_clk cell_16169 ( .C (clk), .D (signal_4874), .Q (signal_21057) ) ;
    buf_clk cell_16175 ( .C (clk), .D (signal_8148), .Q (signal_21063) ) ;
    buf_clk cell_16181 ( .C (clk), .D (signal_5121), .Q (signal_21069) ) ;
    buf_clk cell_16187 ( .C (clk), .D (signal_8404), .Q (signal_21075) ) ;
    buf_clk cell_16193 ( .C (clk), .D (signal_4873), .Q (signal_21081) ) ;
    buf_clk cell_16199 ( .C (clk), .D (signal_8147), .Q (signal_21087) ) ;
    buf_clk cell_16205 ( .C (clk), .D (signal_4651), .Q (signal_21093) ) ;
    buf_clk cell_16211 ( .C (clk), .D (signal_7943), .Q (signal_21099) ) ;
    buf_clk cell_16217 ( .C (clk), .D (signal_4649), .Q (signal_21105) ) ;
    buf_clk cell_16223 ( .C (clk), .D (signal_7941), .Q (signal_21111) ) ;
    buf_clk cell_16229 ( .C (clk), .D (signal_4650), .Q (signal_21117) ) ;
    buf_clk cell_16235 ( .C (clk), .D (signal_7942), .Q (signal_21123) ) ;
    buf_clk cell_16241 ( .C (clk), .D (signal_4879), .Q (signal_21129) ) ;
    buf_clk cell_16247 ( .C (clk), .D (signal_8153), .Q (signal_21135) ) ;
    buf_clk cell_16253 ( .C (clk), .D (signal_4883), .Q (signal_21141) ) ;
    buf_clk cell_16259 ( .C (clk), .D (signal_8157), .Q (signal_21147) ) ;
    buf_clk cell_16265 ( .C (clk), .D (signal_4882), .Q (signal_21153) ) ;
    buf_clk cell_16271 ( .C (clk), .D (signal_8156), .Q (signal_21159) ) ;
    buf_clk cell_16277 ( .C (clk), .D (signal_5128), .Q (signal_21165) ) ;
    buf_clk cell_16283 ( .C (clk), .D (signal_8411), .Q (signal_21171) ) ;
    buf_clk cell_16289 ( .C (clk), .D (signal_4881), .Q (signal_21177) ) ;
    buf_clk cell_16295 ( .C (clk), .D (signal_8155), .Q (signal_21183) ) ;
    buf_clk cell_16301 ( .C (clk), .D (signal_4661), .Q (signal_21189) ) ;
    buf_clk cell_16307 ( .C (clk), .D (signal_7953), .Q (signal_21195) ) ;
    buf_clk cell_16313 ( .C (clk), .D (signal_4659), .Q (signal_21201) ) ;
    buf_clk cell_16319 ( .C (clk), .D (signal_7951), .Q (signal_21207) ) ;
    buf_clk cell_16325 ( .C (clk), .D (signal_4660), .Q (signal_21213) ) ;
    buf_clk cell_16331 ( .C (clk), .D (signal_7952), .Q (signal_21219) ) ;
    buf_clk cell_16337 ( .C (clk), .D (signal_4887), .Q (signal_21225) ) ;
    buf_clk cell_16343 ( .C (clk), .D (signal_8161), .Q (signal_21231) ) ;
    buf_clk cell_16349 ( .C (clk), .D (signal_4891), .Q (signal_21237) ) ;
    buf_clk cell_16355 ( .C (clk), .D (signal_8165), .Q (signal_21243) ) ;
    buf_clk cell_16361 ( .C (clk), .D (signal_4890), .Q (signal_21249) ) ;
    buf_clk cell_16367 ( .C (clk), .D (signal_8164), .Q (signal_21255) ) ;
    buf_clk cell_16373 ( .C (clk), .D (signal_5135), .Q (signal_21261) ) ;
    buf_clk cell_16379 ( .C (clk), .D (signal_8418), .Q (signal_21267) ) ;
    buf_clk cell_16385 ( .C (clk), .D (signal_4889), .Q (signal_21273) ) ;
    buf_clk cell_16391 ( .C (clk), .D (signal_8163), .Q (signal_21279) ) ;
    buf_clk cell_16397 ( .C (clk), .D (signal_4671), .Q (signal_21285) ) ;
    buf_clk cell_16403 ( .C (clk), .D (signal_7963), .Q (signal_21291) ) ;
    buf_clk cell_16409 ( .C (clk), .D (signal_4669), .Q (signal_21297) ) ;
    buf_clk cell_16415 ( .C (clk), .D (signal_7961), .Q (signal_21303) ) ;
    buf_clk cell_16421 ( .C (clk), .D (signal_4670), .Q (signal_21309) ) ;
    buf_clk cell_16427 ( .C (clk), .D (signal_7962), .Q (signal_21315) ) ;
    buf_clk cell_16433 ( .C (clk), .D (signal_4895), .Q (signal_21321) ) ;
    buf_clk cell_16439 ( .C (clk), .D (signal_8169), .Q (signal_21327) ) ;
    buf_clk cell_16445 ( .C (clk), .D (signal_4899), .Q (signal_21333) ) ;
    buf_clk cell_16451 ( .C (clk), .D (signal_8173), .Q (signal_21339) ) ;
    buf_clk cell_16457 ( .C (clk), .D (signal_4898), .Q (signal_21345) ) ;
    buf_clk cell_16463 ( .C (clk), .D (signal_8172), .Q (signal_21351) ) ;
    buf_clk cell_16469 ( .C (clk), .D (signal_5142), .Q (signal_21357) ) ;
    buf_clk cell_16475 ( .C (clk), .D (signal_8425), .Q (signal_21363) ) ;
    buf_clk cell_16481 ( .C (clk), .D (signal_4897), .Q (signal_21369) ) ;
    buf_clk cell_16487 ( .C (clk), .D (signal_8171), .Q (signal_21375) ) ;
    buf_clk cell_16493 ( .C (clk), .D (signal_4681), .Q (signal_21381) ) ;
    buf_clk cell_16499 ( .C (clk), .D (signal_7973), .Q (signal_21387) ) ;
    buf_clk cell_16505 ( .C (clk), .D (signal_4679), .Q (signal_21393) ) ;
    buf_clk cell_16511 ( .C (clk), .D (signal_7971), .Q (signal_21399) ) ;
    buf_clk cell_16517 ( .C (clk), .D (signal_4680), .Q (signal_21405) ) ;
    buf_clk cell_16523 ( .C (clk), .D (signal_7972), .Q (signal_21411) ) ;
    buf_clk cell_16529 ( .C (clk), .D (signal_4696), .Q (signal_21417) ) ;
    buf_clk cell_16535 ( .C (clk), .D (signal_8080), .Q (signal_21423) ) ;
    buf_clk cell_16541 ( .C (clk), .D (signal_4552), .Q (signal_21429) ) ;
    buf_clk cell_16547 ( .C (clk), .D (signal_7884), .Q (signal_21435) ) ;
    buf_clk cell_16553 ( .C (clk), .D (signal_4910), .Q (signal_21441) ) ;
    buf_clk cell_16559 ( .C (clk), .D (signal_8177), .Q (signal_21447) ) ;
    buf_clk cell_16565 ( .C (clk), .D (signal_4914), .Q (signal_21453) ) ;
    buf_clk cell_16571 ( .C (clk), .D (signal_8181), .Q (signal_21459) ) ;
    buf_clk cell_16577 ( .C (clk), .D (signal_4913), .Q (signal_21465) ) ;
    buf_clk cell_16583 ( .C (clk), .D (signal_8180), .Q (signal_21471) ) ;
    buf_clk cell_16589 ( .C (clk), .D (signal_5155), .Q (signal_21477) ) ;
    buf_clk cell_16595 ( .C (clk), .D (signal_8432), .Q (signal_21483) ) ;
    buf_clk cell_16601 ( .C (clk), .D (signal_4912), .Q (signal_21489) ) ;
    buf_clk cell_16607 ( .C (clk), .D (signal_8179), .Q (signal_21495) ) ;
    buf_clk cell_16613 ( .C (clk), .D (signal_4699), .Q (signal_21501) ) ;
    buf_clk cell_16619 ( .C (clk), .D (signal_7983), .Q (signal_21507) ) ;
    buf_clk cell_16625 ( .C (clk), .D (signal_4697), .Q (signal_21513) ) ;
    buf_clk cell_16631 ( .C (clk), .D (signal_7981), .Q (signal_21519) ) ;
    buf_clk cell_16637 ( .C (clk), .D (signal_4698), .Q (signal_21525) ) ;
    buf_clk cell_16643 ( .C (clk), .D (signal_7982), .Q (signal_21531) ) ;
    buf_clk cell_16649 ( .C (clk), .D (signal_4918), .Q (signal_21537) ) ;
    buf_clk cell_16655 ( .C (clk), .D (signal_8185), .Q (signal_21543) ) ;
    buf_clk cell_16661 ( .C (clk), .D (signal_4922), .Q (signal_21549) ) ;
    buf_clk cell_16667 ( .C (clk), .D (signal_8189), .Q (signal_21555) ) ;
    buf_clk cell_16673 ( .C (clk), .D (signal_4921), .Q (signal_21561) ) ;
    buf_clk cell_16679 ( .C (clk), .D (signal_8188), .Q (signal_21567) ) ;
    buf_clk cell_16685 ( .C (clk), .D (signal_5162), .Q (signal_21573) ) ;
    buf_clk cell_16691 ( .C (clk), .D (signal_8439), .Q (signal_21579) ) ;
    buf_clk cell_16697 ( .C (clk), .D (signal_4920), .Q (signal_21585) ) ;
    buf_clk cell_16703 ( .C (clk), .D (signal_8187), .Q (signal_21591) ) ;
    buf_clk cell_16709 ( .C (clk), .D (signal_4709), .Q (signal_21597) ) ;
    buf_clk cell_16715 ( .C (clk), .D (signal_7993), .Q (signal_21603) ) ;
    buf_clk cell_16721 ( .C (clk), .D (signal_4707), .Q (signal_21609) ) ;
    buf_clk cell_16727 ( .C (clk), .D (signal_7991), .Q (signal_21615) ) ;
    buf_clk cell_16733 ( .C (clk), .D (signal_4708), .Q (signal_21621) ) ;
    buf_clk cell_16739 ( .C (clk), .D (signal_7992), .Q (signal_21627) ) ;
    buf_clk cell_16745 ( .C (clk), .D (signal_4926), .Q (signal_21633) ) ;
    buf_clk cell_16751 ( .C (clk), .D (signal_8193), .Q (signal_21639) ) ;
    buf_clk cell_16757 ( .C (clk), .D (signal_4930), .Q (signal_21645) ) ;
    buf_clk cell_16763 ( .C (clk), .D (signal_8197), .Q (signal_21651) ) ;
    buf_clk cell_16769 ( .C (clk), .D (signal_4929), .Q (signal_21657) ) ;
    buf_clk cell_16775 ( .C (clk), .D (signal_8196), .Q (signal_21663) ) ;
    buf_clk cell_16781 ( .C (clk), .D (signal_5169), .Q (signal_21669) ) ;
    buf_clk cell_16787 ( .C (clk), .D (signal_8446), .Q (signal_21675) ) ;
    buf_clk cell_16793 ( .C (clk), .D (signal_4928), .Q (signal_21681) ) ;
    buf_clk cell_16799 ( .C (clk), .D (signal_8195), .Q (signal_21687) ) ;
    buf_clk cell_16805 ( .C (clk), .D (signal_4719), .Q (signal_21693) ) ;
    buf_clk cell_16811 ( .C (clk), .D (signal_8003), .Q (signal_21699) ) ;
    buf_clk cell_16817 ( .C (clk), .D (signal_4717), .Q (signal_21705) ) ;
    buf_clk cell_16823 ( .C (clk), .D (signal_8001), .Q (signal_21711) ) ;
    buf_clk cell_16829 ( .C (clk), .D (signal_4718), .Q (signal_21717) ) ;
    buf_clk cell_16835 ( .C (clk), .D (signal_8002), .Q (signal_21723) ) ;
    buf_clk cell_16841 ( .C (clk), .D (signal_4734), .Q (signal_21729) ) ;
    buf_clk cell_16847 ( .C (clk), .D (signal_8088), .Q (signal_21735) ) ;
    buf_clk cell_16853 ( .C (clk), .D (signal_4562), .Q (signal_21741) ) ;
    buf_clk cell_16859 ( .C (clk), .D (signal_7894), .Q (signal_21747) ) ;
    buf_clk cell_16865 ( .C (clk), .D (signal_4941), .Q (signal_21753) ) ;
    buf_clk cell_16871 ( .C (clk), .D (signal_8201), .Q (signal_21759) ) ;
    buf_clk cell_16877 ( .C (clk), .D (signal_4945), .Q (signal_21765) ) ;
    buf_clk cell_16883 ( .C (clk), .D (signal_8205), .Q (signal_21771) ) ;
    buf_clk cell_16889 ( .C (clk), .D (signal_4944), .Q (signal_21777) ) ;
    buf_clk cell_16895 ( .C (clk), .D (signal_8204), .Q (signal_21783) ) ;
    buf_clk cell_16901 ( .C (clk), .D (signal_5182), .Q (signal_21789) ) ;
    buf_clk cell_16907 ( .C (clk), .D (signal_8453), .Q (signal_21795) ) ;
    buf_clk cell_16913 ( .C (clk), .D (signal_4943), .Q (signal_21801) ) ;
    buf_clk cell_16919 ( .C (clk), .D (signal_8203), .Q (signal_21807) ) ;
    buf_clk cell_16925 ( .C (clk), .D (signal_4737), .Q (signal_21813) ) ;
    buf_clk cell_16931 ( .C (clk), .D (signal_8013), .Q (signal_21819) ) ;
    buf_clk cell_16937 ( .C (clk), .D (signal_4735), .Q (signal_21825) ) ;
    buf_clk cell_16943 ( .C (clk), .D (signal_8011), .Q (signal_21831) ) ;
    buf_clk cell_16949 ( .C (clk), .D (signal_4736), .Q (signal_21837) ) ;
    buf_clk cell_16955 ( .C (clk), .D (signal_8012), .Q (signal_21843) ) ;
    buf_clk cell_16961 ( .C (clk), .D (signal_4949), .Q (signal_21849) ) ;
    buf_clk cell_16967 ( .C (clk), .D (signal_8209), .Q (signal_21855) ) ;
    buf_clk cell_16973 ( .C (clk), .D (signal_4953), .Q (signal_21861) ) ;
    buf_clk cell_16979 ( .C (clk), .D (signal_8213), .Q (signal_21867) ) ;
    buf_clk cell_16985 ( .C (clk), .D (signal_4952), .Q (signal_21873) ) ;
    buf_clk cell_16991 ( .C (clk), .D (signal_8212), .Q (signal_21879) ) ;
    buf_clk cell_16997 ( .C (clk), .D (signal_5189), .Q (signal_21885) ) ;
    buf_clk cell_17003 ( .C (clk), .D (signal_8460), .Q (signal_21891) ) ;
    buf_clk cell_17009 ( .C (clk), .D (signal_4951), .Q (signal_21897) ) ;
    buf_clk cell_17015 ( .C (clk), .D (signal_8211), .Q (signal_21903) ) ;
    buf_clk cell_17021 ( .C (clk), .D (signal_4747), .Q (signal_21909) ) ;
    buf_clk cell_17027 ( .C (clk), .D (signal_8023), .Q (signal_21915) ) ;
    buf_clk cell_17033 ( .C (clk), .D (signal_4745), .Q (signal_21921) ) ;
    buf_clk cell_17039 ( .C (clk), .D (signal_8021), .Q (signal_21927) ) ;
    buf_clk cell_17045 ( .C (clk), .D (signal_4746), .Q (signal_21933) ) ;
    buf_clk cell_17051 ( .C (clk), .D (signal_8022), .Q (signal_21939) ) ;
    buf_clk cell_17057 ( .C (clk), .D (signal_4957), .Q (signal_21945) ) ;
    buf_clk cell_17063 ( .C (clk), .D (signal_8217), .Q (signal_21951) ) ;
    buf_clk cell_17069 ( .C (clk), .D (signal_4961), .Q (signal_21957) ) ;
    buf_clk cell_17075 ( .C (clk), .D (signal_8221), .Q (signal_21963) ) ;
    buf_clk cell_17081 ( .C (clk), .D (signal_4960), .Q (signal_21969) ) ;
    buf_clk cell_17087 ( .C (clk), .D (signal_8220), .Q (signal_21975) ) ;
    buf_clk cell_17093 ( .C (clk), .D (signal_5196), .Q (signal_21981) ) ;
    buf_clk cell_17099 ( .C (clk), .D (signal_8467), .Q (signal_21987) ) ;
    buf_clk cell_17105 ( .C (clk), .D (signal_4959), .Q (signal_21993) ) ;
    buf_clk cell_17111 ( .C (clk), .D (signal_8219), .Q (signal_21999) ) ;
    buf_clk cell_17117 ( .C (clk), .D (signal_4757), .Q (signal_22005) ) ;
    buf_clk cell_17123 ( .C (clk), .D (signal_8033), .Q (signal_22011) ) ;
    buf_clk cell_17129 ( .C (clk), .D (signal_4755), .Q (signal_22017) ) ;
    buf_clk cell_17135 ( .C (clk), .D (signal_8031), .Q (signal_22023) ) ;
    buf_clk cell_17141 ( .C (clk), .D (signal_4756), .Q (signal_22029) ) ;
    buf_clk cell_17147 ( .C (clk), .D (signal_8032), .Q (signal_22035) ) ;
    buf_clk cell_17153 ( .C (clk), .D (signal_4772), .Q (signal_22041) ) ;
    buf_clk cell_17159 ( .C (clk), .D (signal_8096), .Q (signal_22047) ) ;
    buf_clk cell_17165 ( .C (clk), .D (signal_4572), .Q (signal_22053) ) ;
    buf_clk cell_17171 ( .C (clk), .D (signal_7904), .Q (signal_22059) ) ;
    buf_clk cell_17177 ( .C (clk), .D (signal_4780), .Q (signal_22065) ) ;
    buf_clk cell_17183 ( .C (clk), .D (signal_8048), .Q (signal_22071) ) ;
    buf_clk cell_17189 ( .C (clk), .D (signal_4582), .Q (signal_22077) ) ;
    buf_clk cell_17195 ( .C (clk), .D (signal_7844), .Q (signal_22083) ) ;
    buf_clk cell_17201 ( .C (clk), .D (signal_4788), .Q (signal_22089) ) ;
    buf_clk cell_17207 ( .C (clk), .D (signal_8056), .Q (signal_22095) ) ;
    buf_clk cell_17213 ( .C (clk), .D (signal_4592), .Q (signal_22101) ) ;
    buf_clk cell_17219 ( .C (clk), .D (signal_7854), .Q (signal_22107) ) ;
    buf_clk cell_17225 ( .C (clk), .D (signal_4796), .Q (signal_22113) ) ;
    buf_clk cell_17231 ( .C (clk), .D (signal_8064), .Q (signal_22119) ) ;
    buf_clk cell_17237 ( .C (clk), .D (signal_4602), .Q (signal_22125) ) ;
    buf_clk cell_17243 ( .C (clk), .D (signal_7864), .Q (signal_22131) ) ;
    buf_clk cell_17249 ( .C (clk), .D (signal_4804), .Q (signal_22137) ) ;
    buf_clk cell_17255 ( .C (clk), .D (signal_8072), .Q (signal_22143) ) ;
    buf_clk cell_17261 ( .C (clk), .D (signal_4612), .Q (signal_22149) ) ;
    buf_clk cell_17267 ( .C (clk), .D (signal_7874), .Q (signal_22155) ) ;
    buf_clk cell_17273 ( .C (clk), .D (signal_4854), .Q (signal_22161) ) ;
    buf_clk cell_17279 ( .C (clk), .D (signal_8128), .Q (signal_22167) ) ;
    buf_clk cell_17285 ( .C (clk), .D (signal_4622), .Q (signal_22173) ) ;
    buf_clk cell_17291 ( .C (clk), .D (signal_7914), .Q (signal_22179) ) ;
    buf_clk cell_17297 ( .C (clk), .D (signal_4862), .Q (signal_22185) ) ;
    buf_clk cell_17303 ( .C (clk), .D (signal_8136), .Q (signal_22191) ) ;
    buf_clk cell_17309 ( .C (clk), .D (signal_4632), .Q (signal_22197) ) ;
    buf_clk cell_17315 ( .C (clk), .D (signal_7924), .Q (signal_22203) ) ;
    buf_clk cell_17321 ( .C (clk), .D (signal_4870), .Q (signal_22209) ) ;
    buf_clk cell_17327 ( .C (clk), .D (signal_8144), .Q (signal_22215) ) ;
    buf_clk cell_17333 ( .C (clk), .D (signal_4642), .Q (signal_22221) ) ;
    buf_clk cell_17339 ( .C (clk), .D (signal_7934), .Q (signal_22227) ) ;
    buf_clk cell_17345 ( .C (clk), .D (signal_4878), .Q (signal_22233) ) ;
    buf_clk cell_17351 ( .C (clk), .D (signal_8152), .Q (signal_22239) ) ;
    buf_clk cell_17357 ( .C (clk), .D (signal_4652), .Q (signal_22245) ) ;
    buf_clk cell_17363 ( .C (clk), .D (signal_7944), .Q (signal_22251) ) ;
    buf_clk cell_17369 ( .C (clk), .D (signal_4886), .Q (signal_22257) ) ;
    buf_clk cell_17375 ( .C (clk), .D (signal_8160), .Q (signal_22263) ) ;
    buf_clk cell_17381 ( .C (clk), .D (signal_4662), .Q (signal_22269) ) ;
    buf_clk cell_17387 ( .C (clk), .D (signal_7954), .Q (signal_22275) ) ;
    buf_clk cell_17393 ( .C (clk), .D (signal_4894), .Q (signal_22281) ) ;
    buf_clk cell_17399 ( .C (clk), .D (signal_8168), .Q (signal_22287) ) ;
    buf_clk cell_17405 ( .C (clk), .D (signal_4672), .Q (signal_22293) ) ;
    buf_clk cell_17411 ( .C (clk), .D (signal_7964), .Q (signal_22299) ) ;
    buf_clk cell_17417 ( .C (clk), .D (signal_4902), .Q (signal_22305) ) ;
    buf_clk cell_17423 ( .C (clk), .D (signal_8176), .Q (signal_22311) ) ;
    buf_clk cell_17429 ( .C (clk), .D (signal_4682), .Q (signal_22317) ) ;
    buf_clk cell_17435 ( .C (clk), .D (signal_7974), .Q (signal_22323) ) ;
    buf_clk cell_17441 ( .C (clk), .D (signal_4917), .Q (signal_22329) ) ;
    buf_clk cell_17447 ( .C (clk), .D (signal_8184), .Q (signal_22335) ) ;
    buf_clk cell_17453 ( .C (clk), .D (signal_4700), .Q (signal_22341) ) ;
    buf_clk cell_17459 ( .C (clk), .D (signal_7984), .Q (signal_22347) ) ;
    buf_clk cell_17465 ( .C (clk), .D (signal_4925), .Q (signal_22353) ) ;
    buf_clk cell_17471 ( .C (clk), .D (signal_8192), .Q (signal_22359) ) ;
    buf_clk cell_17477 ( .C (clk), .D (signal_4710), .Q (signal_22365) ) ;
    buf_clk cell_17483 ( .C (clk), .D (signal_7994), .Q (signal_22371) ) ;
    buf_clk cell_17489 ( .C (clk), .D (signal_4933), .Q (signal_22377) ) ;
    buf_clk cell_17495 ( .C (clk), .D (signal_8200), .Q (signal_22383) ) ;
    buf_clk cell_17501 ( .C (clk), .D (signal_4720), .Q (signal_22389) ) ;
    buf_clk cell_17507 ( .C (clk), .D (signal_8004), .Q (signal_22395) ) ;
    buf_clk cell_17513 ( .C (clk), .D (signal_4948), .Q (signal_22401) ) ;
    buf_clk cell_17519 ( .C (clk), .D (signal_8208), .Q (signal_22407) ) ;
    buf_clk cell_17525 ( .C (clk), .D (signal_4738), .Q (signal_22413) ) ;
    buf_clk cell_17531 ( .C (clk), .D (signal_8014), .Q (signal_22419) ) ;
    buf_clk cell_17537 ( .C (clk), .D (signal_4956), .Q (signal_22425) ) ;
    buf_clk cell_17543 ( .C (clk), .D (signal_8216), .Q (signal_22431) ) ;
    buf_clk cell_17549 ( .C (clk), .D (signal_4748), .Q (signal_22437) ) ;
    buf_clk cell_17555 ( .C (clk), .D (signal_8024), .Q (signal_22443) ) ;
    buf_clk cell_17561 ( .C (clk), .D (signal_4964), .Q (signal_22449) ) ;
    buf_clk cell_17567 ( .C (clk), .D (signal_8224), .Q (signal_22455) ) ;
    buf_clk cell_17573 ( .C (clk), .D (signal_4758), .Q (signal_22461) ) ;
    buf_clk cell_17579 ( .C (clk), .D (signal_8034), .Q (signal_22467) ) ;
    buf_clk cell_17585 ( .C (clk), .D (signal_4266), .Q (signal_22473) ) ;
    buf_clk cell_17593 ( .C (clk), .D (signal_7571), .Q (signal_22481) ) ;
    buf_clk cell_17601 ( .C (clk), .D (signal_4274), .Q (signal_22489) ) ;
    buf_clk cell_17609 ( .C (clk), .D (signal_7544), .Q (signal_22497) ) ;
    buf_clk cell_17617 ( .C (clk), .D (signal_4282), .Q (signal_22505) ) ;
    buf_clk cell_17625 ( .C (clk), .D (signal_7826), .Q (signal_22513) ) ;
    buf_clk cell_17633 ( .C (clk), .D (signal_4306), .Q (signal_22521) ) ;
    buf_clk cell_17641 ( .C (clk), .D (signal_7772), .Q (signal_22529) ) ;
    buf_clk cell_17649 ( .C (clk), .D (signal_4279), .Q (signal_22537) ) ;
    buf_clk cell_17657 ( .C (clk), .D (signal_7835), .Q (signal_22545) ) ;
    buf_clk cell_17665 ( .C (clk), .D (signal_4280), .Q (signal_22553) ) ;
    buf_clk cell_17673 ( .C (clk), .D (signal_7832), .Q (signal_22561) ) ;
    buf_clk cell_17681 ( .C (clk), .D (signal_4281), .Q (signal_22569) ) ;
    buf_clk cell_17689 ( .C (clk), .D (signal_7829), .Q (signal_22577) ) ;
    buf_clk cell_17697 ( .C (clk), .D (signal_4298), .Q (signal_22585) ) ;
    buf_clk cell_17705 ( .C (clk), .D (signal_7799), .Q (signal_22593) ) ;
    buf_clk cell_17713 ( .C (clk), .D (signal_4259), .Q (signal_22601) ) ;
    buf_clk cell_17721 ( .C (clk), .D (signal_7592), .Q (signal_22609) ) ;
    buf_clk cell_17729 ( .C (clk), .D (signal_4260), .Q (signal_22617) ) ;
    buf_clk cell_17737 ( .C (clk), .D (signal_7589), .Q (signal_22625) ) ;
    buf_clk cell_17745 ( .C (clk), .D (signal_4261), .Q (signal_22633) ) ;
    buf_clk cell_17753 ( .C (clk), .D (signal_7586), .Q (signal_22641) ) ;
    buf_clk cell_17761 ( .C (clk), .D (signal_4262), .Q (signal_22649) ) ;
    buf_clk cell_17769 ( .C (clk), .D (signal_7583), .Q (signal_22657) ) ;
    buf_clk cell_17777 ( .C (clk), .D (signal_4263), .Q (signal_22665) ) ;
    buf_clk cell_17785 ( .C (clk), .D (signal_7580), .Q (signal_22673) ) ;
    buf_clk cell_17793 ( .C (clk), .D (signal_4264), .Q (signal_22681) ) ;
    buf_clk cell_17801 ( .C (clk), .D (signal_7577), .Q (signal_22689) ) ;
    buf_clk cell_17809 ( .C (clk), .D (signal_4265), .Q (signal_22697) ) ;
    buf_clk cell_17817 ( .C (clk), .D (signal_7574), .Q (signal_22705) ) ;
    buf_clk cell_17825 ( .C (clk), .D (signal_4267), .Q (signal_22713) ) ;
    buf_clk cell_17833 ( .C (clk), .D (signal_7568), .Q (signal_22721) ) ;
    buf_clk cell_17841 ( .C (clk), .D (signal_4268), .Q (signal_22729) ) ;
    buf_clk cell_17849 ( .C (clk), .D (signal_7565), .Q (signal_22737) ) ;
    buf_clk cell_17857 ( .C (clk), .D (signal_4269), .Q (signal_22745) ) ;
    buf_clk cell_17865 ( .C (clk), .D (signal_7559), .Q (signal_22753) ) ;
    buf_clk cell_17873 ( .C (clk), .D (signal_4270), .Q (signal_22761) ) ;
    buf_clk cell_17881 ( .C (clk), .D (signal_7556), .Q (signal_22769) ) ;
    buf_clk cell_17889 ( .C (clk), .D (signal_4271), .Q (signal_22777) ) ;
    buf_clk cell_17897 ( .C (clk), .D (signal_7553), .Q (signal_22785) ) ;
    buf_clk cell_17905 ( .C (clk), .D (signal_4272), .Q (signal_22793) ) ;
    buf_clk cell_17913 ( .C (clk), .D (signal_7550), .Q (signal_22801) ) ;
    buf_clk cell_17921 ( .C (clk), .D (signal_4273), .Q (signal_22809) ) ;
    buf_clk cell_17929 ( .C (clk), .D (signal_7547), .Q (signal_22817) ) ;
    buf_clk cell_17937 ( .C (clk), .D (signal_4275), .Q (signal_22825) ) ;
    buf_clk cell_17945 ( .C (clk), .D (signal_7541), .Q (signal_22833) ) ;
    buf_clk cell_17953 ( .C (clk), .D (signal_4276), .Q (signal_22841) ) ;
    buf_clk cell_17961 ( .C (clk), .D (signal_7538), .Q (signal_22849) ) ;
    buf_clk cell_17969 ( .C (clk), .D (signal_4277), .Q (signal_22857) ) ;
    buf_clk cell_17977 ( .C (clk), .D (signal_7535), .Q (signal_22865) ) ;
    buf_clk cell_17985 ( .C (clk), .D (signal_4278), .Q (signal_22873) ) ;
    buf_clk cell_17993 ( .C (clk), .D (signal_7532), .Q (signal_22881) ) ;
    buf_clk cell_18001 ( .C (clk), .D (signal_4314), .Q (signal_22889) ) ;
    buf_clk cell_18009 ( .C (clk), .D (signal_7745), .Q (signal_22897) ) ;
    buf_clk cell_18017 ( .C (clk), .D (signal_4305), .Q (signal_22905) ) ;
    buf_clk cell_18025 ( .C (clk), .D (signal_7775), .Q (signal_22913) ) ;
    buf_clk cell_18033 ( .C (clk), .D (signal_4338), .Q (signal_22921) ) ;
    buf_clk cell_18041 ( .C (clk), .D (signal_7691), .Q (signal_22929) ) ;
    buf_clk cell_18049 ( .C (clk), .D (signal_4307), .Q (signal_22937) ) ;
    buf_clk cell_18057 ( .C (clk), .D (signal_7769), .Q (signal_22945) ) ;
    buf_clk cell_18065 ( .C (clk), .D (signal_4308), .Q (signal_22953) ) ;
    buf_clk cell_18073 ( .C (clk), .D (signal_7766), .Q (signal_22961) ) ;
    buf_clk cell_18081 ( .C (clk), .D (signal_4309), .Q (signal_22969) ) ;
    buf_clk cell_18089 ( .C (clk), .D (signal_7760), .Q (signal_22977) ) ;
    buf_clk cell_18097 ( .C (clk), .D (signal_4310), .Q (signal_22985) ) ;
    buf_clk cell_18105 ( .C (clk), .D (signal_7757), .Q (signal_22993) ) ;
    buf_clk cell_18113 ( .C (clk), .D (signal_4311), .Q (signal_23001) ) ;
    buf_clk cell_18121 ( .C (clk), .D (signal_7754), .Q (signal_23009) ) ;
    buf_clk cell_18129 ( .C (clk), .D (signal_4312), .Q (signal_23017) ) ;
    buf_clk cell_18137 ( .C (clk), .D (signal_7751), .Q (signal_23025) ) ;
    buf_clk cell_18145 ( .C (clk), .D (signal_4291), .Q (signal_23033) ) ;
    buf_clk cell_18153 ( .C (clk), .D (signal_7820), .Q (signal_23041) ) ;
    buf_clk cell_18161 ( .C (clk), .D (signal_4292), .Q (signal_23049) ) ;
    buf_clk cell_18169 ( .C (clk), .D (signal_7817), .Q (signal_23057) ) ;
    buf_clk cell_18177 ( .C (clk), .D (signal_4293), .Q (signal_23065) ) ;
    buf_clk cell_18185 ( .C (clk), .D (signal_7814), .Q (signal_23073) ) ;
    buf_clk cell_18193 ( .C (clk), .D (signal_4294), .Q (signal_23081) ) ;
    buf_clk cell_18201 ( .C (clk), .D (signal_7811), .Q (signal_23089) ) ;
    buf_clk cell_18209 ( .C (clk), .D (signal_4313), .Q (signal_23097) ) ;
    buf_clk cell_18217 ( .C (clk), .D (signal_7748), .Q (signal_23105) ) ;
    buf_clk cell_18225 ( .C (clk), .D (signal_4295), .Q (signal_23113) ) ;
    buf_clk cell_18233 ( .C (clk), .D (signal_7808), .Q (signal_23121) ) ;
    buf_clk cell_18241 ( .C (clk), .D (signal_4296), .Q (signal_23129) ) ;
    buf_clk cell_18249 ( .C (clk), .D (signal_7805), .Q (signal_23137) ) ;
    buf_clk cell_18257 ( .C (clk), .D (signal_4297), .Q (signal_23145) ) ;
    buf_clk cell_18265 ( .C (clk), .D (signal_7802), .Q (signal_23153) ) ;
    buf_clk cell_18273 ( .C (clk), .D (signal_4330), .Q (signal_23161) ) ;
    buf_clk cell_18281 ( .C (clk), .D (signal_7715), .Q (signal_23169) ) ;
    buf_clk cell_18289 ( .C (clk), .D (signal_4299), .Q (signal_23177) ) ;
    buf_clk cell_18297 ( .C (clk), .D (signal_7793), .Q (signal_23185) ) ;
    buf_clk cell_18305 ( .C (clk), .D (signal_4300), .Q (signal_23193) ) ;
    buf_clk cell_18313 ( .C (clk), .D (signal_7790), .Q (signal_23201) ) ;
    buf_clk cell_18321 ( .C (clk), .D (signal_4301), .Q (signal_23209) ) ;
    buf_clk cell_18329 ( .C (clk), .D (signal_7787), .Q (signal_23217) ) ;
    buf_clk cell_18337 ( .C (clk), .D (signal_4302), .Q (signal_23225) ) ;
    buf_clk cell_18345 ( .C (clk), .D (signal_7784), .Q (signal_23233) ) ;
    buf_clk cell_18353 ( .C (clk), .D (signal_4303), .Q (signal_23241) ) ;
    buf_clk cell_18361 ( .C (clk), .D (signal_7781), .Q (signal_23249) ) ;
    buf_clk cell_18369 ( .C (clk), .D (signal_4304), .Q (signal_23257) ) ;
    buf_clk cell_18377 ( .C (clk), .D (signal_7778), .Q (signal_23265) ) ;
    buf_clk cell_18385 ( .C (clk), .D (signal_4346), .Q (signal_23273) ) ;
    buf_clk cell_18393 ( .C (clk), .D (signal_7664), .Q (signal_23281) ) ;
    buf_clk cell_18405 ( .C (clk), .D (signal_4337), .Q (signal_23293) ) ;
    buf_clk cell_18413 ( .C (clk), .D (signal_7694), .Q (signal_23301) ) ;
    buf_clk cell_18421 ( .C (clk), .D (signal_4339), .Q (signal_23309) ) ;
    buf_clk cell_18429 ( .C (clk), .D (signal_7685), .Q (signal_23317) ) ;
    buf_clk cell_18437 ( .C (clk), .D (signal_4340), .Q (signal_23325) ) ;
    buf_clk cell_18445 ( .C (clk), .D (signal_7682), .Q (signal_23333) ) ;
    buf_clk cell_18453 ( .C (clk), .D (signal_4341), .Q (signal_23341) ) ;
    buf_clk cell_18461 ( .C (clk), .D (signal_7679), .Q (signal_23349) ) ;
    buf_clk cell_18469 ( .C (clk), .D (signal_4342), .Q (signal_23357) ) ;
    buf_clk cell_18477 ( .C (clk), .D (signal_7676), .Q (signal_23365) ) ;
    buf_clk cell_18485 ( .C (clk), .D (signal_4343), .Q (signal_23373) ) ;
    buf_clk cell_18493 ( .C (clk), .D (signal_7673), .Q (signal_23381) ) ;
    buf_clk cell_18501 ( .C (clk), .D (signal_4344), .Q (signal_23389) ) ;
    buf_clk cell_18509 ( .C (clk), .D (signal_7670), .Q (signal_23397) ) ;
    buf_clk cell_18517 ( .C (clk), .D (signal_4323), .Q (signal_23405) ) ;
    buf_clk cell_18525 ( .C (clk), .D (signal_7739), .Q (signal_23413) ) ;
    buf_clk cell_18533 ( .C (clk), .D (signal_4324), .Q (signal_23421) ) ;
    buf_clk cell_18541 ( .C (clk), .D (signal_7736), .Q (signal_23429) ) ;
    buf_clk cell_18549 ( .C (clk), .D (signal_4325), .Q (signal_23437) ) ;
    buf_clk cell_18557 ( .C (clk), .D (signal_7733), .Q (signal_23445) ) ;
    buf_clk cell_18565 ( .C (clk), .D (signal_4326), .Q (signal_23453) ) ;
    buf_clk cell_18573 ( .C (clk), .D (signal_7730), .Q (signal_23461) ) ;
    buf_clk cell_18581 ( .C (clk), .D (signal_4345), .Q (signal_23469) ) ;
    buf_clk cell_18589 ( .C (clk), .D (signal_7667), .Q (signal_23477) ) ;
    buf_clk cell_18597 ( .C (clk), .D (signal_4327), .Q (signal_23485) ) ;
    buf_clk cell_18605 ( .C (clk), .D (signal_7727), .Q (signal_23493) ) ;
    buf_clk cell_18613 ( .C (clk), .D (signal_4328), .Q (signal_23501) ) ;
    buf_clk cell_18621 ( .C (clk), .D (signal_7724), .Q (signal_23509) ) ;
    buf_clk cell_18629 ( .C (clk), .D (signal_4329), .Q (signal_23517) ) ;
    buf_clk cell_18637 ( .C (clk), .D (signal_7718), .Q (signal_23525) ) ;
    buf_clk cell_18649 ( .C (clk), .D (signal_4331), .Q (signal_23537) ) ;
    buf_clk cell_18657 ( .C (clk), .D (signal_7712), .Q (signal_23545) ) ;
    buf_clk cell_18665 ( .C (clk), .D (signal_4332), .Q (signal_23553) ) ;
    buf_clk cell_18673 ( .C (clk), .D (signal_7709), .Q (signal_23561) ) ;
    buf_clk cell_18681 ( .C (clk), .D (signal_4333), .Q (signal_23569) ) ;
    buf_clk cell_18689 ( .C (clk), .D (signal_7706), .Q (signal_23577) ) ;
    buf_clk cell_18697 ( .C (clk), .D (signal_4334), .Q (signal_23585) ) ;
    buf_clk cell_18705 ( .C (clk), .D (signal_7703), .Q (signal_23593) ) ;
    buf_clk cell_18713 ( .C (clk), .D (signal_4335), .Q (signal_23601) ) ;
    buf_clk cell_18721 ( .C (clk), .D (signal_7700), .Q (signal_23609) ) ;
    buf_clk cell_18729 ( .C (clk), .D (signal_4336), .Q (signal_23617) ) ;
    buf_clk cell_18737 ( .C (clk), .D (signal_7697), .Q (signal_23625) ) ;
    buf_clk cell_18749 ( .C (clk), .D (signal_4369), .Q (signal_23637) ) ;
    buf_clk cell_18757 ( .C (clk), .D (signal_7838), .Q (signal_23645) ) ;
    buf_clk cell_18765 ( .C (clk), .D (signal_4371), .Q (signal_23653) ) ;
    buf_clk cell_18773 ( .C (clk), .D (signal_7796), .Q (signal_23661) ) ;
    buf_clk cell_18781 ( .C (clk), .D (signal_4372), .Q (signal_23669) ) ;
    buf_clk cell_18789 ( .C (clk), .D (signal_7763), .Q (signal_23677) ) ;
    buf_clk cell_18797 ( .C (clk), .D (signal_4373), .Q (signal_23685) ) ;
    buf_clk cell_18805 ( .C (clk), .D (signal_7742), .Q (signal_23693) ) ;
    buf_clk cell_18813 ( .C (clk), .D (signal_4374), .Q (signal_23701) ) ;
    buf_clk cell_18821 ( .C (clk), .D (signal_7721), .Q (signal_23709) ) ;
    buf_clk cell_18829 ( .C (clk), .D (signal_4375), .Q (signal_23717) ) ;
    buf_clk cell_18837 ( .C (clk), .D (signal_7688), .Q (signal_23725) ) ;
    buf_clk cell_18845 ( .C (clk), .D (signal_4376), .Q (signal_23733) ) ;
    buf_clk cell_18853 ( .C (clk), .D (signal_7655), .Q (signal_23741) ) ;
    buf_clk cell_18861 ( .C (clk), .D (signal_4355), .Q (signal_23749) ) ;
    buf_clk cell_18869 ( .C (clk), .D (signal_7634), .Q (signal_23757) ) ;
    buf_clk cell_18877 ( .C (clk), .D (signal_4356), .Q (signal_23765) ) ;
    buf_clk cell_18885 ( .C (clk), .D (signal_7631), .Q (signal_23773) ) ;
    buf_clk cell_18893 ( .C (clk), .D (signal_4357), .Q (signal_23781) ) ;
    buf_clk cell_18901 ( .C (clk), .D (signal_7628), .Q (signal_23789) ) ;
    buf_clk cell_18909 ( .C (clk), .D (signal_4358), .Q (signal_23797) ) ;
    buf_clk cell_18917 ( .C (clk), .D (signal_7625), .Q (signal_23805) ) ;
    buf_clk cell_18925 ( .C (clk), .D (signal_4377), .Q (signal_23813) ) ;
    buf_clk cell_18933 ( .C (clk), .D (signal_7622), .Q (signal_23821) ) ;
    buf_clk cell_18941 ( .C (clk), .D (signal_4359), .Q (signal_23829) ) ;
    buf_clk cell_18949 ( .C (clk), .D (signal_7619), .Q (signal_23837) ) ;
    buf_clk cell_18957 ( .C (clk), .D (signal_4360), .Q (signal_23845) ) ;
    buf_clk cell_18965 ( .C (clk), .D (signal_7616), .Q (signal_23853) ) ;
    buf_clk cell_18973 ( .C (clk), .D (signal_4361), .Q (signal_23861) ) ;
    buf_clk cell_18981 ( .C (clk), .D (signal_7613), .Q (signal_23869) ) ;
    buf_clk cell_18989 ( .C (clk), .D (signal_4363), .Q (signal_23877) ) ;
    buf_clk cell_18997 ( .C (clk), .D (signal_7607), .Q (signal_23885) ) ;
    buf_clk cell_19005 ( .C (clk), .D (signal_4364), .Q (signal_23893) ) ;
    buf_clk cell_19013 ( .C (clk), .D (signal_7604), .Q (signal_23901) ) ;
    buf_clk cell_19021 ( .C (clk), .D (signal_4365), .Q (signal_23909) ) ;
    buf_clk cell_19029 ( .C (clk), .D (signal_7601), .Q (signal_23917) ) ;
    buf_clk cell_19037 ( .C (clk), .D (signal_4366), .Q (signal_23925) ) ;
    buf_clk cell_19045 ( .C (clk), .D (signal_7598), .Q (signal_23933) ) ;
    buf_clk cell_19053 ( .C (clk), .D (signal_4367), .Q (signal_23941) ) ;
    buf_clk cell_19061 ( .C (clk), .D (signal_7595), .Q (signal_23949) ) ;
    buf_clk cell_19069 ( .C (clk), .D (signal_4368), .Q (signal_23957) ) ;
    buf_clk cell_19077 ( .C (clk), .D (signal_7562), .Q (signal_23965) ) ;
    buf_clk cell_19085 ( .C (clk), .D (signal_3612), .Q (signal_23973) ) ;
    buf_clk cell_19093 ( .C (clk), .D (signal_3610), .Q (signal_23981) ) ;
    buf_clk cell_19101 ( .C (clk), .D (signal_3607), .Q (signal_23989) ) ;
    buf_clk cell_19109 ( .C (clk), .D (signal_3608), .Q (signal_23997) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4569 ( .a ({signal_8073, signal_4689}), .b ({signal_8075, signal_4691}), .clk (clk), .r (Fresh[0]), .c ({signal_8253, signal_4805}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4570 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_8078, signal_4694}), .clk (clk), .r (Fresh[1]), .c ({signal_8254, signal_4806}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4571 ( .a ({signal_7883, signal_4551}), .b ({signal_8077, signal_4693}), .clk (clk), .r (Fresh[2]), .c ({signal_8255, signal_4807}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4572 ( .a ({signal_8074, signal_4690}), .b ({signal_8079, signal_4695}), .clk (clk), .r (Fresh[3]), .c ({signal_8256, signal_4808}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4573 ( .a ({signal_7881, signal_4549}), .b ({signal_8076, signal_4692}), .clk (clk), .r (Fresh[4]), .c ({signal_8257, signal_4809}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4574 ( .a ({signal_7884, signal_4552}), .b ({signal_8080, signal_4696}), .clk (clk), .r (Fresh[5]), .c ({signal_8258, signal_4810}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4575 ( .a ({signal_8081, signal_4727}), .b ({signal_8083, signal_4729}), .clk (clk), .r (Fresh[6]), .c ({signal_8259, signal_4811}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4576 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_8086, signal_4732}), .clk (clk), .r (Fresh[7]), .c ({signal_8260, signal_4812}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4577 ( .a ({signal_7893, signal_4561}), .b ({signal_8085, signal_4731}), .clk (clk), .r (Fresh[8]), .c ({signal_8261, signal_4813}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4578 ( .a ({signal_8082, signal_4728}), .b ({signal_8087, signal_4733}), .clk (clk), .r (Fresh[9]), .c ({signal_8262, signal_4814}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4579 ( .a ({signal_7891, signal_4559}), .b ({signal_8084, signal_4730}), .clk (clk), .r (Fresh[10]), .c ({signal_8263, signal_4815}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4580 ( .a ({signal_7894, signal_4562}), .b ({signal_8088, signal_4734}), .clk (clk), .r (Fresh[11]), .c ({signal_8264, signal_4816}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4581 ( .a ({signal_8089, signal_4765}), .b ({signal_8091, signal_4767}), .clk (clk), .r (Fresh[12]), .c ({signal_8265, signal_4817}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4582 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_8094, signal_4770}), .clk (clk), .r (Fresh[13]), .c ({signal_8266, signal_4818}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4583 ( .a ({signal_7903, signal_4571}), .b ({signal_8093, signal_4769}), .clk (clk), .r (Fresh[14]), .c ({signal_8267, signal_4819}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4584 ( .a ({signal_8090, signal_4766}), .b ({signal_8095, signal_4771}), .clk (clk), .r (Fresh[15]), .c ({signal_8268, signal_4820}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4585 ( .a ({signal_7901, signal_4569}), .b ({signal_8092, signal_4768}), .clk (clk), .r (Fresh[16]), .c ({signal_8269, signal_4821}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4586 ( .a ({signal_7904, signal_4572}), .b ({signal_8096, signal_4772}), .clk (clk), .r (Fresh[17]), .c ({signal_8270, signal_4822}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4587 ( .a ({signal_8041, signal_4773}), .b ({signal_8043, signal_4775}), .clk (clk), .r (Fresh[18]), .c ({signal_8097, signal_4823}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4588 ( .a ({signal_7610, signal_4362}), .b ({signal_8046, signal_4778}), .clk (clk), .r (Fresh[19]), .c ({signal_8098, signal_4824}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4589 ( .a ({signal_7843, signal_4581}), .b ({signal_8045, signal_4777}), .clk (clk), .r (Fresh[20]), .c ({signal_8099, signal_4825}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4590 ( .a ({signal_8042, signal_4774}), .b ({signal_8047, signal_4779}), .clk (clk), .r (Fresh[21]), .c ({signal_8100, signal_4826}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4591 ( .a ({signal_7841, signal_4579}), .b ({signal_8044, signal_4776}), .clk (clk), .r (Fresh[22]), .c ({signal_8101, signal_4827}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4592 ( .a ({signal_7844, signal_4582}), .b ({signal_8048, signal_4780}), .clk (clk), .r (Fresh[23]), .c ({signal_8102, signal_4828}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4593 ( .a ({signal_8049, signal_4781}), .b ({signal_8051, signal_4783}), .clk (clk), .r (Fresh[24]), .c ({signal_8103, signal_4829}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4594 ( .a ({signal_7823, signal_4370}), .b ({signal_8054, signal_4786}), .clk (clk), .r (Fresh[25]), .c ({signal_8104, signal_4830}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4595 ( .a ({signal_7853, signal_4591}), .b ({signal_8053, signal_4785}), .clk (clk), .r (Fresh[26]), .c ({signal_8105, signal_4831}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4596 ( .a ({signal_8050, signal_4782}), .b ({signal_8055, signal_4787}), .clk (clk), .r (Fresh[27]), .c ({signal_8106, signal_4832}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4597 ( .a ({signal_7851, signal_4589}), .b ({signal_8052, signal_4784}), .clk (clk), .r (Fresh[28]), .c ({signal_8107, signal_4833}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4598 ( .a ({signal_7854, signal_4592}), .b ({signal_8056, signal_4788}), .clk (clk), .r (Fresh[29]), .c ({signal_8108, signal_4834}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4599 ( .a ({signal_8057, signal_4789}), .b ({signal_8059, signal_4791}), .clk (clk), .r (Fresh[30]), .c ({signal_8109, signal_4835}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4600 ( .a ({signal_7529, signal_4378}), .b ({signal_8062, signal_4794}), .clk (clk), .r (Fresh[31]), .c ({signal_8110, signal_4836}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4601 ( .a ({signal_7863, signal_4601}), .b ({signal_8061, signal_4793}), .clk (clk), .r (Fresh[32]), .c ({signal_8111, signal_4837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4602 ( .a ({signal_8058, signal_4790}), .b ({signal_8063, signal_4795}), .clk (clk), .r (Fresh[33]), .c ({signal_8112, signal_4838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4603 ( .a ({signal_7861, signal_4599}), .b ({signal_8060, signal_4792}), .clk (clk), .r (Fresh[34]), .c ({signal_8113, signal_4839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4604 ( .a ({signal_7864, signal_4602}), .b ({signal_8064, signal_4796}), .clk (clk), .r (Fresh[35]), .c ({signal_8114, signal_4840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4605 ( .a ({signal_8065, signal_4797}), .b ({signal_8067, signal_4799}), .clk (clk), .r (Fresh[36]), .c ({signal_8115, signal_4841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4606 ( .a ({signal_7637, signal_4354}), .b ({signal_8070, signal_4802}), .clk (clk), .r (Fresh[37]), .c ({signal_8116, signal_4842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4607 ( .a ({signal_7873, signal_4611}), .b ({signal_8069, signal_4801}), .clk (clk), .r (Fresh[38]), .c ({signal_8117, signal_4843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4608 ( .a ({signal_8066, signal_4798}), .b ({signal_8071, signal_4803}), .clk (clk), .r (Fresh[39]), .c ({signal_8118, signal_4844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4609 ( .a ({signal_7871, signal_4609}), .b ({signal_8068, signal_4800}), .clk (clk), .r (Fresh[40]), .c ({signal_8119, signal_4845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4610 ( .a ({signal_7874, signal_4612}), .b ({signal_8072, signal_4804}), .clk (clk), .r (Fresh[41]), .c ({signal_8120, signal_4846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4764 ( .a ({signal_8121, signal_4847}), .b ({signal_8123, signal_4849}), .clk (clk), .r (Fresh[42]), .c ({signal_8292, signal_5000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4765 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_8126, signal_4852}), .clk (clk), .r (Fresh[43]), .c ({signal_8293, signal_5001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4766 ( .a ({signal_7913, signal_4621}), .b ({signal_8125, signal_4851}), .clk (clk), .r (Fresh[44]), .c ({signal_8294, signal_5002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4767 ( .a ({signal_8122, signal_4848}), .b ({signal_8127, signal_4853}), .clk (clk), .r (Fresh[45]), .c ({signal_8295, signal_5003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4768 ( .a ({signal_7911, signal_4619}), .b ({signal_8124, signal_4850}), .clk (clk), .r (Fresh[46]), .c ({signal_8296, signal_5004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4769 ( .a ({signal_7914, signal_4622}), .b ({signal_8128, signal_4854}), .clk (clk), .r (Fresh[47]), .c ({signal_8297, signal_5005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4770 ( .a ({signal_8129, signal_4855}), .b ({signal_8131, signal_4857}), .clk (clk), .r (Fresh[48]), .c ({signal_8298, signal_5006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4771 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_8134, signal_4860}), .clk (clk), .r (Fresh[49]), .c ({signal_8299, signal_5007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4772 ( .a ({signal_7923, signal_4631}), .b ({signal_8133, signal_4859}), .clk (clk), .r (Fresh[50]), .c ({signal_8300, signal_5008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4773 ( .a ({signal_8130, signal_4856}), .b ({signal_8135, signal_4861}), .clk (clk), .r (Fresh[51]), .c ({signal_8301, signal_5009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4774 ( .a ({signal_7921, signal_4629}), .b ({signal_8132, signal_4858}), .clk (clk), .r (Fresh[52]), .c ({signal_8302, signal_5010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4775 ( .a ({signal_7924, signal_4632}), .b ({signal_8136, signal_4862}), .clk (clk), .r (Fresh[53]), .c ({signal_8303, signal_5011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4776 ( .a ({signal_8137, signal_4863}), .b ({signal_8139, signal_4865}), .clk (clk), .r (Fresh[54]), .c ({signal_8304, signal_5012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4777 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_8142, signal_4868}), .clk (clk), .r (Fresh[55]), .c ({signal_8305, signal_5013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4778 ( .a ({signal_7933, signal_4641}), .b ({signal_8141, signal_4867}), .clk (clk), .r (Fresh[56]), .c ({signal_8306, signal_5014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4779 ( .a ({signal_8138, signal_4864}), .b ({signal_8143, signal_4869}), .clk (clk), .r (Fresh[57]), .c ({signal_8307, signal_5015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4780 ( .a ({signal_7931, signal_4639}), .b ({signal_8140, signal_4866}), .clk (clk), .r (Fresh[58]), .c ({signal_8308, signal_5016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4781 ( .a ({signal_7934, signal_4642}), .b ({signal_8144, signal_4870}), .clk (clk), .r (Fresh[59]), .c ({signal_8309, signal_5017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4782 ( .a ({signal_8145, signal_4871}), .b ({signal_8147, signal_4873}), .clk (clk), .r (Fresh[60]), .c ({signal_8310, signal_5018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4783 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_8150, signal_4876}), .clk (clk), .r (Fresh[61]), .c ({signal_8311, signal_5019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4784 ( .a ({signal_7943, signal_4651}), .b ({signal_8149, signal_4875}), .clk (clk), .r (Fresh[62]), .c ({signal_8312, signal_5020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4785 ( .a ({signal_8146, signal_4872}), .b ({signal_8151, signal_4877}), .clk (clk), .r (Fresh[63]), .c ({signal_8313, signal_5021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4786 ( .a ({signal_7941, signal_4649}), .b ({signal_8148, signal_4874}), .clk (clk), .r (Fresh[64]), .c ({signal_8314, signal_5022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4787 ( .a ({signal_7944, signal_4652}), .b ({signal_8152, signal_4878}), .clk (clk), .r (Fresh[65]), .c ({signal_8315, signal_5023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4788 ( .a ({signal_8153, signal_4879}), .b ({signal_8155, signal_4881}), .clk (clk), .r (Fresh[66]), .c ({signal_8316, signal_5024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4789 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_8158, signal_4884}), .clk (clk), .r (Fresh[67]), .c ({signal_8317, signal_5025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4790 ( .a ({signal_7953, signal_4661}), .b ({signal_8157, signal_4883}), .clk (clk), .r (Fresh[68]), .c ({signal_8318, signal_5026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4791 ( .a ({signal_8154, signal_4880}), .b ({signal_8159, signal_4885}), .clk (clk), .r (Fresh[69]), .c ({signal_8319, signal_5027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4792 ( .a ({signal_7951, signal_4659}), .b ({signal_8156, signal_4882}), .clk (clk), .r (Fresh[70]), .c ({signal_8320, signal_5028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4793 ( .a ({signal_7954, signal_4662}), .b ({signal_8160, signal_4886}), .clk (clk), .r (Fresh[71]), .c ({signal_8321, signal_5029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4794 ( .a ({signal_8161, signal_4887}), .b ({signal_8163, signal_4889}), .clk (clk), .r (Fresh[72]), .c ({signal_8322, signal_5030}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4795 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_8166, signal_4892}), .clk (clk), .r (Fresh[73]), .c ({signal_8323, signal_5031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4796 ( .a ({signal_7963, signal_4671}), .b ({signal_8165, signal_4891}), .clk (clk), .r (Fresh[74]), .c ({signal_8324, signal_5032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4797 ( .a ({signal_8162, signal_4888}), .b ({signal_8167, signal_4893}), .clk (clk), .r (Fresh[75]), .c ({signal_8325, signal_5033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4798 ( .a ({signal_7961, signal_4669}), .b ({signal_8164, signal_4890}), .clk (clk), .r (Fresh[76]), .c ({signal_8326, signal_5034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4799 ( .a ({signal_7964, signal_4672}), .b ({signal_8168, signal_4894}), .clk (clk), .r (Fresh[77]), .c ({signal_8327, signal_5035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4800 ( .a ({signal_8169, signal_4895}), .b ({signal_8171, signal_4897}), .clk (clk), .r (Fresh[78]), .c ({signal_8328, signal_5036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4801 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_8174, signal_4900}), .clk (clk), .r (Fresh[79]), .c ({signal_8329, signal_5037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4802 ( .a ({signal_7973, signal_4681}), .b ({signal_8173, signal_4899}), .clk (clk), .r (Fresh[80]), .c ({signal_8330, signal_5038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4803 ( .a ({signal_8170, signal_4896}), .b ({signal_8175, signal_4901}), .clk (clk), .r (Fresh[81]), .c ({signal_8331, signal_5039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4804 ( .a ({signal_7971, signal_4679}), .b ({signal_8172, signal_4898}), .clk (clk), .r (Fresh[82]), .c ({signal_8332, signal_5040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4805 ( .a ({signal_7974, signal_4682}), .b ({signal_8176, signal_4902}), .clk (clk), .r (Fresh[83]), .c ({signal_8333, signal_5041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4806 ( .a ({signal_8271, signal_4903}), .b ({signal_8276, signal_4908}), .clk (clk), .r (Fresh[84]), .c ({signal_8497, signal_5042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4807 ( .a ({signal_8274, signal_4906}), .b ({signal_8275, signal_4907}), .clk (clk), .r (Fresh[85]), .c ({signal_8498, signal_5043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4808 ( .a ({signal_7882, signal_4550}), .b ({signal_8272, signal_4904}), .clk (clk), .r (Fresh[86]), .c ({signal_8499, signal_5044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4809 ( .a ({signal_8177, signal_4910}), .b ({signal_8179, signal_4912}), .clk (clk), .r (Fresh[87]), .c ({signal_8334, signal_5045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4810 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_8182, signal_4915}), .clk (clk), .r (Fresh[88]), .c ({signal_8335, signal_5046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4811 ( .a ({signal_7983, signal_4699}), .b ({signal_8181, signal_4914}), .clk (clk), .r (Fresh[89]), .c ({signal_8336, signal_5047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4812 ( .a ({signal_8178, signal_4911}), .b ({signal_8183, signal_4916}), .clk (clk), .r (Fresh[90]), .c ({signal_8337, signal_5048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4813 ( .a ({signal_7981, signal_4697}), .b ({signal_8180, signal_4913}), .clk (clk), .r (Fresh[91]), .c ({signal_8338, signal_5049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4814 ( .a ({signal_7984, signal_4700}), .b ({signal_8184, signal_4917}), .clk (clk), .r (Fresh[92]), .c ({signal_8339, signal_5050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4815 ( .a ({signal_8185, signal_4918}), .b ({signal_8187, signal_4920}), .clk (clk), .r (Fresh[93]), .c ({signal_8340, signal_5051}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4816 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_8190, signal_4923}), .clk (clk), .r (Fresh[94]), .c ({signal_8341, signal_5052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4817 ( .a ({signal_7993, signal_4709}), .b ({signal_8189, signal_4922}), .clk (clk), .r (Fresh[95]), .c ({signal_8342, signal_5053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4818 ( .a ({signal_8186, signal_4919}), .b ({signal_8191, signal_4924}), .clk (clk), .r (Fresh[96]), .c ({signal_8343, signal_5054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4819 ( .a ({signal_7991, signal_4707}), .b ({signal_8188, signal_4921}), .clk (clk), .r (Fresh[97]), .c ({signal_8344, signal_5055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4820 ( .a ({signal_7994, signal_4710}), .b ({signal_8192, signal_4925}), .clk (clk), .r (Fresh[98]), .c ({signal_8345, signal_5056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4821 ( .a ({signal_8193, signal_4926}), .b ({signal_8195, signal_4928}), .clk (clk), .r (Fresh[99]), .c ({signal_8346, signal_5057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4822 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8198, signal_4931}), .clk (clk), .r (Fresh[100]), .c ({signal_8347, signal_5058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4823 ( .a ({signal_8003, signal_4719}), .b ({signal_8197, signal_4930}), .clk (clk), .r (Fresh[101]), .c ({signal_8348, signal_5059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4824 ( .a ({signal_8194, signal_4927}), .b ({signal_8199, signal_4932}), .clk (clk), .r (Fresh[102]), .c ({signal_8349, signal_5060}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4825 ( .a ({signal_8001, signal_4717}), .b ({signal_8196, signal_4929}), .clk (clk), .r (Fresh[103]), .c ({signal_8350, signal_5061}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4826 ( .a ({signal_8004, signal_4720}), .b ({signal_8200, signal_4933}), .clk (clk), .r (Fresh[104]), .c ({signal_8351, signal_5062}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4827 ( .a ({signal_8278, signal_4934}), .b ({signal_8283, signal_4939}), .clk (clk), .r (Fresh[105]), .c ({signal_8500, signal_5063}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4828 ( .a ({signal_8281, signal_4937}), .b ({signal_8282, signal_4938}), .clk (clk), .r (Fresh[106]), .c ({signal_8501, signal_5064}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4829 ( .a ({signal_7892, signal_4560}), .b ({signal_8279, signal_4935}), .clk (clk), .r (Fresh[107]), .c ({signal_8502, signal_5065}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4830 ( .a ({signal_8201, signal_4941}), .b ({signal_8203, signal_4943}), .clk (clk), .r (Fresh[108]), .c ({signal_8352, signal_5066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4831 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8206, signal_4946}), .clk (clk), .r (Fresh[109]), .c ({signal_8353, signal_5067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4832 ( .a ({signal_8013, signal_4737}), .b ({signal_8205, signal_4945}), .clk (clk), .r (Fresh[110]), .c ({signal_8354, signal_5068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4833 ( .a ({signal_8202, signal_4942}), .b ({signal_8207, signal_4947}), .clk (clk), .r (Fresh[111]), .c ({signal_8355, signal_5069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4834 ( .a ({signal_8011, signal_4735}), .b ({signal_8204, signal_4944}), .clk (clk), .r (Fresh[112]), .c ({signal_8356, signal_5070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4835 ( .a ({signal_8014, signal_4738}), .b ({signal_8208, signal_4948}), .clk (clk), .r (Fresh[113]), .c ({signal_8357, signal_5071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4836 ( .a ({signal_8209, signal_4949}), .b ({signal_8211, signal_4951}), .clk (clk), .r (Fresh[114]), .c ({signal_8358, signal_5072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4837 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8214, signal_4954}), .clk (clk), .r (Fresh[115]), .c ({signal_8359, signal_5073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4838 ( .a ({signal_8023, signal_4747}), .b ({signal_8213, signal_4953}), .clk (clk), .r (Fresh[116]), .c ({signal_8360, signal_5074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4839 ( .a ({signal_8210, signal_4950}), .b ({signal_8215, signal_4955}), .clk (clk), .r (Fresh[117]), .c ({signal_8361, signal_5075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4840 ( .a ({signal_8021, signal_4745}), .b ({signal_8212, signal_4952}), .clk (clk), .r (Fresh[118]), .c ({signal_8362, signal_5076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4841 ( .a ({signal_8024, signal_4748}), .b ({signal_8216, signal_4956}), .clk (clk), .r (Fresh[119]), .c ({signal_8363, signal_5077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4842 ( .a ({signal_8217, signal_4957}), .b ({signal_8219, signal_4959}), .clk (clk), .r (Fresh[120]), .c ({signal_8364, signal_5078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4843 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8222, signal_4962}), .clk (clk), .r (Fresh[121]), .c ({signal_8365, signal_5079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4844 ( .a ({signal_8033, signal_4757}), .b ({signal_8221, signal_4961}), .clk (clk), .r (Fresh[122]), .c ({signal_8366, signal_5080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4845 ( .a ({signal_8218, signal_4958}), .b ({signal_8223, signal_4963}), .clk (clk), .r (Fresh[123]), .c ({signal_8367, signal_5081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4846 ( .a ({signal_8031, signal_4755}), .b ({signal_8220, signal_4960}), .clk (clk), .r (Fresh[124]), .c ({signal_8368, signal_5082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4847 ( .a ({signal_8034, signal_4758}), .b ({signal_8224, signal_4964}), .clk (clk), .r (Fresh[125]), .c ({signal_8369, signal_5083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4848 ( .a ({signal_8285, signal_4965}), .b ({signal_8290, signal_4970}), .clk (clk), .r (Fresh[126]), .c ({signal_8503, signal_5084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4849 ( .a ({signal_8288, signal_4968}), .b ({signal_8289, signal_4969}), .clk (clk), .r (Fresh[127]), .c ({signal_8504, signal_5085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4850 ( .a ({signal_7902, signal_4570}), .b ({signal_8286, signal_4966}), .clk (clk), .r (Fresh[128]), .c ({signal_8505, signal_5086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4851 ( .a ({signal_8225, signal_4972}), .b ({signal_8230, signal_4977}), .clk (clk), .r (Fresh[129]), .c ({signal_8370, signal_5087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4852 ( .a ({signal_8228, signal_4975}), .b ({signal_8229, signal_4976}), .clk (clk), .r (Fresh[130]), .c ({signal_8371, signal_5088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4853 ( .a ({signal_7842, signal_4580}), .b ({signal_8226, signal_4973}), .clk (clk), .r (Fresh[131]), .c ({signal_8372, signal_5089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4854 ( .a ({signal_8232, signal_4979}), .b ({signal_8237, signal_4984}), .clk (clk), .r (Fresh[132]), .c ({signal_8373, signal_5090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4855 ( .a ({signal_8235, signal_4982}), .b ({signal_8236, signal_4983}), .clk (clk), .r (Fresh[133]), .c ({signal_8374, signal_5091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4856 ( .a ({signal_7852, signal_4590}), .b ({signal_8233, signal_4980}), .clk (clk), .r (Fresh[134]), .c ({signal_8375, signal_5092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4857 ( .a ({signal_8239, signal_4986}), .b ({signal_8244, signal_4991}), .clk (clk), .r (Fresh[135]), .c ({signal_8376, signal_5093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4858 ( .a ({signal_8242, signal_4989}), .b ({signal_8243, signal_4990}), .clk (clk), .r (Fresh[136]), .c ({signal_8377, signal_5094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4859 ( .a ({signal_7862, signal_4600}), .b ({signal_8240, signal_4987}), .clk (clk), .r (Fresh[137]), .c ({signal_8378, signal_5095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4860 ( .a ({signal_8246, signal_4993}), .b ({signal_8251, signal_4998}), .clk (clk), .r (Fresh[138]), .c ({signal_8379, signal_5096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4861 ( .a ({signal_8249, signal_4996}), .b ({signal_8250, signal_4997}), .clk (clk), .r (Fresh[139]), .c ({signal_8380, signal_5097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4862 ( .a ({signal_7872, signal_4610}), .b ({signal_8247, signal_4994}), .clk (clk), .r (Fresh[140]), .c ({signal_8381, signal_5098}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4914 ( .a ({signal_12472, signal_12470}), .b ({signal_8253, signal_4805}), .c ({signal_8508, signal_5150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4915 ( .a ({signal_8253, signal_4805}), .b ({signal_8254, signal_4806}), .c ({signal_8509, signal_5151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4916 ( .a ({signal_12476, signal_12474}), .b ({signal_8255, signal_4807}), .c ({signal_8510, signal_5152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4917 ( .a ({signal_8257, signal_4809}), .b ({signal_8258, signal_4810}), .c ({signal_8511, signal_5153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4941 ( .a ({signal_12480, signal_12478}), .b ({signal_8259, signal_4811}), .c ({signal_8514, signal_5177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4942 ( .a ({signal_8259, signal_4811}), .b ({signal_8260, signal_4812}), .c ({signal_8515, signal_5178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4943 ( .a ({signal_12484, signal_12482}), .b ({signal_8261, signal_4813}), .c ({signal_8516, signal_5179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4944 ( .a ({signal_8263, signal_4815}), .b ({signal_8264, signal_4816}), .c ({signal_8517, signal_5180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4968 ( .a ({signal_12488, signal_12486}), .b ({signal_8265, signal_4817}), .c ({signal_8520, signal_5204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4969 ( .a ({signal_8265, signal_4817}), .b ({signal_8266, signal_4818}), .c ({signal_8521, signal_5205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4970 ( .a ({signal_12492, signal_12490}), .b ({signal_8267, signal_4819}), .c ({signal_8522, signal_5206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4971 ( .a ({signal_8269, signal_4821}), .b ({signal_8270, signal_4822}), .c ({signal_8523, signal_5207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4974 ( .a ({signal_12496, signal_12494}), .b ({signal_8097, signal_4823}), .c ({signal_8475, signal_5210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4975 ( .a ({signal_8097, signal_4823}), .b ({signal_8098, signal_4824}), .c ({signal_8476, signal_5211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4976 ( .a ({signal_12500, signal_12498}), .b ({signal_8099, signal_4825}), .c ({signal_8477, signal_5212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4977 ( .a ({signal_8101, signal_4827}), .b ({signal_8102, signal_4828}), .c ({signal_8478, signal_5213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4980 ( .a ({signal_12504, signal_12502}), .b ({signal_8103, signal_4829}), .c ({signal_8481, signal_5216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4981 ( .a ({signal_8103, signal_4829}), .b ({signal_8104, signal_4830}), .c ({signal_8482, signal_5217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4982 ( .a ({signal_12508, signal_12506}), .b ({signal_8105, signal_4831}), .c ({signal_8483, signal_5218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4983 ( .a ({signal_8107, signal_4833}), .b ({signal_8108, signal_4834}), .c ({signal_8484, signal_5219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4986 ( .a ({signal_12512, signal_12510}), .b ({signal_8109, signal_4835}), .c ({signal_8487, signal_5222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4987 ( .a ({signal_8109, signal_4835}), .b ({signal_8110, signal_4836}), .c ({signal_8488, signal_5223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4988 ( .a ({signal_12516, signal_12514}), .b ({signal_8111, signal_4837}), .c ({signal_8489, signal_5224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4989 ( .a ({signal_8113, signal_4839}), .b ({signal_8114, signal_4840}), .c ({signal_8490, signal_5225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4992 ( .a ({signal_12520, signal_12518}), .b ({signal_8115, signal_4841}), .c ({signal_8493, signal_5228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4993 ( .a ({signal_8115, signal_4841}), .b ({signal_8116, signal_4842}), .c ({signal_8494, signal_5229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4994 ( .a ({signal_12524, signal_12522}), .b ({signal_8117, signal_4843}), .c ({signal_8495, signal_5230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4995 ( .a ({signal_8119, signal_4845}), .b ({signal_8120, signal_4846}), .c ({signal_8496, signal_5231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4996 ( .a ({signal_8382, signal_5099}), .b ({signal_8387, signal_5104}), .clk (clk), .r (Fresh[141]), .c ({signal_8524, signal_5232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4997 ( .a ({signal_8385, signal_5102}), .b ({signal_8386, signal_5103}), .clk (clk), .r (Fresh[142]), .c ({signal_8525, signal_5233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4998 ( .a ({signal_7912, signal_4620}), .b ({signal_8383, signal_5100}), .clk (clk), .r (Fresh[143]), .c ({signal_8526, signal_5234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_4999 ( .a ({signal_8389, signal_5106}), .b ({signal_8394, signal_5111}), .clk (clk), .r (Fresh[144]), .c ({signal_8527, signal_5235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5000 ( .a ({signal_8392, signal_5109}), .b ({signal_8393, signal_5110}), .clk (clk), .r (Fresh[145]), .c ({signal_8528, signal_5236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5001 ( .a ({signal_7922, signal_4630}), .b ({signal_8390, signal_5107}), .clk (clk), .r (Fresh[146]), .c ({signal_8529, signal_5237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5002 ( .a ({signal_8396, signal_5113}), .b ({signal_8401, signal_5118}), .clk (clk), .r (Fresh[147]), .c ({signal_8530, signal_5238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5003 ( .a ({signal_8399, signal_5116}), .b ({signal_8400, signal_5117}), .clk (clk), .r (Fresh[148]), .c ({signal_8531, signal_5239}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5004 ( .a ({signal_7932, signal_4640}), .b ({signal_8397, signal_5114}), .clk (clk), .r (Fresh[149]), .c ({signal_8532, signal_5240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5005 ( .a ({signal_8403, signal_5120}), .b ({signal_8408, signal_5125}), .clk (clk), .r (Fresh[150]), .c ({signal_8533, signal_5241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5006 ( .a ({signal_8406, signal_5123}), .b ({signal_8407, signal_5124}), .clk (clk), .r (Fresh[151]), .c ({signal_8534, signal_5242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5007 ( .a ({signal_7942, signal_4650}), .b ({signal_8404, signal_5121}), .clk (clk), .r (Fresh[152]), .c ({signal_8535, signal_5243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5008 ( .a ({signal_8410, signal_5127}), .b ({signal_8415, signal_5132}), .clk (clk), .r (Fresh[153]), .c ({signal_8536, signal_5244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5009 ( .a ({signal_8413, signal_5130}), .b ({signal_8414, signal_5131}), .clk (clk), .r (Fresh[154]), .c ({signal_8537, signal_5245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5010 ( .a ({signal_7952, signal_4660}), .b ({signal_8411, signal_5128}), .clk (clk), .r (Fresh[155]), .c ({signal_8538, signal_5246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5011 ( .a ({signal_8417, signal_5134}), .b ({signal_8422, signal_5139}), .clk (clk), .r (Fresh[156]), .c ({signal_8539, signal_5247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5012 ( .a ({signal_8420, signal_5137}), .b ({signal_8421, signal_5138}), .clk (clk), .r (Fresh[157]), .c ({signal_8540, signal_5248}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5013 ( .a ({signal_7962, signal_4670}), .b ({signal_8418, signal_5135}), .clk (clk), .r (Fresh[158]), .c ({signal_8541, signal_5249}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5014 ( .a ({signal_8424, signal_5141}), .b ({signal_8429, signal_5146}), .clk (clk), .r (Fresh[159]), .c ({signal_8542, signal_5250}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5015 ( .a ({signal_8427, signal_5144}), .b ({signal_8428, signal_5145}), .clk (clk), .r (Fresh[160]), .c ({signal_8543, signal_5251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5016 ( .a ({signal_7972, signal_4680}), .b ({signal_8425, signal_5142}), .clk (clk), .r (Fresh[161]), .c ({signal_8544, signal_5252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5017 ( .a ({signal_8431, signal_5154}), .b ({signal_8436, signal_5159}), .clk (clk), .r (Fresh[162]), .c ({signal_8545, signal_5253}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5018 ( .a ({signal_8434, signal_5157}), .b ({signal_8435, signal_5158}), .clk (clk), .r (Fresh[163]), .c ({signal_8546, signal_5254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5019 ( .a ({signal_7982, signal_4698}), .b ({signal_8432, signal_5155}), .clk (clk), .r (Fresh[164]), .c ({signal_8547, signal_5255}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5020 ( .a ({signal_8438, signal_5161}), .b ({signal_8443, signal_5166}), .clk (clk), .r (Fresh[165]), .c ({signal_8548, signal_5256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5021 ( .a ({signal_8441, signal_5164}), .b ({signal_8442, signal_5165}), .clk (clk), .r (Fresh[166]), .c ({signal_8549, signal_5257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5022 ( .a ({signal_7992, signal_4708}), .b ({signal_8439, signal_5162}), .clk (clk), .r (Fresh[167]), .c ({signal_8550, signal_5258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5023 ( .a ({signal_8445, signal_5168}), .b ({signal_8450, signal_5173}), .clk (clk), .r (Fresh[168]), .c ({signal_8551, signal_5259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5024 ( .a ({signal_8448, signal_5171}), .b ({signal_8449, signal_5172}), .clk (clk), .r (Fresh[169]), .c ({signal_8552, signal_5260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5025 ( .a ({signal_8002, signal_4718}), .b ({signal_8446, signal_5169}), .clk (clk), .r (Fresh[170]), .c ({signal_8553, signal_5261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5026 ( .a ({signal_8452, signal_5181}), .b ({signal_8457, signal_5186}), .clk (clk), .r (Fresh[171]), .c ({signal_8554, signal_5262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5027 ( .a ({signal_8455, signal_5184}), .b ({signal_8456, signal_5185}), .clk (clk), .r (Fresh[172]), .c ({signal_8555, signal_5263}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5028 ( .a ({signal_8012, signal_4736}), .b ({signal_8453, signal_5182}), .clk (clk), .r (Fresh[173]), .c ({signal_8556, signal_5264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5029 ( .a ({signal_8459, signal_5188}), .b ({signal_8464, signal_5193}), .clk (clk), .r (Fresh[174]), .c ({signal_8557, signal_5265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5030 ( .a ({signal_8462, signal_5191}), .b ({signal_8463, signal_5192}), .clk (clk), .r (Fresh[175]), .c ({signal_8558, signal_5266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5031 ( .a ({signal_8022, signal_4746}), .b ({signal_8460, signal_5189}), .clk (clk), .r (Fresh[176]), .c ({signal_8559, signal_5267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5032 ( .a ({signal_8466, signal_5195}), .b ({signal_8471, signal_5200}), .clk (clk), .r (Fresh[177]), .c ({signal_8560, signal_5268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5033 ( .a ({signal_8469, signal_5198}), .b ({signal_8470, signal_5199}), .clk (clk), .r (Fresh[178]), .c ({signal_8561, signal_5269}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5034 ( .a ({signal_8032, signal_4756}), .b ({signal_8467, signal_5196}), .clk (clk), .r (Fresh[179]), .c ({signal_8562, signal_5270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5037 ( .a ({signal_12528, signal_12526}), .b ({signal_8292, signal_5000}), .c ({signal_8565, signal_5273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5038 ( .a ({signal_8292, signal_5000}), .b ({signal_8293, signal_5001}), .c ({signal_8566, signal_5274}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5039 ( .a ({signal_12532, signal_12530}), .b ({signal_8294, signal_5002}), .c ({signal_8567, signal_5275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5040 ( .a ({signal_8296, signal_5004}), .b ({signal_8297, signal_5005}), .c ({signal_8568, signal_5276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5043 ( .a ({signal_12536, signal_12534}), .b ({signal_8298, signal_5006}), .c ({signal_8571, signal_5279}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5044 ( .a ({signal_8298, signal_5006}), .b ({signal_8299, signal_5007}), .c ({signal_8572, signal_5280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5045 ( .a ({signal_12540, signal_12538}), .b ({signal_8300, signal_5008}), .c ({signal_8573, signal_5281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5046 ( .a ({signal_8302, signal_5010}), .b ({signal_8303, signal_5011}), .c ({signal_8574, signal_5282}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5049 ( .a ({signal_12544, signal_12542}), .b ({signal_8304, signal_5012}), .c ({signal_8577, signal_5285}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5050 ( .a ({signal_8304, signal_5012}), .b ({signal_8305, signal_5013}), .c ({signal_8578, signal_5286}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5051 ( .a ({signal_12548, signal_12546}), .b ({signal_8306, signal_5014}), .c ({signal_8579, signal_5287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5052 ( .a ({signal_8308, signal_5016}), .b ({signal_8309, signal_5017}), .c ({signal_8580, signal_5288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5055 ( .a ({signal_12552, signal_12550}), .b ({signal_8310, signal_5018}), .c ({signal_8583, signal_5291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5056 ( .a ({signal_8310, signal_5018}), .b ({signal_8311, signal_5019}), .c ({signal_8584, signal_5292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5057 ( .a ({signal_12556, signal_12554}), .b ({signal_8312, signal_5020}), .c ({signal_8585, signal_5293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5058 ( .a ({signal_8314, signal_5022}), .b ({signal_8315, signal_5023}), .c ({signal_8586, signal_5294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5061 ( .a ({signal_12560, signal_12558}), .b ({signal_8316, signal_5024}), .c ({signal_8589, signal_5297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5062 ( .a ({signal_8316, signal_5024}), .b ({signal_8317, signal_5025}), .c ({signal_8590, signal_5298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5063 ( .a ({signal_12564, signal_12562}), .b ({signal_8318, signal_5026}), .c ({signal_8591, signal_5299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5064 ( .a ({signal_8320, signal_5028}), .b ({signal_8321, signal_5029}), .c ({signal_8592, signal_5300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5067 ( .a ({signal_12568, signal_12566}), .b ({signal_8322, signal_5030}), .c ({signal_8595, signal_5303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5068 ( .a ({signal_8322, signal_5030}), .b ({signal_8323, signal_5031}), .c ({signal_8596, signal_5304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5069 ( .a ({signal_12572, signal_12570}), .b ({signal_8324, signal_5032}), .c ({signal_8597, signal_5305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5070 ( .a ({signal_8326, signal_5034}), .b ({signal_8327, signal_5035}), .c ({signal_8598, signal_5306}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5073 ( .a ({signal_12576, signal_12574}), .b ({signal_8328, signal_5036}), .c ({signal_8601, signal_5309}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5074 ( .a ({signal_8328, signal_5036}), .b ({signal_8329, signal_5037}), .c ({signal_8602, signal_5310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5075 ( .a ({signal_12580, signal_12578}), .b ({signal_8330, signal_5038}), .c ({signal_8603, signal_5311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5076 ( .a ({signal_8332, signal_5040}), .b ({signal_8333, signal_5041}), .c ({signal_8604, signal_5312}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5077 ( .a ({signal_8255, signal_4807}), .b ({signal_8498, signal_5043}), .c ({signal_8661, signal_5313}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5078 ( .a ({signal_8257, signal_4809}), .b ({signal_8499, signal_5044}), .c ({signal_8662, signal_5314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5079 ( .a ({signal_8497, signal_5042}), .b ({signal_8508, signal_5150}), .c ({signal_8663, signal_5315}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5080 ( .a ({signal_12584, signal_12582}), .b ({signal_8509, signal_5151}), .c ({signal_8664, signal_5316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5081 ( .a ({signal_8256, signal_4808}), .b ({signal_8510, signal_5152}), .c ({signal_8665, signal_5317}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5084 ( .a ({signal_12588, signal_12586}), .b ({signal_8334, signal_5045}), .c ({signal_8607, signal_5320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5085 ( .a ({signal_8334, signal_5045}), .b ({signal_8335, signal_5046}), .c ({signal_8608, signal_5321}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5086 ( .a ({signal_12592, signal_12590}), .b ({signal_8336, signal_5047}), .c ({signal_8609, signal_5322}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5087 ( .a ({signal_8338, signal_5049}), .b ({signal_8339, signal_5050}), .c ({signal_8610, signal_5323}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5090 ( .a ({signal_12596, signal_12594}), .b ({signal_8340, signal_5051}), .c ({signal_8613, signal_5326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5091 ( .a ({signal_8340, signal_5051}), .b ({signal_8341, signal_5052}), .c ({signal_8614, signal_5327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5092 ( .a ({signal_12600, signal_12598}), .b ({signal_8342, signal_5053}), .c ({signal_8615, signal_5328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5093 ( .a ({signal_8344, signal_5055}), .b ({signal_8345, signal_5056}), .c ({signal_8616, signal_5329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5096 ( .a ({signal_12604, signal_12602}), .b ({signal_8346, signal_5057}), .c ({signal_8619, signal_5332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5097 ( .a ({signal_8346, signal_5057}), .b ({signal_8347, signal_5058}), .c ({signal_8620, signal_5333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5098 ( .a ({signal_12608, signal_12606}), .b ({signal_8348, signal_5059}), .c ({signal_8621, signal_5334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5099 ( .a ({signal_8350, signal_5061}), .b ({signal_8351, signal_5062}), .c ({signal_8622, signal_5335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5100 ( .a ({signal_8261, signal_4813}), .b ({signal_8501, signal_5064}), .c ({signal_8666, signal_5336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5101 ( .a ({signal_8263, signal_4815}), .b ({signal_8502, signal_5065}), .c ({signal_8667, signal_5337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5102 ( .a ({signal_8500, signal_5063}), .b ({signal_8514, signal_5177}), .c ({signal_8668, signal_5338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5103 ( .a ({signal_12612, signal_12610}), .b ({signal_8515, signal_5178}), .c ({signal_8669, signal_5339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5104 ( .a ({signal_8262, signal_4814}), .b ({signal_8516, signal_5179}), .c ({signal_8670, signal_5340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5107 ( .a ({signal_12616, signal_12614}), .b ({signal_8352, signal_5066}), .c ({signal_8625, signal_5343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5108 ( .a ({signal_8352, signal_5066}), .b ({signal_8353, signal_5067}), .c ({signal_8626, signal_5344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5109 ( .a ({signal_12620, signal_12618}), .b ({signal_8354, signal_5068}), .c ({signal_8627, signal_5345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5110 ( .a ({signal_8356, signal_5070}), .b ({signal_8357, signal_5071}), .c ({signal_8628, signal_5346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5113 ( .a ({signal_12624, signal_12622}), .b ({signal_8358, signal_5072}), .c ({signal_8631, signal_5349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5114 ( .a ({signal_8358, signal_5072}), .b ({signal_8359, signal_5073}), .c ({signal_8632, signal_5350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5115 ( .a ({signal_12628, signal_12626}), .b ({signal_8360, signal_5074}), .c ({signal_8633, signal_5351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5116 ( .a ({signal_8362, signal_5076}), .b ({signal_8363, signal_5077}), .c ({signal_8634, signal_5352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5119 ( .a ({signal_12632, signal_12630}), .b ({signal_8364, signal_5078}), .c ({signal_8637, signal_5355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5120 ( .a ({signal_8364, signal_5078}), .b ({signal_8365, signal_5079}), .c ({signal_8638, signal_5356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5121 ( .a ({signal_12636, signal_12634}), .b ({signal_8366, signal_5080}), .c ({signal_8639, signal_5357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5122 ( .a ({signal_8368, signal_5082}), .b ({signal_8369, signal_5083}), .c ({signal_8640, signal_5358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5123 ( .a ({signal_8267, signal_4819}), .b ({signal_8504, signal_5085}), .c ({signal_8671, signal_5359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5124 ( .a ({signal_8269, signal_4821}), .b ({signal_8505, signal_5086}), .c ({signal_8672, signal_5360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5125 ( .a ({signal_8503, signal_5084}), .b ({signal_8520, signal_5204}), .c ({signal_8673, signal_5361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5126 ( .a ({signal_12640, signal_12638}), .b ({signal_8521, signal_5205}), .c ({signal_8674, signal_5362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5127 ( .a ({signal_8268, signal_4820}), .b ({signal_8522, signal_5206}), .c ({signal_8675, signal_5363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5128 ( .a ({signal_8099, signal_4825}), .b ({signal_8371, signal_5088}), .c ({signal_8641, signal_5364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5129 ( .a ({signal_8101, signal_4827}), .b ({signal_8372, signal_5089}), .c ({signal_8642, signal_5365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5130 ( .a ({signal_8370, signal_5087}), .b ({signal_8475, signal_5210}), .c ({signal_8643, signal_5366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5131 ( .a ({signal_12644, signal_12642}), .b ({signal_8476, signal_5211}), .c ({signal_8644, signal_5367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5132 ( .a ({signal_8100, signal_4826}), .b ({signal_8477, signal_5212}), .c ({signal_8645, signal_5368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5133 ( .a ({signal_8105, signal_4831}), .b ({signal_8374, signal_5091}), .c ({signal_8646, signal_5369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5134 ( .a ({signal_8107, signal_4833}), .b ({signal_8375, signal_5092}), .c ({signal_8647, signal_5370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5135 ( .a ({signal_8373, signal_5090}), .b ({signal_8481, signal_5216}), .c ({signal_8648, signal_5371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5136 ( .a ({signal_12648, signal_12646}), .b ({signal_8482, signal_5217}), .c ({signal_8649, signal_5372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5137 ( .a ({signal_8106, signal_4832}), .b ({signal_8483, signal_5218}), .c ({signal_8650, signal_5373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5138 ( .a ({signal_8111, signal_4837}), .b ({signal_8377, signal_5094}), .c ({signal_8651, signal_5374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5139 ( .a ({signal_8113, signal_4839}), .b ({signal_8378, signal_5095}), .c ({signal_8652, signal_5375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5140 ( .a ({signal_8376, signal_5093}), .b ({signal_8487, signal_5222}), .c ({signal_8653, signal_5376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5141 ( .a ({signal_12652, signal_12650}), .b ({signal_8488, signal_5223}), .c ({signal_8654, signal_5377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5142 ( .a ({signal_8112, signal_4838}), .b ({signal_8489, signal_5224}), .c ({signal_8655, signal_5378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5143 ( .a ({signal_8117, signal_4843}), .b ({signal_8380, signal_5097}), .c ({signal_8656, signal_5379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5144 ( .a ({signal_8119, signal_4845}), .b ({signal_8381, signal_5098}), .c ({signal_8657, signal_5380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5145 ( .a ({signal_8379, signal_5096}), .b ({signal_8493, signal_5228}), .c ({signal_8658, signal_5381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5146 ( .a ({signal_12656, signal_12654}), .b ({signal_8494, signal_5229}), .c ({signal_8659, signal_5382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5147 ( .a ({signal_8118, signal_4844}), .b ({signal_8495, signal_5230}), .c ({signal_8660, signal_5383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5148 ( .a ({signal_8294, signal_5002}), .b ({signal_8525, signal_5233}), .c ({signal_8676, signal_5384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5149 ( .a ({signal_8296, signal_5004}), .b ({signal_8526, signal_5234}), .c ({signal_8677, signal_5385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5150 ( .a ({signal_8524, signal_5232}), .b ({signal_8565, signal_5273}), .c ({signal_8678, signal_5386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5151 ( .a ({signal_12660, signal_12658}), .b ({signal_8566, signal_5274}), .c ({signal_8679, signal_5387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5152 ( .a ({signal_8295, signal_5003}), .b ({signal_8567, signal_5275}), .c ({signal_8680, signal_5388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5153 ( .a ({signal_8300, signal_5008}), .b ({signal_8528, signal_5236}), .c ({signal_8681, signal_5389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5154 ( .a ({signal_8302, signal_5010}), .b ({signal_8529, signal_5237}), .c ({signal_8682, signal_5390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5155 ( .a ({signal_8527, signal_5235}), .b ({signal_8571, signal_5279}), .c ({signal_8683, signal_5391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5156 ( .a ({signal_12664, signal_12662}), .b ({signal_8572, signal_5280}), .c ({signal_8684, signal_5392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5157 ( .a ({signal_8301, signal_5009}), .b ({signal_8573, signal_5281}), .c ({signal_8685, signal_5393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5158 ( .a ({signal_8306, signal_5014}), .b ({signal_8531, signal_5239}), .c ({signal_8686, signal_5394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5159 ( .a ({signal_8308, signal_5016}), .b ({signal_8532, signal_5240}), .c ({signal_8687, signal_5395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5160 ( .a ({signal_8530, signal_5238}), .b ({signal_8577, signal_5285}), .c ({signal_8688, signal_5396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5161 ( .a ({signal_12668, signal_12666}), .b ({signal_8578, signal_5286}), .c ({signal_8689, signal_5397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5162 ( .a ({signal_8307, signal_5015}), .b ({signal_8579, signal_5287}), .c ({signal_8690, signal_5398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5163 ( .a ({signal_8312, signal_5020}), .b ({signal_8534, signal_5242}), .c ({signal_8691, signal_5399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5164 ( .a ({signal_8314, signal_5022}), .b ({signal_8535, signal_5243}), .c ({signal_8692, signal_5400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5165 ( .a ({signal_8533, signal_5241}), .b ({signal_8583, signal_5291}), .c ({signal_8693, signal_5401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5166 ( .a ({signal_12672, signal_12670}), .b ({signal_8584, signal_5292}), .c ({signal_8694, signal_5402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5167 ( .a ({signal_8313, signal_5021}), .b ({signal_8585, signal_5293}), .c ({signal_8695, signal_5403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5168 ( .a ({signal_8318, signal_5026}), .b ({signal_8537, signal_5245}), .c ({signal_8696, signal_5404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5169 ( .a ({signal_8320, signal_5028}), .b ({signal_8538, signal_5246}), .c ({signal_8697, signal_5405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5170 ( .a ({signal_8536, signal_5244}), .b ({signal_8589, signal_5297}), .c ({signal_8698, signal_5406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5171 ( .a ({signal_12676, signal_12674}), .b ({signal_8590, signal_5298}), .c ({signal_8699, signal_5407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5172 ( .a ({signal_8319, signal_5027}), .b ({signal_8591, signal_5299}), .c ({signal_8700, signal_5408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5173 ( .a ({signal_8324, signal_5032}), .b ({signal_8540, signal_5248}), .c ({signal_8701, signal_5409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5174 ( .a ({signal_8326, signal_5034}), .b ({signal_8541, signal_5249}), .c ({signal_8702, signal_5410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5175 ( .a ({signal_8539, signal_5247}), .b ({signal_8595, signal_5303}), .c ({signal_8703, signal_5411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5176 ( .a ({signal_12680, signal_12678}), .b ({signal_8596, signal_5304}), .c ({signal_8704, signal_5412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5177 ( .a ({signal_8325, signal_5033}), .b ({signal_8597, signal_5305}), .c ({signal_8705, signal_5413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5178 ( .a ({signal_8330, signal_5038}), .b ({signal_8543, signal_5251}), .c ({signal_8706, signal_5414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5179 ( .a ({signal_8332, signal_5040}), .b ({signal_8544, signal_5252}), .c ({signal_8707, signal_5415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5180 ( .a ({signal_8542, signal_5250}), .b ({signal_8601, signal_5309}), .c ({signal_8708, signal_5416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5181 ( .a ({signal_12684, signal_12682}), .b ({signal_8602, signal_5310}), .c ({signal_8709, signal_5417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5182 ( .a ({signal_8331, signal_5039}), .b ({signal_8603, signal_5311}), .c ({signal_8710, signal_5418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5183 ( .a ({signal_8661, signal_5313}), .b ({signal_8662, signal_5314}), .c ({signal_8757, signal_5419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5184 ( .a ({signal_8511, signal_5153}), .b ({signal_8663, signal_5315}), .c ({signal_8758, signal_5420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5185 ( .a ({signal_8662, signal_5314}), .b ({signal_8664, signal_5316}), .c ({signal_8759, signal_5421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5186 ( .a ({signal_8511, signal_5153}), .b ({signal_8665, signal_5317}), .c ({signal_8760, signal_5422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5187 ( .a ({signal_8336, signal_5047}), .b ({signal_8546, signal_5254}), .c ({signal_8711, signal_5423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5188 ( .a ({signal_8338, signal_5049}), .b ({signal_8547, signal_5255}), .c ({signal_8712, signal_5424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5189 ( .a ({signal_8545, signal_5253}), .b ({signal_8607, signal_5320}), .c ({signal_8713, signal_5425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5190 ( .a ({signal_12688, signal_12686}), .b ({signal_8608, signal_5321}), .c ({signal_8714, signal_5426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5191 ( .a ({signal_8337, signal_5048}), .b ({signal_8609, signal_5322}), .c ({signal_8715, signal_5427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5192 ( .a ({signal_8342, signal_5053}), .b ({signal_8549, signal_5257}), .c ({signal_8716, signal_5428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5193 ( .a ({signal_8344, signal_5055}), .b ({signal_8550, signal_5258}), .c ({signal_8717, signal_5429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5194 ( .a ({signal_8548, signal_5256}), .b ({signal_8613, signal_5326}), .c ({signal_8718, signal_5430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5195 ( .a ({signal_12692, signal_12690}), .b ({signal_8614, signal_5327}), .c ({signal_8719, signal_5431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5196 ( .a ({signal_8343, signal_5054}), .b ({signal_8615, signal_5328}), .c ({signal_8720, signal_5432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5197 ( .a ({signal_8348, signal_5059}), .b ({signal_8552, signal_5260}), .c ({signal_8721, signal_5433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5198 ( .a ({signal_8350, signal_5061}), .b ({signal_8553, signal_5261}), .c ({signal_8722, signal_5434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5199 ( .a ({signal_8551, signal_5259}), .b ({signal_8619, signal_5332}), .c ({signal_8723, signal_5435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5200 ( .a ({signal_12696, signal_12694}), .b ({signal_8620, signal_5333}), .c ({signal_8724, signal_5436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5201 ( .a ({signal_8349, signal_5060}), .b ({signal_8621, signal_5334}), .c ({signal_8725, signal_5437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5202 ( .a ({signal_8666, signal_5336}), .b ({signal_8667, signal_5337}), .c ({signal_8761, signal_5438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5203 ( .a ({signal_8517, signal_5180}), .b ({signal_8668, signal_5338}), .c ({signal_8762, signal_5439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5204 ( .a ({signal_8667, signal_5337}), .b ({signal_8669, signal_5339}), .c ({signal_8763, signal_5440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5205 ( .a ({signal_8517, signal_5180}), .b ({signal_8670, signal_5340}), .c ({signal_8764, signal_5441}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5206 ( .a ({signal_8354, signal_5068}), .b ({signal_8555, signal_5263}), .c ({signal_8726, signal_5442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5207 ( .a ({signal_8356, signal_5070}), .b ({signal_8556, signal_5264}), .c ({signal_8727, signal_5443}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5208 ( .a ({signal_8554, signal_5262}), .b ({signal_8625, signal_5343}), .c ({signal_8728, signal_5444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5209 ( .a ({signal_12700, signal_12698}), .b ({signal_8626, signal_5344}), .c ({signal_8729, signal_5445}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5210 ( .a ({signal_8355, signal_5069}), .b ({signal_8627, signal_5345}), .c ({signal_8730, signal_5446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5211 ( .a ({signal_8360, signal_5074}), .b ({signal_8558, signal_5266}), .c ({signal_8731, signal_5447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5212 ( .a ({signal_8362, signal_5076}), .b ({signal_8559, signal_5267}), .c ({signal_8732, signal_5448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5213 ( .a ({signal_8557, signal_5265}), .b ({signal_8631, signal_5349}), .c ({signal_8733, signal_5449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5214 ( .a ({signal_12704, signal_12702}), .b ({signal_8632, signal_5350}), .c ({signal_8734, signal_5450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5215 ( .a ({signal_8361, signal_5075}), .b ({signal_8633, signal_5351}), .c ({signal_8735, signal_5451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5216 ( .a ({signal_8366, signal_5080}), .b ({signal_8561, signal_5269}), .c ({signal_8736, signal_5452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5217 ( .a ({signal_8368, signal_5082}), .b ({signal_8562, signal_5270}), .c ({signal_8737, signal_5453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5218 ( .a ({signal_8560, signal_5268}), .b ({signal_8637, signal_5355}), .c ({signal_8738, signal_5454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5219 ( .a ({signal_12708, signal_12706}), .b ({signal_8638, signal_5356}), .c ({signal_8739, signal_5455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5220 ( .a ({signal_8367, signal_5081}), .b ({signal_8639, signal_5357}), .c ({signal_8740, signal_5456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5221 ( .a ({signal_8671, signal_5359}), .b ({signal_8672, signal_5360}), .c ({signal_8765, signal_5457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5222 ( .a ({signal_8523, signal_5207}), .b ({signal_8673, signal_5361}), .c ({signal_8766, signal_5458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5223 ( .a ({signal_8672, signal_5360}), .b ({signal_8674, signal_5362}), .c ({signal_8767, signal_5459}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5224 ( .a ({signal_8523, signal_5207}), .b ({signal_8675, signal_5363}), .c ({signal_8768, signal_5460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5225 ( .a ({signal_8641, signal_5364}), .b ({signal_8642, signal_5365}), .c ({signal_8741, signal_5461}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5226 ( .a ({signal_8478, signal_5213}), .b ({signal_8643, signal_5366}), .c ({signal_8742, signal_5462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5227 ( .a ({signal_8642, signal_5365}), .b ({signal_8644, signal_5367}), .c ({signal_8743, signal_5463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5228 ( .a ({signal_8478, signal_5213}), .b ({signal_8645, signal_5368}), .c ({signal_8744, signal_5464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5229 ( .a ({signal_8646, signal_5369}), .b ({signal_8647, signal_5370}), .c ({signal_8745, signal_5465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5230 ( .a ({signal_8484, signal_5219}), .b ({signal_8648, signal_5371}), .c ({signal_8746, signal_5466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5231 ( .a ({signal_8647, signal_5370}), .b ({signal_8649, signal_5372}), .c ({signal_8747, signal_5467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5232 ( .a ({signal_8484, signal_5219}), .b ({signal_8650, signal_5373}), .c ({signal_8748, signal_5468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5233 ( .a ({signal_8651, signal_5374}), .b ({signal_8652, signal_5375}), .c ({signal_8749, signal_5469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5234 ( .a ({signal_8490, signal_5225}), .b ({signal_8653, signal_5376}), .c ({signal_8750, signal_5470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5235 ( .a ({signal_8652, signal_5375}), .b ({signal_8654, signal_5377}), .c ({signal_8751, signal_5471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5236 ( .a ({signal_8490, signal_5225}), .b ({signal_8655, signal_5378}), .c ({signal_8752, signal_5472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5237 ( .a ({signal_8656, signal_5379}), .b ({signal_8657, signal_5380}), .c ({signal_8753, signal_5473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5238 ( .a ({signal_8496, signal_5231}), .b ({signal_8658, signal_5381}), .c ({signal_8754, signal_5474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5239 ( .a ({signal_8657, signal_5380}), .b ({signal_8659, signal_5382}), .c ({signal_8755, signal_5475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5240 ( .a ({signal_8496, signal_5231}), .b ({signal_8660, signal_5383}), .c ({signal_8756, signal_5476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5255 ( .a ({signal_8676, signal_5384}), .b ({signal_8677, signal_5385}), .c ({signal_8777, signal_5491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5256 ( .a ({signal_8568, signal_5276}), .b ({signal_8678, signal_5386}), .c ({signal_8778, signal_5492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5257 ( .a ({signal_8677, signal_5385}), .b ({signal_8679, signal_5387}), .c ({signal_8779, signal_5493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5258 ( .a ({signal_8568, signal_5276}), .b ({signal_8680, signal_5388}), .c ({signal_8780, signal_5494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5259 ( .a ({signal_8681, signal_5389}), .b ({signal_8682, signal_5390}), .c ({signal_8781, signal_5495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5260 ( .a ({signal_8574, signal_5282}), .b ({signal_8683, signal_5391}), .c ({signal_8782, signal_5496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5261 ( .a ({signal_8682, signal_5390}), .b ({signal_8684, signal_5392}), .c ({signal_8783, signal_5497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5262 ( .a ({signal_8574, signal_5282}), .b ({signal_8685, signal_5393}), .c ({signal_8784, signal_5498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5263 ( .a ({signal_8686, signal_5394}), .b ({signal_8687, signal_5395}), .c ({signal_8785, signal_5499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5264 ( .a ({signal_8580, signal_5288}), .b ({signal_8688, signal_5396}), .c ({signal_8786, signal_5500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5265 ( .a ({signal_8687, signal_5395}), .b ({signal_8689, signal_5397}), .c ({signal_8787, signal_5501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5266 ( .a ({signal_8580, signal_5288}), .b ({signal_8690, signal_5398}), .c ({signal_8788, signal_5502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5267 ( .a ({signal_8691, signal_5399}), .b ({signal_8692, signal_5400}), .c ({signal_8789, signal_5503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5268 ( .a ({signal_8586, signal_5294}), .b ({signal_8693, signal_5401}), .c ({signal_8790, signal_5504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5269 ( .a ({signal_8692, signal_5400}), .b ({signal_8694, signal_5402}), .c ({signal_8791, signal_5505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5270 ( .a ({signal_8586, signal_5294}), .b ({signal_8695, signal_5403}), .c ({signal_8792, signal_5506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5271 ( .a ({signal_8696, signal_5404}), .b ({signal_8697, signal_5405}), .c ({signal_8793, signal_5507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5272 ( .a ({signal_8592, signal_5300}), .b ({signal_8698, signal_5406}), .c ({signal_8794, signal_5508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5273 ( .a ({signal_8697, signal_5405}), .b ({signal_8699, signal_5407}), .c ({signal_8795, signal_5509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5274 ( .a ({signal_8592, signal_5300}), .b ({signal_8700, signal_5408}), .c ({signal_8796, signal_5510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5275 ( .a ({signal_8701, signal_5409}), .b ({signal_8702, signal_5410}), .c ({signal_8797, signal_5511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5276 ( .a ({signal_8598, signal_5306}), .b ({signal_8703, signal_5411}), .c ({signal_8798, signal_5512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5277 ( .a ({signal_8702, signal_5410}), .b ({signal_8704, signal_5412}), .c ({signal_8799, signal_5513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5278 ( .a ({signal_8598, signal_5306}), .b ({signal_8705, signal_5413}), .c ({signal_8800, signal_5514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5279 ( .a ({signal_8706, signal_5414}), .b ({signal_8707, signal_5415}), .c ({signal_8801, signal_5515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5280 ( .a ({signal_8604, signal_5312}), .b ({signal_8708, signal_5416}), .c ({signal_8802, signal_5516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5281 ( .a ({signal_8707, signal_5415}), .b ({signal_8709, signal_5417}), .c ({signal_8803, signal_5517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5282 ( .a ({signal_8604, signal_5312}), .b ({signal_8710, signal_5418}), .c ({signal_8804, signal_5518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5283 ( .a ({signal_12712, signal_12710}), .b ({signal_8757, signal_5419}), .c ({signal_8843, signal_5519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5284 ( .a ({signal_8758, signal_5420}), .b ({signal_8759, signal_5421}), .c ({signal_8844, signal_5520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5285 ( .a ({signal_8711, signal_5423}), .b ({signal_8712, signal_5424}), .c ({signal_8805, signal_5521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5286 ( .a ({signal_8610, signal_5323}), .b ({signal_8713, signal_5425}), .c ({signal_8806, signal_5522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5287 ( .a ({signal_8712, signal_5424}), .b ({signal_8714, signal_5426}), .c ({signal_8807, signal_5523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5288 ( .a ({signal_8610, signal_5323}), .b ({signal_8715, signal_5427}), .c ({signal_8808, signal_5524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5289 ( .a ({signal_8716, signal_5428}), .b ({signal_8717, signal_5429}), .c ({signal_8809, signal_5525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5290 ( .a ({signal_8616, signal_5329}), .b ({signal_8718, signal_5430}), .c ({signal_8810, signal_5526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5291 ( .a ({signal_8717, signal_5429}), .b ({signal_8719, signal_5431}), .c ({signal_8811, signal_5527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5292 ( .a ({signal_8616, signal_5329}), .b ({signal_8720, signal_5432}), .c ({signal_8812, signal_5528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5293 ( .a ({signal_8721, signal_5433}), .b ({signal_8722, signal_5434}), .c ({signal_8813, signal_5529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5294 ( .a ({signal_8622, signal_5335}), .b ({signal_8723, signal_5435}), .c ({signal_8814, signal_5530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5295 ( .a ({signal_8722, signal_5434}), .b ({signal_8724, signal_5436}), .c ({signal_8815, signal_5531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5296 ( .a ({signal_8622, signal_5335}), .b ({signal_8725, signal_5437}), .c ({signal_8816, signal_5532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5297 ( .a ({signal_12716, signal_12714}), .b ({signal_8761, signal_5438}), .c ({signal_8845, signal_5533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5298 ( .a ({signal_8762, signal_5439}), .b ({signal_8763, signal_5440}), .c ({signal_8846, signal_5534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5299 ( .a ({signal_8726, signal_5442}), .b ({signal_8727, signal_5443}), .c ({signal_8817, signal_5535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5300 ( .a ({signal_8628, signal_5346}), .b ({signal_8728, signal_5444}), .c ({signal_8818, signal_5536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5301 ( .a ({signal_8727, signal_5443}), .b ({signal_8729, signal_5445}), .c ({signal_8819, signal_5537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5302 ( .a ({signal_8628, signal_5346}), .b ({signal_8730, signal_5446}), .c ({signal_8820, signal_5538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5303 ( .a ({signal_8731, signal_5447}), .b ({signal_8732, signal_5448}), .c ({signal_8821, signal_5539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5304 ( .a ({signal_8634, signal_5352}), .b ({signal_8733, signal_5449}), .c ({signal_8822, signal_5540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5305 ( .a ({signal_8732, signal_5448}), .b ({signal_8734, signal_5450}), .c ({signal_8823, signal_5541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5306 ( .a ({signal_8634, signal_5352}), .b ({signal_8735, signal_5451}), .c ({signal_8824, signal_5542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5307 ( .a ({signal_8736, signal_5452}), .b ({signal_8737, signal_5453}), .c ({signal_8825, signal_5543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5308 ( .a ({signal_8640, signal_5358}), .b ({signal_8738, signal_5454}), .c ({signal_8826, signal_5544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5309 ( .a ({signal_8737, signal_5453}), .b ({signal_8739, signal_5455}), .c ({signal_8827, signal_5545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5310 ( .a ({signal_8640, signal_5358}), .b ({signal_8740, signal_5456}), .c ({signal_8828, signal_5546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5311 ( .a ({signal_12720, signal_12718}), .b ({signal_8765, signal_5457}), .c ({signal_8847, signal_5547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5312 ( .a ({signal_8766, signal_5458}), .b ({signal_8767, signal_5459}), .c ({signal_8848, signal_5548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5313 ( .a ({signal_12724, signal_12722}), .b ({signal_8741, signal_5461}), .c ({signal_8829, signal_5549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5314 ( .a ({signal_8742, signal_5462}), .b ({signal_8743, signal_5463}), .c ({signal_8830, signal_5550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5315 ( .a ({signal_12728, signal_12726}), .b ({signal_8745, signal_5465}), .c ({signal_8831, signal_5551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5316 ( .a ({signal_8746, signal_5466}), .b ({signal_8747, signal_5467}), .c ({signal_8832, signal_5552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5317 ( .a ({signal_12732, signal_12730}), .b ({signal_8749, signal_5469}), .c ({signal_8833, signal_5553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5318 ( .a ({signal_8750, signal_5470}), .b ({signal_8751, signal_5471}), .c ({signal_8834, signal_5554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5319 ( .a ({signal_12736, signal_12734}), .b ({signal_8753, signal_5473}), .c ({signal_8835, signal_5555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5320 ( .a ({signal_8754, signal_5474}), .b ({signal_8755, signal_5475}), .c ({signal_8836, signal_5556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5354 ( .a ({signal_12740, signal_12738}), .b ({signal_8777, signal_5491}), .c ({signal_8879, signal_5590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5355 ( .a ({signal_8778, signal_5492}), .b ({signal_8779, signal_5493}), .c ({signal_8880, signal_5591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5356 ( .a ({signal_12744, signal_12742}), .b ({signal_8781, signal_5495}), .c ({signal_8881, signal_5592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5357 ( .a ({signal_8782, signal_5496}), .b ({signal_8783, signal_5497}), .c ({signal_8882, signal_5593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5358 ( .a ({signal_12748, signal_12746}), .b ({signal_8785, signal_5499}), .c ({signal_8883, signal_5594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5359 ( .a ({signal_8786, signal_5500}), .b ({signal_8787, signal_5501}), .c ({signal_8884, signal_5595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5360 ( .a ({signal_12752, signal_12750}), .b ({signal_8789, signal_5503}), .c ({signal_8885, signal_5596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5361 ( .a ({signal_8790, signal_5504}), .b ({signal_8791, signal_5505}), .c ({signal_8886, signal_5597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5362 ( .a ({signal_12756, signal_12754}), .b ({signal_8793, signal_5507}), .c ({signal_8887, signal_5598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5363 ( .a ({signal_8794, signal_5508}), .b ({signal_8795, signal_5509}), .c ({signal_8888, signal_5599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5364 ( .a ({signal_12760, signal_12758}), .b ({signal_8797, signal_5511}), .c ({signal_8889, signal_5600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5365 ( .a ({signal_8798, signal_5512}), .b ({signal_8799, signal_5513}), .c ({signal_8890, signal_5601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5366 ( .a ({signal_12764, signal_12762}), .b ({signal_8801, signal_5515}), .c ({signal_8891, signal_5602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5367 ( .a ({signal_8802, signal_5516}), .b ({signal_8803, signal_5517}), .c ({signal_8892, signal_5603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5368 ( .a ({signal_8760, signal_5422}), .b ({signal_8843, signal_5519}), .c ({signal_8924, signal_5604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5372 ( .a ({signal_12768, signal_12766}), .b ({signal_8805, signal_5521}), .c ({signal_8893, signal_5608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5373 ( .a ({signal_8806, signal_5522}), .b ({signal_8807, signal_5523}), .c ({signal_8894, signal_5609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5374 ( .a ({signal_12772, signal_12770}), .b ({signal_8809, signal_5525}), .c ({signal_8895, signal_5610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5375 ( .a ({signal_8810, signal_5526}), .b ({signal_8811, signal_5527}), .c ({signal_8896, signal_5611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5376 ( .a ({signal_12776, signal_12774}), .b ({signal_8813, signal_5529}), .c ({signal_8897, signal_5612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5377 ( .a ({signal_8814, signal_5530}), .b ({signal_8815, signal_5531}), .c ({signal_8898, signal_5613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5378 ( .a ({signal_8764, signal_5441}), .b ({signal_8845, signal_5533}), .c ({signal_8928, signal_5614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5382 ( .a ({signal_12780, signal_12778}), .b ({signal_8817, signal_5535}), .c ({signal_8899, signal_5618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5383 ( .a ({signal_8818, signal_5536}), .b ({signal_8819, signal_5537}), .c ({signal_8900, signal_5619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5384 ( .a ({signal_12784, signal_12782}), .b ({signal_8821, signal_5539}), .c ({signal_8901, signal_5620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5385 ( .a ({signal_8822, signal_5540}), .b ({signal_8823, signal_5541}), .c ({signal_8902, signal_5621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5386 ( .a ({signal_12788, signal_12786}), .b ({signal_8825, signal_5543}), .c ({signal_8903, signal_5622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5387 ( .a ({signal_8826, signal_5544}), .b ({signal_8827, signal_5545}), .c ({signal_8904, signal_5623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5388 ( .a ({signal_8768, signal_5460}), .b ({signal_8847, signal_5547}), .c ({signal_8932, signal_5624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5392 ( .a ({signal_8744, signal_5464}), .b ({signal_8829, signal_5549}), .c ({signal_8905, signal_5628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5396 ( .a ({signal_8748, signal_5468}), .b ({signal_8831, signal_5551}), .c ({signal_8909, signal_5632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5400 ( .a ({signal_8752, signal_5472}), .b ({signal_8833, signal_5553}), .c ({signal_8913, signal_5636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5404 ( .a ({signal_8756, signal_5476}), .b ({signal_8835, signal_5555}), .c ({signal_8917, signal_5640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5449 ( .a ({signal_8780, signal_5494}), .b ({signal_8879, signal_5590}), .c ({signal_8965, signal_5685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5453 ( .a ({signal_8784, signal_5498}), .b ({signal_8881, signal_5592}), .c ({signal_8969, signal_5689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5457 ( .a ({signal_8788, signal_5502}), .b ({signal_8883, signal_5594}), .c ({signal_8973, signal_5693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5461 ( .a ({signal_8792, signal_5506}), .b ({signal_8885, signal_5596}), .c ({signal_8977, signal_5697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5465 ( .a ({signal_8796, signal_5510}), .b ({signal_8887, signal_5598}), .c ({signal_8981, signal_5701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5469 ( .a ({signal_8800, signal_5514}), .b ({signal_8889, signal_5600}), .c ({signal_8985, signal_5705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5473 ( .a ({signal_8804, signal_5518}), .b ({signal_8891, signal_5602}), .c ({signal_8989, signal_5709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5478 ( .a ({signal_8808, signal_5524}), .b ({signal_8893, signal_5608}), .c ({signal_8993, signal_5714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5482 ( .a ({signal_8812, signal_5528}), .b ({signal_8895, signal_5610}), .c ({signal_8997, signal_5718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5486 ( .a ({signal_8816, signal_5532}), .b ({signal_8897, signal_5612}), .c ({signal_9001, signal_5722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5491 ( .a ({signal_8820, signal_5538}), .b ({signal_8899, signal_5618}), .c ({signal_9005, signal_5727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5495 ( .a ({signal_8824, signal_5542}), .b ({signal_8901, signal_5620}), .c ({signal_9009, signal_5731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5499 ( .a ({signal_8828, signal_5546}), .b ({signal_8903, signal_5622}), .c ({signal_9013, signal_5735}) ) ;
    buf_clk cell_7582 ( .C (clk), .D (signal_12469), .Q (signal_12470) ) ;
    buf_clk cell_7584 ( .C (clk), .D (signal_12471), .Q (signal_12472) ) ;
    buf_clk cell_7586 ( .C (clk), .D (signal_12473), .Q (signal_12474) ) ;
    buf_clk cell_7588 ( .C (clk), .D (signal_12475), .Q (signal_12476) ) ;
    buf_clk cell_7590 ( .C (clk), .D (signal_12477), .Q (signal_12478) ) ;
    buf_clk cell_7592 ( .C (clk), .D (signal_12479), .Q (signal_12480) ) ;
    buf_clk cell_7594 ( .C (clk), .D (signal_12481), .Q (signal_12482) ) ;
    buf_clk cell_7596 ( .C (clk), .D (signal_12483), .Q (signal_12484) ) ;
    buf_clk cell_7598 ( .C (clk), .D (signal_12485), .Q (signal_12486) ) ;
    buf_clk cell_7600 ( .C (clk), .D (signal_12487), .Q (signal_12488) ) ;
    buf_clk cell_7602 ( .C (clk), .D (signal_12489), .Q (signal_12490) ) ;
    buf_clk cell_7604 ( .C (clk), .D (signal_12491), .Q (signal_12492) ) ;
    buf_clk cell_7606 ( .C (clk), .D (signal_12493), .Q (signal_12494) ) ;
    buf_clk cell_7608 ( .C (clk), .D (signal_12495), .Q (signal_12496) ) ;
    buf_clk cell_7610 ( .C (clk), .D (signal_12497), .Q (signal_12498) ) ;
    buf_clk cell_7612 ( .C (clk), .D (signal_12499), .Q (signal_12500) ) ;
    buf_clk cell_7614 ( .C (clk), .D (signal_12501), .Q (signal_12502) ) ;
    buf_clk cell_7616 ( .C (clk), .D (signal_12503), .Q (signal_12504) ) ;
    buf_clk cell_7618 ( .C (clk), .D (signal_12505), .Q (signal_12506) ) ;
    buf_clk cell_7620 ( .C (clk), .D (signal_12507), .Q (signal_12508) ) ;
    buf_clk cell_7622 ( .C (clk), .D (signal_12509), .Q (signal_12510) ) ;
    buf_clk cell_7624 ( .C (clk), .D (signal_12511), .Q (signal_12512) ) ;
    buf_clk cell_7626 ( .C (clk), .D (signal_12513), .Q (signal_12514) ) ;
    buf_clk cell_7628 ( .C (clk), .D (signal_12515), .Q (signal_12516) ) ;
    buf_clk cell_7630 ( .C (clk), .D (signal_12517), .Q (signal_12518) ) ;
    buf_clk cell_7632 ( .C (clk), .D (signal_12519), .Q (signal_12520) ) ;
    buf_clk cell_7634 ( .C (clk), .D (signal_12521), .Q (signal_12522) ) ;
    buf_clk cell_7636 ( .C (clk), .D (signal_12523), .Q (signal_12524) ) ;
    buf_clk cell_7638 ( .C (clk), .D (signal_12525), .Q (signal_12526) ) ;
    buf_clk cell_7640 ( .C (clk), .D (signal_12527), .Q (signal_12528) ) ;
    buf_clk cell_7642 ( .C (clk), .D (signal_12529), .Q (signal_12530) ) ;
    buf_clk cell_7644 ( .C (clk), .D (signal_12531), .Q (signal_12532) ) ;
    buf_clk cell_7646 ( .C (clk), .D (signal_12533), .Q (signal_12534) ) ;
    buf_clk cell_7648 ( .C (clk), .D (signal_12535), .Q (signal_12536) ) ;
    buf_clk cell_7650 ( .C (clk), .D (signal_12537), .Q (signal_12538) ) ;
    buf_clk cell_7652 ( .C (clk), .D (signal_12539), .Q (signal_12540) ) ;
    buf_clk cell_7654 ( .C (clk), .D (signal_12541), .Q (signal_12542) ) ;
    buf_clk cell_7656 ( .C (clk), .D (signal_12543), .Q (signal_12544) ) ;
    buf_clk cell_7658 ( .C (clk), .D (signal_12545), .Q (signal_12546) ) ;
    buf_clk cell_7660 ( .C (clk), .D (signal_12547), .Q (signal_12548) ) ;
    buf_clk cell_7662 ( .C (clk), .D (signal_12549), .Q (signal_12550) ) ;
    buf_clk cell_7664 ( .C (clk), .D (signal_12551), .Q (signal_12552) ) ;
    buf_clk cell_7666 ( .C (clk), .D (signal_12553), .Q (signal_12554) ) ;
    buf_clk cell_7668 ( .C (clk), .D (signal_12555), .Q (signal_12556) ) ;
    buf_clk cell_7670 ( .C (clk), .D (signal_12557), .Q (signal_12558) ) ;
    buf_clk cell_7672 ( .C (clk), .D (signal_12559), .Q (signal_12560) ) ;
    buf_clk cell_7674 ( .C (clk), .D (signal_12561), .Q (signal_12562) ) ;
    buf_clk cell_7676 ( .C (clk), .D (signal_12563), .Q (signal_12564) ) ;
    buf_clk cell_7678 ( .C (clk), .D (signal_12565), .Q (signal_12566) ) ;
    buf_clk cell_7680 ( .C (clk), .D (signal_12567), .Q (signal_12568) ) ;
    buf_clk cell_7682 ( .C (clk), .D (signal_12569), .Q (signal_12570) ) ;
    buf_clk cell_7684 ( .C (clk), .D (signal_12571), .Q (signal_12572) ) ;
    buf_clk cell_7686 ( .C (clk), .D (signal_12573), .Q (signal_12574) ) ;
    buf_clk cell_7688 ( .C (clk), .D (signal_12575), .Q (signal_12576) ) ;
    buf_clk cell_7690 ( .C (clk), .D (signal_12577), .Q (signal_12578) ) ;
    buf_clk cell_7692 ( .C (clk), .D (signal_12579), .Q (signal_12580) ) ;
    buf_clk cell_7694 ( .C (clk), .D (signal_12581), .Q (signal_12582) ) ;
    buf_clk cell_7696 ( .C (clk), .D (signal_12583), .Q (signal_12584) ) ;
    buf_clk cell_7698 ( .C (clk), .D (signal_12585), .Q (signal_12586) ) ;
    buf_clk cell_7700 ( .C (clk), .D (signal_12587), .Q (signal_12588) ) ;
    buf_clk cell_7702 ( .C (clk), .D (signal_12589), .Q (signal_12590) ) ;
    buf_clk cell_7704 ( .C (clk), .D (signal_12591), .Q (signal_12592) ) ;
    buf_clk cell_7706 ( .C (clk), .D (signal_12593), .Q (signal_12594) ) ;
    buf_clk cell_7708 ( .C (clk), .D (signal_12595), .Q (signal_12596) ) ;
    buf_clk cell_7710 ( .C (clk), .D (signal_12597), .Q (signal_12598) ) ;
    buf_clk cell_7712 ( .C (clk), .D (signal_12599), .Q (signal_12600) ) ;
    buf_clk cell_7714 ( .C (clk), .D (signal_12601), .Q (signal_12602) ) ;
    buf_clk cell_7716 ( .C (clk), .D (signal_12603), .Q (signal_12604) ) ;
    buf_clk cell_7718 ( .C (clk), .D (signal_12605), .Q (signal_12606) ) ;
    buf_clk cell_7720 ( .C (clk), .D (signal_12607), .Q (signal_12608) ) ;
    buf_clk cell_7722 ( .C (clk), .D (signal_12609), .Q (signal_12610) ) ;
    buf_clk cell_7724 ( .C (clk), .D (signal_12611), .Q (signal_12612) ) ;
    buf_clk cell_7726 ( .C (clk), .D (signal_12613), .Q (signal_12614) ) ;
    buf_clk cell_7728 ( .C (clk), .D (signal_12615), .Q (signal_12616) ) ;
    buf_clk cell_7730 ( .C (clk), .D (signal_12617), .Q (signal_12618) ) ;
    buf_clk cell_7732 ( .C (clk), .D (signal_12619), .Q (signal_12620) ) ;
    buf_clk cell_7734 ( .C (clk), .D (signal_12621), .Q (signal_12622) ) ;
    buf_clk cell_7736 ( .C (clk), .D (signal_12623), .Q (signal_12624) ) ;
    buf_clk cell_7738 ( .C (clk), .D (signal_12625), .Q (signal_12626) ) ;
    buf_clk cell_7740 ( .C (clk), .D (signal_12627), .Q (signal_12628) ) ;
    buf_clk cell_7742 ( .C (clk), .D (signal_12629), .Q (signal_12630) ) ;
    buf_clk cell_7744 ( .C (clk), .D (signal_12631), .Q (signal_12632) ) ;
    buf_clk cell_7746 ( .C (clk), .D (signal_12633), .Q (signal_12634) ) ;
    buf_clk cell_7748 ( .C (clk), .D (signal_12635), .Q (signal_12636) ) ;
    buf_clk cell_7750 ( .C (clk), .D (signal_12637), .Q (signal_12638) ) ;
    buf_clk cell_7752 ( .C (clk), .D (signal_12639), .Q (signal_12640) ) ;
    buf_clk cell_7754 ( .C (clk), .D (signal_12641), .Q (signal_12642) ) ;
    buf_clk cell_7756 ( .C (clk), .D (signal_12643), .Q (signal_12644) ) ;
    buf_clk cell_7758 ( .C (clk), .D (signal_12645), .Q (signal_12646) ) ;
    buf_clk cell_7760 ( .C (clk), .D (signal_12647), .Q (signal_12648) ) ;
    buf_clk cell_7762 ( .C (clk), .D (signal_12649), .Q (signal_12650) ) ;
    buf_clk cell_7764 ( .C (clk), .D (signal_12651), .Q (signal_12652) ) ;
    buf_clk cell_7766 ( .C (clk), .D (signal_12653), .Q (signal_12654) ) ;
    buf_clk cell_7768 ( .C (clk), .D (signal_12655), .Q (signal_12656) ) ;
    buf_clk cell_7770 ( .C (clk), .D (signal_12657), .Q (signal_12658) ) ;
    buf_clk cell_7772 ( .C (clk), .D (signal_12659), .Q (signal_12660) ) ;
    buf_clk cell_7774 ( .C (clk), .D (signal_12661), .Q (signal_12662) ) ;
    buf_clk cell_7776 ( .C (clk), .D (signal_12663), .Q (signal_12664) ) ;
    buf_clk cell_7778 ( .C (clk), .D (signal_12665), .Q (signal_12666) ) ;
    buf_clk cell_7780 ( .C (clk), .D (signal_12667), .Q (signal_12668) ) ;
    buf_clk cell_7782 ( .C (clk), .D (signal_12669), .Q (signal_12670) ) ;
    buf_clk cell_7784 ( .C (clk), .D (signal_12671), .Q (signal_12672) ) ;
    buf_clk cell_7786 ( .C (clk), .D (signal_12673), .Q (signal_12674) ) ;
    buf_clk cell_7788 ( .C (clk), .D (signal_12675), .Q (signal_12676) ) ;
    buf_clk cell_7790 ( .C (clk), .D (signal_12677), .Q (signal_12678) ) ;
    buf_clk cell_7792 ( .C (clk), .D (signal_12679), .Q (signal_12680) ) ;
    buf_clk cell_7794 ( .C (clk), .D (signal_12681), .Q (signal_12682) ) ;
    buf_clk cell_7796 ( .C (clk), .D (signal_12683), .Q (signal_12684) ) ;
    buf_clk cell_7798 ( .C (clk), .D (signal_12685), .Q (signal_12686) ) ;
    buf_clk cell_7800 ( .C (clk), .D (signal_12687), .Q (signal_12688) ) ;
    buf_clk cell_7802 ( .C (clk), .D (signal_12689), .Q (signal_12690) ) ;
    buf_clk cell_7804 ( .C (clk), .D (signal_12691), .Q (signal_12692) ) ;
    buf_clk cell_7806 ( .C (clk), .D (signal_12693), .Q (signal_12694) ) ;
    buf_clk cell_7808 ( .C (clk), .D (signal_12695), .Q (signal_12696) ) ;
    buf_clk cell_7810 ( .C (clk), .D (signal_12697), .Q (signal_12698) ) ;
    buf_clk cell_7812 ( .C (clk), .D (signal_12699), .Q (signal_12700) ) ;
    buf_clk cell_7814 ( .C (clk), .D (signal_12701), .Q (signal_12702) ) ;
    buf_clk cell_7816 ( .C (clk), .D (signal_12703), .Q (signal_12704) ) ;
    buf_clk cell_7818 ( .C (clk), .D (signal_12705), .Q (signal_12706) ) ;
    buf_clk cell_7820 ( .C (clk), .D (signal_12707), .Q (signal_12708) ) ;
    buf_clk cell_7822 ( .C (clk), .D (signal_12709), .Q (signal_12710) ) ;
    buf_clk cell_7824 ( .C (clk), .D (signal_12711), .Q (signal_12712) ) ;
    buf_clk cell_7826 ( .C (clk), .D (signal_12713), .Q (signal_12714) ) ;
    buf_clk cell_7828 ( .C (clk), .D (signal_12715), .Q (signal_12716) ) ;
    buf_clk cell_7830 ( .C (clk), .D (signal_12717), .Q (signal_12718) ) ;
    buf_clk cell_7832 ( .C (clk), .D (signal_12719), .Q (signal_12720) ) ;
    buf_clk cell_7834 ( .C (clk), .D (signal_12721), .Q (signal_12722) ) ;
    buf_clk cell_7836 ( .C (clk), .D (signal_12723), .Q (signal_12724) ) ;
    buf_clk cell_7838 ( .C (clk), .D (signal_12725), .Q (signal_12726) ) ;
    buf_clk cell_7840 ( .C (clk), .D (signal_12727), .Q (signal_12728) ) ;
    buf_clk cell_7842 ( .C (clk), .D (signal_12729), .Q (signal_12730) ) ;
    buf_clk cell_7844 ( .C (clk), .D (signal_12731), .Q (signal_12732) ) ;
    buf_clk cell_7846 ( .C (clk), .D (signal_12733), .Q (signal_12734) ) ;
    buf_clk cell_7848 ( .C (clk), .D (signal_12735), .Q (signal_12736) ) ;
    buf_clk cell_7850 ( .C (clk), .D (signal_12737), .Q (signal_12738) ) ;
    buf_clk cell_7852 ( .C (clk), .D (signal_12739), .Q (signal_12740) ) ;
    buf_clk cell_7854 ( .C (clk), .D (signal_12741), .Q (signal_12742) ) ;
    buf_clk cell_7856 ( .C (clk), .D (signal_12743), .Q (signal_12744) ) ;
    buf_clk cell_7858 ( .C (clk), .D (signal_12745), .Q (signal_12746) ) ;
    buf_clk cell_7860 ( .C (clk), .D (signal_12747), .Q (signal_12748) ) ;
    buf_clk cell_7862 ( .C (clk), .D (signal_12749), .Q (signal_12750) ) ;
    buf_clk cell_7864 ( .C (clk), .D (signal_12751), .Q (signal_12752) ) ;
    buf_clk cell_7866 ( .C (clk), .D (signal_12753), .Q (signal_12754) ) ;
    buf_clk cell_7868 ( .C (clk), .D (signal_12755), .Q (signal_12756) ) ;
    buf_clk cell_7870 ( .C (clk), .D (signal_12757), .Q (signal_12758) ) ;
    buf_clk cell_7872 ( .C (clk), .D (signal_12759), .Q (signal_12760) ) ;
    buf_clk cell_7874 ( .C (clk), .D (signal_12761), .Q (signal_12762) ) ;
    buf_clk cell_7876 ( .C (clk), .D (signal_12763), .Q (signal_12764) ) ;
    buf_clk cell_7878 ( .C (clk), .D (signal_12765), .Q (signal_12766) ) ;
    buf_clk cell_7880 ( .C (clk), .D (signal_12767), .Q (signal_12768) ) ;
    buf_clk cell_7882 ( .C (clk), .D (signal_12769), .Q (signal_12770) ) ;
    buf_clk cell_7884 ( .C (clk), .D (signal_12771), .Q (signal_12772) ) ;
    buf_clk cell_7886 ( .C (clk), .D (signal_12773), .Q (signal_12774) ) ;
    buf_clk cell_7888 ( .C (clk), .D (signal_12775), .Q (signal_12776) ) ;
    buf_clk cell_7890 ( .C (clk), .D (signal_12777), .Q (signal_12778) ) ;
    buf_clk cell_7892 ( .C (clk), .D (signal_12779), .Q (signal_12780) ) ;
    buf_clk cell_7894 ( .C (clk), .D (signal_12781), .Q (signal_12782) ) ;
    buf_clk cell_7896 ( .C (clk), .D (signal_12783), .Q (signal_12784) ) ;
    buf_clk cell_7898 ( .C (clk), .D (signal_12785), .Q (signal_12786) ) ;
    buf_clk cell_7900 ( .C (clk), .D (signal_12787), .Q (signal_12788) ) ;
    buf_clk cell_8542 ( .C (clk), .D (signal_13429), .Q (signal_13430) ) ;
    buf_clk cell_8550 ( .C (clk), .D (signal_13437), .Q (signal_13438) ) ;
    buf_clk cell_8558 ( .C (clk), .D (signal_13445), .Q (signal_13446) ) ;
    buf_clk cell_8566 ( .C (clk), .D (signal_13453), .Q (signal_13454) ) ;
    buf_clk cell_8574 ( .C (clk), .D (signal_13461), .Q (signal_13462) ) ;
    buf_clk cell_8582 ( .C (clk), .D (signal_13469), .Q (signal_13470) ) ;
    buf_clk cell_8590 ( .C (clk), .D (signal_13477), .Q (signal_13478) ) ;
    buf_clk cell_8598 ( .C (clk), .D (signal_13485), .Q (signal_13486) ) ;
    buf_clk cell_8606 ( .C (clk), .D (signal_13493), .Q (signal_13494) ) ;
    buf_clk cell_8614 ( .C (clk), .D (signal_13501), .Q (signal_13502) ) ;
    buf_clk cell_8622 ( .C (clk), .D (signal_13509), .Q (signal_13510) ) ;
    buf_clk cell_8630 ( .C (clk), .D (signal_13517), .Q (signal_13518) ) ;
    buf_clk cell_8638 ( .C (clk), .D (signal_13525), .Q (signal_13526) ) ;
    buf_clk cell_8646 ( .C (clk), .D (signal_13533), .Q (signal_13534) ) ;
    buf_clk cell_8654 ( .C (clk), .D (signal_13541), .Q (signal_13542) ) ;
    buf_clk cell_8662 ( .C (clk), .D (signal_13549), .Q (signal_13550) ) ;
    buf_clk cell_8670 ( .C (clk), .D (signal_13557), .Q (signal_13558) ) ;
    buf_clk cell_8678 ( .C (clk), .D (signal_13565), .Q (signal_13566) ) ;
    buf_clk cell_8686 ( .C (clk), .D (signal_13573), .Q (signal_13574) ) ;
    buf_clk cell_8694 ( .C (clk), .D (signal_13581), .Q (signal_13582) ) ;
    buf_clk cell_8702 ( .C (clk), .D (signal_13589), .Q (signal_13590) ) ;
    buf_clk cell_8710 ( .C (clk), .D (signal_13597), .Q (signal_13598) ) ;
    buf_clk cell_8718 ( .C (clk), .D (signal_13605), .Q (signal_13606) ) ;
    buf_clk cell_8726 ( .C (clk), .D (signal_13613), .Q (signal_13614) ) ;
    buf_clk cell_8734 ( .C (clk), .D (signal_13621), .Q (signal_13622) ) ;
    buf_clk cell_8742 ( .C (clk), .D (signal_13629), .Q (signal_13630) ) ;
    buf_clk cell_8750 ( .C (clk), .D (signal_13637), .Q (signal_13638) ) ;
    buf_clk cell_8758 ( .C (clk), .D (signal_13645), .Q (signal_13646) ) ;
    buf_clk cell_8766 ( .C (clk), .D (signal_13653), .Q (signal_13654) ) ;
    buf_clk cell_8774 ( .C (clk), .D (signal_13661), .Q (signal_13662) ) ;
    buf_clk cell_8782 ( .C (clk), .D (signal_13669), .Q (signal_13670) ) ;
    buf_clk cell_8790 ( .C (clk), .D (signal_13677), .Q (signal_13678) ) ;
    buf_clk cell_8798 ( .C (clk), .D (signal_13685), .Q (signal_13686) ) ;
    buf_clk cell_8806 ( .C (clk), .D (signal_13693), .Q (signal_13694) ) ;
    buf_clk cell_8814 ( .C (clk), .D (signal_13701), .Q (signal_13702) ) ;
    buf_clk cell_8822 ( .C (clk), .D (signal_13709), .Q (signal_13710) ) ;
    buf_clk cell_8830 ( .C (clk), .D (signal_13717), .Q (signal_13718) ) ;
    buf_clk cell_8838 ( .C (clk), .D (signal_13725), .Q (signal_13726) ) ;
    buf_clk cell_8846 ( .C (clk), .D (signal_13733), .Q (signal_13734) ) ;
    buf_clk cell_8854 ( .C (clk), .D (signal_13741), .Q (signal_13742) ) ;
    buf_clk cell_8862 ( .C (clk), .D (signal_13749), .Q (signal_13750) ) ;
    buf_clk cell_8870 ( .C (clk), .D (signal_13757), .Q (signal_13758) ) ;
    buf_clk cell_8878 ( .C (clk), .D (signal_13765), .Q (signal_13766) ) ;
    buf_clk cell_8886 ( .C (clk), .D (signal_13773), .Q (signal_13774) ) ;
    buf_clk cell_8894 ( .C (clk), .D (signal_13781), .Q (signal_13782) ) ;
    buf_clk cell_8902 ( .C (clk), .D (signal_13789), .Q (signal_13790) ) ;
    buf_clk cell_8910 ( .C (clk), .D (signal_13797), .Q (signal_13798) ) ;
    buf_clk cell_8918 ( .C (clk), .D (signal_13805), .Q (signal_13806) ) ;
    buf_clk cell_8926 ( .C (clk), .D (signal_13813), .Q (signal_13814) ) ;
    buf_clk cell_8934 ( .C (clk), .D (signal_13821), .Q (signal_13822) ) ;
    buf_clk cell_8942 ( .C (clk), .D (signal_13829), .Q (signal_13830) ) ;
    buf_clk cell_8950 ( .C (clk), .D (signal_13837), .Q (signal_13838) ) ;
    buf_clk cell_8958 ( .C (clk), .D (signal_13845), .Q (signal_13846) ) ;
    buf_clk cell_8966 ( .C (clk), .D (signal_13853), .Q (signal_13854) ) ;
    buf_clk cell_8974 ( .C (clk), .D (signal_13861), .Q (signal_13862) ) ;
    buf_clk cell_8982 ( .C (clk), .D (signal_13869), .Q (signal_13870) ) ;
    buf_clk cell_8990 ( .C (clk), .D (signal_13877), .Q (signal_13878) ) ;
    buf_clk cell_8998 ( .C (clk), .D (signal_13885), .Q (signal_13886) ) ;
    buf_clk cell_9006 ( .C (clk), .D (signal_13893), .Q (signal_13894) ) ;
    buf_clk cell_9014 ( .C (clk), .D (signal_13901), .Q (signal_13902) ) ;
    buf_clk cell_9022 ( .C (clk), .D (signal_13909), .Q (signal_13910) ) ;
    buf_clk cell_9030 ( .C (clk), .D (signal_13917), .Q (signal_13918) ) ;
    buf_clk cell_9038 ( .C (clk), .D (signal_13925), .Q (signal_13926) ) ;
    buf_clk cell_9046 ( .C (clk), .D (signal_13933), .Q (signal_13934) ) ;
    buf_clk cell_9054 ( .C (clk), .D (signal_13941), .Q (signal_13942) ) ;
    buf_clk cell_9062 ( .C (clk), .D (signal_13949), .Q (signal_13950) ) ;
    buf_clk cell_9070 ( .C (clk), .D (signal_13957), .Q (signal_13958) ) ;
    buf_clk cell_9078 ( .C (clk), .D (signal_13965), .Q (signal_13966) ) ;
    buf_clk cell_9086 ( .C (clk), .D (signal_13973), .Q (signal_13974) ) ;
    buf_clk cell_9094 ( .C (clk), .D (signal_13981), .Q (signal_13982) ) ;
    buf_clk cell_9102 ( .C (clk), .D (signal_13989), .Q (signal_13990) ) ;
    buf_clk cell_9110 ( .C (clk), .D (signal_13997), .Q (signal_13998) ) ;
    buf_clk cell_9118 ( .C (clk), .D (signal_14005), .Q (signal_14006) ) ;
    buf_clk cell_9126 ( .C (clk), .D (signal_14013), .Q (signal_14014) ) ;
    buf_clk cell_9134 ( .C (clk), .D (signal_14021), .Q (signal_14022) ) ;
    buf_clk cell_9142 ( .C (clk), .D (signal_14029), .Q (signal_14030) ) ;
    buf_clk cell_9150 ( .C (clk), .D (signal_14037), .Q (signal_14038) ) ;
    buf_clk cell_9158 ( .C (clk), .D (signal_14045), .Q (signal_14046) ) ;
    buf_clk cell_9166 ( .C (clk), .D (signal_14053), .Q (signal_14054) ) ;
    buf_clk cell_9174 ( .C (clk), .D (signal_14061), .Q (signal_14062) ) ;
    buf_clk cell_9182 ( .C (clk), .D (signal_14069), .Q (signal_14070) ) ;
    buf_clk cell_9190 ( .C (clk), .D (signal_14077), .Q (signal_14078) ) ;
    buf_clk cell_9198 ( .C (clk), .D (signal_14085), .Q (signal_14086) ) ;
    buf_clk cell_9206 ( .C (clk), .D (signal_14093), .Q (signal_14094) ) ;
    buf_clk cell_9214 ( .C (clk), .D (signal_14101), .Q (signal_14102) ) ;
    buf_clk cell_9222 ( .C (clk), .D (signal_14109), .Q (signal_14110) ) ;
    buf_clk cell_9230 ( .C (clk), .D (signal_14117), .Q (signal_14118) ) ;
    buf_clk cell_9238 ( .C (clk), .D (signal_14125), .Q (signal_14126) ) ;
    buf_clk cell_9246 ( .C (clk), .D (signal_14133), .Q (signal_14134) ) ;
    buf_clk cell_9254 ( .C (clk), .D (signal_14141), .Q (signal_14142) ) ;
    buf_clk cell_9262 ( .C (clk), .D (signal_14149), .Q (signal_14150) ) ;
    buf_clk cell_9270 ( .C (clk), .D (signal_14157), .Q (signal_14158) ) ;
    buf_clk cell_9278 ( .C (clk), .D (signal_14165), .Q (signal_14166) ) ;
    buf_clk cell_9286 ( .C (clk), .D (signal_14173), .Q (signal_14174) ) ;
    buf_clk cell_9294 ( .C (clk), .D (signal_14181), .Q (signal_14182) ) ;
    buf_clk cell_9302 ( .C (clk), .D (signal_14189), .Q (signal_14190) ) ;
    buf_clk cell_9310 ( .C (clk), .D (signal_14197), .Q (signal_14198) ) ;
    buf_clk cell_9318 ( .C (clk), .D (signal_14205), .Q (signal_14206) ) ;
    buf_clk cell_9326 ( .C (clk), .D (signal_14213), .Q (signal_14214) ) ;
    buf_clk cell_9334 ( .C (clk), .D (signal_14221), .Q (signal_14222) ) ;
    buf_clk cell_9342 ( .C (clk), .D (signal_14229), .Q (signal_14230) ) ;
    buf_clk cell_9350 ( .C (clk), .D (signal_14237), .Q (signal_14238) ) ;
    buf_clk cell_9358 ( .C (clk), .D (signal_14245), .Q (signal_14246) ) ;
    buf_clk cell_9366 ( .C (clk), .D (signal_14253), .Q (signal_14254) ) ;
    buf_clk cell_9374 ( .C (clk), .D (signal_14261), .Q (signal_14262) ) ;
    buf_clk cell_9382 ( .C (clk), .D (signal_14269), .Q (signal_14270) ) ;
    buf_clk cell_9390 ( .C (clk), .D (signal_14277), .Q (signal_14278) ) ;
    buf_clk cell_9398 ( .C (clk), .D (signal_14285), .Q (signal_14286) ) ;
    buf_clk cell_9406 ( .C (clk), .D (signal_14293), .Q (signal_14294) ) ;
    buf_clk cell_9414 ( .C (clk), .D (signal_14301), .Q (signal_14302) ) ;
    buf_clk cell_9422 ( .C (clk), .D (signal_14309), .Q (signal_14310) ) ;
    buf_clk cell_9430 ( .C (clk), .D (signal_14317), .Q (signal_14318) ) ;
    buf_clk cell_9438 ( .C (clk), .D (signal_14325), .Q (signal_14326) ) ;
    buf_clk cell_9446 ( .C (clk), .D (signal_14333), .Q (signal_14334) ) ;
    buf_clk cell_9454 ( .C (clk), .D (signal_14341), .Q (signal_14342) ) ;
    buf_clk cell_9462 ( .C (clk), .D (signal_14349), .Q (signal_14350) ) ;
    buf_clk cell_9470 ( .C (clk), .D (signal_14357), .Q (signal_14358) ) ;
    buf_clk cell_9478 ( .C (clk), .D (signal_14365), .Q (signal_14366) ) ;
    buf_clk cell_9486 ( .C (clk), .D (signal_14373), .Q (signal_14374) ) ;
    buf_clk cell_9494 ( .C (clk), .D (signal_14381), .Q (signal_14382) ) ;
    buf_clk cell_9502 ( .C (clk), .D (signal_14389), .Q (signal_14390) ) ;
    buf_clk cell_9510 ( .C (clk), .D (signal_14397), .Q (signal_14398) ) ;
    buf_clk cell_9518 ( .C (clk), .D (signal_14405), .Q (signal_14406) ) ;
    buf_clk cell_9526 ( .C (clk), .D (signal_14413), .Q (signal_14414) ) ;
    buf_clk cell_9534 ( .C (clk), .D (signal_14421), .Q (signal_14422) ) ;
    buf_clk cell_9542 ( .C (clk), .D (signal_14429), .Q (signal_14430) ) ;
    buf_clk cell_9550 ( .C (clk), .D (signal_14437), .Q (signal_14438) ) ;
    buf_clk cell_9558 ( .C (clk), .D (signal_14445), .Q (signal_14446) ) ;
    buf_clk cell_9566 ( .C (clk), .D (signal_14453), .Q (signal_14454) ) ;
    buf_clk cell_9574 ( .C (clk), .D (signal_14461), .Q (signal_14462) ) ;
    buf_clk cell_9582 ( .C (clk), .D (signal_14469), .Q (signal_14470) ) ;
    buf_clk cell_9590 ( .C (clk), .D (signal_14477), .Q (signal_14478) ) ;
    buf_clk cell_9598 ( .C (clk), .D (signal_14485), .Q (signal_14486) ) ;
    buf_clk cell_9606 ( .C (clk), .D (signal_14493), .Q (signal_14494) ) ;
    buf_clk cell_9614 ( .C (clk), .D (signal_14501), .Q (signal_14502) ) ;
    buf_clk cell_9622 ( .C (clk), .D (signal_14509), .Q (signal_14510) ) ;
    buf_clk cell_9630 ( .C (clk), .D (signal_14517), .Q (signal_14518) ) ;
    buf_clk cell_9638 ( .C (clk), .D (signal_14525), .Q (signal_14526) ) ;
    buf_clk cell_9646 ( .C (clk), .D (signal_14533), .Q (signal_14534) ) ;
    buf_clk cell_9654 ( .C (clk), .D (signal_14541), .Q (signal_14542) ) ;
    buf_clk cell_9662 ( .C (clk), .D (signal_14549), .Q (signal_14550) ) ;
    buf_clk cell_9670 ( .C (clk), .D (signal_14557), .Q (signal_14558) ) ;
    buf_clk cell_9678 ( .C (clk), .D (signal_14565), .Q (signal_14566) ) ;
    buf_clk cell_9686 ( .C (clk), .D (signal_14573), .Q (signal_14574) ) ;
    buf_clk cell_9694 ( .C (clk), .D (signal_14581), .Q (signal_14582) ) ;
    buf_clk cell_9702 ( .C (clk), .D (signal_14589), .Q (signal_14590) ) ;
    buf_clk cell_9710 ( .C (clk), .D (signal_14597), .Q (signal_14598) ) ;
    buf_clk cell_9718 ( .C (clk), .D (signal_14605), .Q (signal_14606) ) ;
    buf_clk cell_9726 ( .C (clk), .D (signal_14613), .Q (signal_14614) ) ;
    buf_clk cell_9734 ( .C (clk), .D (signal_14621), .Q (signal_14622) ) ;
    buf_clk cell_9742 ( .C (clk), .D (signal_14629), .Q (signal_14630) ) ;
    buf_clk cell_9750 ( .C (clk), .D (signal_14637), .Q (signal_14638) ) ;
    buf_clk cell_9758 ( .C (clk), .D (signal_14645), .Q (signal_14646) ) ;
    buf_clk cell_9766 ( .C (clk), .D (signal_14653), .Q (signal_14654) ) ;
    buf_clk cell_9774 ( .C (clk), .D (signal_14661), .Q (signal_14662) ) ;
    buf_clk cell_9782 ( .C (clk), .D (signal_14669), .Q (signal_14670) ) ;
    buf_clk cell_9790 ( .C (clk), .D (signal_14677), .Q (signal_14678) ) ;
    buf_clk cell_9798 ( .C (clk), .D (signal_14685), .Q (signal_14686) ) ;
    buf_clk cell_9806 ( .C (clk), .D (signal_14693), .Q (signal_14694) ) ;
    buf_clk cell_9814 ( .C (clk), .D (signal_14701), .Q (signal_14702) ) ;
    buf_clk cell_9822 ( .C (clk), .D (signal_14709), .Q (signal_14710) ) ;
    buf_clk cell_9830 ( .C (clk), .D (signal_14717), .Q (signal_14718) ) ;
    buf_clk cell_9838 ( .C (clk), .D (signal_14725), .Q (signal_14726) ) ;
    buf_clk cell_9846 ( .C (clk), .D (signal_14733), .Q (signal_14734) ) ;
    buf_clk cell_9854 ( .C (clk), .D (signal_14741), .Q (signal_14742) ) ;
    buf_clk cell_9862 ( .C (clk), .D (signal_14749), .Q (signal_14750) ) ;
    buf_clk cell_9870 ( .C (clk), .D (signal_14757), .Q (signal_14758) ) ;
    buf_clk cell_9878 ( .C (clk), .D (signal_14765), .Q (signal_14766) ) ;
    buf_clk cell_9886 ( .C (clk), .D (signal_14773), .Q (signal_14774) ) ;
    buf_clk cell_9894 ( .C (clk), .D (signal_14781), .Q (signal_14782) ) ;
    buf_clk cell_9902 ( .C (clk), .D (signal_14789), .Q (signal_14790) ) ;
    buf_clk cell_9910 ( .C (clk), .D (signal_14797), .Q (signal_14798) ) ;
    buf_clk cell_9918 ( .C (clk), .D (signal_14805), .Q (signal_14806) ) ;
    buf_clk cell_9926 ( .C (clk), .D (signal_14813), .Q (signal_14814) ) ;
    buf_clk cell_9934 ( .C (clk), .D (signal_14821), .Q (signal_14822) ) ;
    buf_clk cell_9942 ( .C (clk), .D (signal_14829), .Q (signal_14830) ) ;
    buf_clk cell_9950 ( .C (clk), .D (signal_14837), .Q (signal_14838) ) ;
    buf_clk cell_9958 ( .C (clk), .D (signal_14845), .Q (signal_14846) ) ;
    buf_clk cell_9966 ( .C (clk), .D (signal_14853), .Q (signal_14854) ) ;
    buf_clk cell_9974 ( .C (clk), .D (signal_14861), .Q (signal_14862) ) ;
    buf_clk cell_9982 ( .C (clk), .D (signal_14869), .Q (signal_14870) ) ;
    buf_clk cell_9990 ( .C (clk), .D (signal_14877), .Q (signal_14878) ) ;
    buf_clk cell_9998 ( .C (clk), .D (signal_14885), .Q (signal_14886) ) ;
    buf_clk cell_10006 ( .C (clk), .D (signal_14893), .Q (signal_14894) ) ;
    buf_clk cell_10014 ( .C (clk), .D (signal_14901), .Q (signal_14902) ) ;
    buf_clk cell_10022 ( .C (clk), .D (signal_14909), .Q (signal_14910) ) ;
    buf_clk cell_10030 ( .C (clk), .D (signal_14917), .Q (signal_14918) ) ;
    buf_clk cell_10038 ( .C (clk), .D (signal_14925), .Q (signal_14926) ) ;
    buf_clk cell_10046 ( .C (clk), .D (signal_14933), .Q (signal_14934) ) ;
    buf_clk cell_10054 ( .C (clk), .D (signal_14941), .Q (signal_14942) ) ;
    buf_clk cell_10062 ( .C (clk), .D (signal_14949), .Q (signal_14950) ) ;
    buf_clk cell_10070 ( .C (clk), .D (signal_14957), .Q (signal_14958) ) ;
    buf_clk cell_10078 ( .C (clk), .D (signal_14965), .Q (signal_14966) ) ;
    buf_clk cell_10086 ( .C (clk), .D (signal_14973), .Q (signal_14974) ) ;
    buf_clk cell_10094 ( .C (clk), .D (signal_14981), .Q (signal_14982) ) ;
    buf_clk cell_10102 ( .C (clk), .D (signal_14989), .Q (signal_14990) ) ;
    buf_clk cell_10110 ( .C (clk), .D (signal_14997), .Q (signal_14998) ) ;
    buf_clk cell_10118 ( .C (clk), .D (signal_15005), .Q (signal_15006) ) ;
    buf_clk cell_10126 ( .C (clk), .D (signal_15013), .Q (signal_15014) ) ;
    buf_clk cell_10134 ( .C (clk), .D (signal_15021), .Q (signal_15022) ) ;
    buf_clk cell_10142 ( .C (clk), .D (signal_15029), .Q (signal_15030) ) ;
    buf_clk cell_10150 ( .C (clk), .D (signal_15037), .Q (signal_15038) ) ;
    buf_clk cell_10158 ( .C (clk), .D (signal_15045), .Q (signal_15046) ) ;
    buf_clk cell_10166 ( .C (clk), .D (signal_15053), .Q (signal_15054) ) ;
    buf_clk cell_10174 ( .C (clk), .D (signal_15061), .Q (signal_15062) ) ;
    buf_clk cell_10182 ( .C (clk), .D (signal_15069), .Q (signal_15070) ) ;
    buf_clk cell_10190 ( .C (clk), .D (signal_15077), .Q (signal_15078) ) ;
    buf_clk cell_10198 ( .C (clk), .D (signal_15085), .Q (signal_15086) ) ;
    buf_clk cell_10206 ( .C (clk), .D (signal_15093), .Q (signal_15094) ) ;
    buf_clk cell_10214 ( .C (clk), .D (signal_15101), .Q (signal_15102) ) ;
    buf_clk cell_10222 ( .C (clk), .D (signal_15109), .Q (signal_15110) ) ;
    buf_clk cell_10230 ( .C (clk), .D (signal_15117), .Q (signal_15118) ) ;
    buf_clk cell_10238 ( .C (clk), .D (signal_15125), .Q (signal_15126) ) ;
    buf_clk cell_10246 ( .C (clk), .D (signal_15133), .Q (signal_15134) ) ;
    buf_clk cell_10254 ( .C (clk), .D (signal_15141), .Q (signal_15142) ) ;
    buf_clk cell_10262 ( .C (clk), .D (signal_15149), .Q (signal_15150) ) ;
    buf_clk cell_10270 ( .C (clk), .D (signal_15157), .Q (signal_15158) ) ;
    buf_clk cell_10278 ( .C (clk), .D (signal_15165), .Q (signal_15166) ) ;
    buf_clk cell_10286 ( .C (clk), .D (signal_15173), .Q (signal_15174) ) ;
    buf_clk cell_10294 ( .C (clk), .D (signal_15181), .Q (signal_15182) ) ;
    buf_clk cell_10302 ( .C (clk), .D (signal_15189), .Q (signal_15190) ) ;
    buf_clk cell_10310 ( .C (clk), .D (signal_15197), .Q (signal_15198) ) ;
    buf_clk cell_10318 ( .C (clk), .D (signal_15205), .Q (signal_15206) ) ;
    buf_clk cell_10326 ( .C (clk), .D (signal_15213), .Q (signal_15214) ) ;
    buf_clk cell_10334 ( .C (clk), .D (signal_15221), .Q (signal_15222) ) ;
    buf_clk cell_10342 ( .C (clk), .D (signal_15229), .Q (signal_15230) ) ;
    buf_clk cell_10350 ( .C (clk), .D (signal_15237), .Q (signal_15238) ) ;
    buf_clk cell_10358 ( .C (clk), .D (signal_15245), .Q (signal_15246) ) ;
    buf_clk cell_10366 ( .C (clk), .D (signal_15253), .Q (signal_15254) ) ;
    buf_clk cell_10374 ( .C (clk), .D (signal_15261), .Q (signal_15262) ) ;
    buf_clk cell_10382 ( .C (clk), .D (signal_15269), .Q (signal_15270) ) ;
    buf_clk cell_10390 ( .C (clk), .D (signal_15277), .Q (signal_15278) ) ;
    buf_clk cell_10398 ( .C (clk), .D (signal_15285), .Q (signal_15286) ) ;
    buf_clk cell_10406 ( .C (clk), .D (signal_15293), .Q (signal_15294) ) ;
    buf_clk cell_10414 ( .C (clk), .D (signal_15301), .Q (signal_15302) ) ;
    buf_clk cell_10422 ( .C (clk), .D (signal_15309), .Q (signal_15310) ) ;
    buf_clk cell_10430 ( .C (clk), .D (signal_15317), .Q (signal_15318) ) ;
    buf_clk cell_10438 ( .C (clk), .D (signal_15325), .Q (signal_15326) ) ;
    buf_clk cell_10446 ( .C (clk), .D (signal_15333), .Q (signal_15334) ) ;
    buf_clk cell_10454 ( .C (clk), .D (signal_15341), .Q (signal_15342) ) ;
    buf_clk cell_10462 ( .C (clk), .D (signal_15349), .Q (signal_15350) ) ;
    buf_clk cell_10470 ( .C (clk), .D (signal_15357), .Q (signal_15358) ) ;
    buf_clk cell_10478 ( .C (clk), .D (signal_15365), .Q (signal_15366) ) ;
    buf_clk cell_10486 ( .C (clk), .D (signal_15373), .Q (signal_15374) ) ;
    buf_clk cell_10494 ( .C (clk), .D (signal_15381), .Q (signal_15382) ) ;
    buf_clk cell_10502 ( .C (clk), .D (signal_15389), .Q (signal_15390) ) ;
    buf_clk cell_10510 ( .C (clk), .D (signal_15397), .Q (signal_15398) ) ;
    buf_clk cell_10518 ( .C (clk), .D (signal_15405), .Q (signal_15406) ) ;
    buf_clk cell_10526 ( .C (clk), .D (signal_15413), .Q (signal_15414) ) ;
    buf_clk cell_10534 ( .C (clk), .D (signal_15421), .Q (signal_15422) ) ;
    buf_clk cell_10542 ( .C (clk), .D (signal_15429), .Q (signal_15430) ) ;
    buf_clk cell_10550 ( .C (clk), .D (signal_15437), .Q (signal_15438) ) ;
    buf_clk cell_10558 ( .C (clk), .D (signal_15445), .Q (signal_15446) ) ;
    buf_clk cell_10566 ( .C (clk), .D (signal_15453), .Q (signal_15454) ) ;
    buf_clk cell_10574 ( .C (clk), .D (signal_15461), .Q (signal_15462) ) ;
    buf_clk cell_10582 ( .C (clk), .D (signal_15469), .Q (signal_15470) ) ;
    buf_clk cell_10590 ( .C (clk), .D (signal_15477), .Q (signal_15478) ) ;
    buf_clk cell_10598 ( .C (clk), .D (signal_15485), .Q (signal_15486) ) ;
    buf_clk cell_10606 ( .C (clk), .D (signal_15493), .Q (signal_15494) ) ;
    buf_clk cell_10614 ( .C (clk), .D (signal_15501), .Q (signal_15502) ) ;
    buf_clk cell_10622 ( .C (clk), .D (signal_15509), .Q (signal_15510) ) ;
    buf_clk cell_10630 ( .C (clk), .D (signal_15517), .Q (signal_15518) ) ;
    buf_clk cell_10638 ( .C (clk), .D (signal_15525), .Q (signal_15526) ) ;
    buf_clk cell_10646 ( .C (clk), .D (signal_15533), .Q (signal_15534) ) ;
    buf_clk cell_10654 ( .C (clk), .D (signal_15541), .Q (signal_15542) ) ;
    buf_clk cell_10662 ( .C (clk), .D (signal_15549), .Q (signal_15550) ) ;
    buf_clk cell_10670 ( .C (clk), .D (signal_15557), .Q (signal_15558) ) ;
    buf_clk cell_10678 ( .C (clk), .D (signal_15565), .Q (signal_15566) ) ;
    buf_clk cell_10686 ( .C (clk), .D (signal_15573), .Q (signal_15574) ) ;
    buf_clk cell_10694 ( .C (clk), .D (signal_15581), .Q (signal_15582) ) ;
    buf_clk cell_10702 ( .C (clk), .D (signal_15589), .Q (signal_15590) ) ;
    buf_clk cell_10710 ( .C (clk), .D (signal_15597), .Q (signal_15598) ) ;
    buf_clk cell_10718 ( .C (clk), .D (signal_15605), .Q (signal_15606) ) ;
    buf_clk cell_10726 ( .C (clk), .D (signal_15613), .Q (signal_15614) ) ;
    buf_clk cell_10734 ( .C (clk), .D (signal_15621), .Q (signal_15622) ) ;
    buf_clk cell_10742 ( .C (clk), .D (signal_15629), .Q (signal_15630) ) ;
    buf_clk cell_10750 ( .C (clk), .D (signal_15637), .Q (signal_15638) ) ;
    buf_clk cell_10758 ( .C (clk), .D (signal_15645), .Q (signal_15646) ) ;
    buf_clk cell_10766 ( .C (clk), .D (signal_15653), .Q (signal_15654) ) ;
    buf_clk cell_10774 ( .C (clk), .D (signal_15661), .Q (signal_15662) ) ;
    buf_clk cell_10782 ( .C (clk), .D (signal_15669), .Q (signal_15670) ) ;
    buf_clk cell_10790 ( .C (clk), .D (signal_15677), .Q (signal_15678) ) ;
    buf_clk cell_10798 ( .C (clk), .D (signal_15685), .Q (signal_15686) ) ;
    buf_clk cell_10806 ( .C (clk), .D (signal_15693), .Q (signal_15694) ) ;
    buf_clk cell_10814 ( .C (clk), .D (signal_15701), .Q (signal_15702) ) ;
    buf_clk cell_10822 ( .C (clk), .D (signal_15709), .Q (signal_15710) ) ;
    buf_clk cell_10830 ( .C (clk), .D (signal_15717), .Q (signal_15718) ) ;
    buf_clk cell_10838 ( .C (clk), .D (signal_15725), .Q (signal_15726) ) ;
    buf_clk cell_10846 ( .C (clk), .D (signal_15733), .Q (signal_15734) ) ;
    buf_clk cell_10854 ( .C (clk), .D (signal_15741), .Q (signal_15742) ) ;
    buf_clk cell_10862 ( .C (clk), .D (signal_15749), .Q (signal_15750) ) ;
    buf_clk cell_10870 ( .C (clk), .D (signal_15757), .Q (signal_15758) ) ;
    buf_clk cell_10878 ( .C (clk), .D (signal_15765), .Q (signal_15766) ) ;
    buf_clk cell_10886 ( .C (clk), .D (signal_15773), .Q (signal_15774) ) ;
    buf_clk cell_10894 ( .C (clk), .D (signal_15781), .Q (signal_15782) ) ;
    buf_clk cell_10902 ( .C (clk), .D (signal_15789), .Q (signal_15790) ) ;
    buf_clk cell_10910 ( .C (clk), .D (signal_15797), .Q (signal_15798) ) ;
    buf_clk cell_10918 ( .C (clk), .D (signal_15805), .Q (signal_15806) ) ;
    buf_clk cell_10926 ( .C (clk), .D (signal_15813), .Q (signal_15814) ) ;
    buf_clk cell_10934 ( .C (clk), .D (signal_15821), .Q (signal_15822) ) ;
    buf_clk cell_10942 ( .C (clk), .D (signal_15829), .Q (signal_15830) ) ;
    buf_clk cell_10950 ( .C (clk), .D (signal_15837), .Q (signal_15838) ) ;
    buf_clk cell_10958 ( .C (clk), .D (signal_15845), .Q (signal_15846) ) ;
    buf_clk cell_10966 ( .C (clk), .D (signal_15853), .Q (signal_15854) ) ;
    buf_clk cell_10974 ( .C (clk), .D (signal_15861), .Q (signal_15862) ) ;
    buf_clk cell_10982 ( .C (clk), .D (signal_15869), .Q (signal_15870) ) ;
    buf_clk cell_10990 ( .C (clk), .D (signal_15877), .Q (signal_15878) ) ;
    buf_clk cell_10998 ( .C (clk), .D (signal_15885), .Q (signal_15886) ) ;
    buf_clk cell_11006 ( .C (clk), .D (signal_15893), .Q (signal_15894) ) ;
    buf_clk cell_11014 ( .C (clk), .D (signal_15901), .Q (signal_15902) ) ;
    buf_clk cell_11022 ( .C (clk), .D (signal_15909), .Q (signal_15910) ) ;
    buf_clk cell_11030 ( .C (clk), .D (signal_15917), .Q (signal_15918) ) ;
    buf_clk cell_11038 ( .C (clk), .D (signal_15925), .Q (signal_15926) ) ;
    buf_clk cell_11046 ( .C (clk), .D (signal_15933), .Q (signal_15934) ) ;
    buf_clk cell_11054 ( .C (clk), .D (signal_15941), .Q (signal_15942) ) ;
    buf_clk cell_11062 ( .C (clk), .D (signal_15949), .Q (signal_15950) ) ;
    buf_clk cell_11070 ( .C (clk), .D (signal_15957), .Q (signal_15958) ) ;
    buf_clk cell_11078 ( .C (clk), .D (signal_15965), .Q (signal_15966) ) ;
    buf_clk cell_11086 ( .C (clk), .D (signal_15973), .Q (signal_15974) ) ;
    buf_clk cell_11094 ( .C (clk), .D (signal_15981), .Q (signal_15982) ) ;
    buf_clk cell_11102 ( .C (clk), .D (signal_15989), .Q (signal_15990) ) ;
    buf_clk cell_11110 ( .C (clk), .D (signal_15997), .Q (signal_15998) ) ;
    buf_clk cell_11118 ( .C (clk), .D (signal_16005), .Q (signal_16006) ) ;
    buf_clk cell_11126 ( .C (clk), .D (signal_16013), .Q (signal_16014) ) ;
    buf_clk cell_11134 ( .C (clk), .D (signal_16021), .Q (signal_16022) ) ;
    buf_clk cell_11142 ( .C (clk), .D (signal_16029), .Q (signal_16030) ) ;
    buf_clk cell_11150 ( .C (clk), .D (signal_16037), .Q (signal_16038) ) ;
    buf_clk cell_11158 ( .C (clk), .D (signal_16045), .Q (signal_16046) ) ;
    buf_clk cell_11166 ( .C (clk), .D (signal_16053), .Q (signal_16054) ) ;
    buf_clk cell_11174 ( .C (clk), .D (signal_16061), .Q (signal_16062) ) ;
    buf_clk cell_11182 ( .C (clk), .D (signal_16069), .Q (signal_16070) ) ;
    buf_clk cell_11190 ( .C (clk), .D (signal_16077), .Q (signal_16078) ) ;
    buf_clk cell_11198 ( .C (clk), .D (signal_16085), .Q (signal_16086) ) ;
    buf_clk cell_11206 ( .C (clk), .D (signal_16093), .Q (signal_16094) ) ;
    buf_clk cell_11214 ( .C (clk), .D (signal_16101), .Q (signal_16102) ) ;
    buf_clk cell_11222 ( .C (clk), .D (signal_16109), .Q (signal_16110) ) ;
    buf_clk cell_11230 ( .C (clk), .D (signal_16117), .Q (signal_16118) ) ;
    buf_clk cell_11238 ( .C (clk), .D (signal_16125), .Q (signal_16126) ) ;
    buf_clk cell_11246 ( .C (clk), .D (signal_16133), .Q (signal_16134) ) ;
    buf_clk cell_11254 ( .C (clk), .D (signal_16141), .Q (signal_16142) ) ;
    buf_clk cell_11262 ( .C (clk), .D (signal_16149), .Q (signal_16150) ) ;
    buf_clk cell_11270 ( .C (clk), .D (signal_16157), .Q (signal_16158) ) ;
    buf_clk cell_11278 ( .C (clk), .D (signal_16165), .Q (signal_16166) ) ;
    buf_clk cell_11286 ( .C (clk), .D (signal_16173), .Q (signal_16174) ) ;
    buf_clk cell_11294 ( .C (clk), .D (signal_16181), .Q (signal_16182) ) ;
    buf_clk cell_11302 ( .C (clk), .D (signal_16189), .Q (signal_16190) ) ;
    buf_clk cell_11310 ( .C (clk), .D (signal_16197), .Q (signal_16198) ) ;
    buf_clk cell_11318 ( .C (clk), .D (signal_16205), .Q (signal_16206) ) ;
    buf_clk cell_11326 ( .C (clk), .D (signal_16213), .Q (signal_16214) ) ;
    buf_clk cell_11334 ( .C (clk), .D (signal_16221), .Q (signal_16222) ) ;
    buf_clk cell_11342 ( .C (clk), .D (signal_16229), .Q (signal_16230) ) ;
    buf_clk cell_11350 ( .C (clk), .D (signal_16237), .Q (signal_16238) ) ;
    buf_clk cell_11358 ( .C (clk), .D (signal_16245), .Q (signal_16246) ) ;
    buf_clk cell_11366 ( .C (clk), .D (signal_16253), .Q (signal_16254) ) ;
    buf_clk cell_11374 ( .C (clk), .D (signal_16261), .Q (signal_16262) ) ;
    buf_clk cell_11382 ( .C (clk), .D (signal_16269), .Q (signal_16270) ) ;
    buf_clk cell_11390 ( .C (clk), .D (signal_16277), .Q (signal_16278) ) ;
    buf_clk cell_11398 ( .C (clk), .D (signal_16285), .Q (signal_16286) ) ;
    buf_clk cell_11406 ( .C (clk), .D (signal_16293), .Q (signal_16294) ) ;
    buf_clk cell_11414 ( .C (clk), .D (signal_16301), .Q (signal_16302) ) ;
    buf_clk cell_11422 ( .C (clk), .D (signal_16309), .Q (signal_16310) ) ;
    buf_clk cell_11430 ( .C (clk), .D (signal_16317), .Q (signal_16318) ) ;
    buf_clk cell_11438 ( .C (clk), .D (signal_16325), .Q (signal_16326) ) ;
    buf_clk cell_11446 ( .C (clk), .D (signal_16333), .Q (signal_16334) ) ;
    buf_clk cell_11454 ( .C (clk), .D (signal_16341), .Q (signal_16342) ) ;
    buf_clk cell_11462 ( .C (clk), .D (signal_16349), .Q (signal_16350) ) ;
    buf_clk cell_11470 ( .C (clk), .D (signal_16357), .Q (signal_16358) ) ;
    buf_clk cell_11478 ( .C (clk), .D (signal_16365), .Q (signal_16366) ) ;
    buf_clk cell_11486 ( .C (clk), .D (signal_16373), .Q (signal_16374) ) ;
    buf_clk cell_11494 ( .C (clk), .D (signal_16381), .Q (signal_16382) ) ;
    buf_clk cell_11502 ( .C (clk), .D (signal_16389), .Q (signal_16390) ) ;
    buf_clk cell_11510 ( .C (clk), .D (signal_16397), .Q (signal_16398) ) ;
    buf_clk cell_11518 ( .C (clk), .D (signal_16405), .Q (signal_16406) ) ;
    buf_clk cell_11526 ( .C (clk), .D (signal_16413), .Q (signal_16414) ) ;
    buf_clk cell_11534 ( .C (clk), .D (signal_16421), .Q (signal_16422) ) ;
    buf_clk cell_11542 ( .C (clk), .D (signal_16429), .Q (signal_16430) ) ;
    buf_clk cell_11550 ( .C (clk), .D (signal_16437), .Q (signal_16438) ) ;
    buf_clk cell_11558 ( .C (clk), .D (signal_16445), .Q (signal_16446) ) ;
    buf_clk cell_11566 ( .C (clk), .D (signal_16453), .Q (signal_16454) ) ;
    buf_clk cell_11574 ( .C (clk), .D (signal_16461), .Q (signal_16462) ) ;
    buf_clk cell_11582 ( .C (clk), .D (signal_16469), .Q (signal_16470) ) ;
    buf_clk cell_11590 ( .C (clk), .D (signal_16477), .Q (signal_16478) ) ;
    buf_clk cell_11598 ( .C (clk), .D (signal_16485), .Q (signal_16486) ) ;
    buf_clk cell_11606 ( .C (clk), .D (signal_16493), .Q (signal_16494) ) ;
    buf_clk cell_11614 ( .C (clk), .D (signal_16501), .Q (signal_16502) ) ;
    buf_clk cell_11622 ( .C (clk), .D (signal_16509), .Q (signal_16510) ) ;
    buf_clk cell_11630 ( .C (clk), .D (signal_16517), .Q (signal_16518) ) ;
    buf_clk cell_11638 ( .C (clk), .D (signal_16525), .Q (signal_16526) ) ;
    buf_clk cell_11646 ( .C (clk), .D (signal_16533), .Q (signal_16534) ) ;
    buf_clk cell_11654 ( .C (clk), .D (signal_16541), .Q (signal_16542) ) ;
    buf_clk cell_11662 ( .C (clk), .D (signal_16549), .Q (signal_16550) ) ;
    buf_clk cell_11670 ( .C (clk), .D (signal_16557), .Q (signal_16558) ) ;
    buf_clk cell_11678 ( .C (clk), .D (signal_16565), .Q (signal_16566) ) ;
    buf_clk cell_11686 ( .C (clk), .D (signal_16573), .Q (signal_16574) ) ;
    buf_clk cell_11694 ( .C (clk), .D (signal_16581), .Q (signal_16582) ) ;
    buf_clk cell_11702 ( .C (clk), .D (signal_16589), .Q (signal_16590) ) ;
    buf_clk cell_11710 ( .C (clk), .D (signal_16597), .Q (signal_16598) ) ;
    buf_clk cell_11718 ( .C (clk), .D (signal_16605), .Q (signal_16606) ) ;
    buf_clk cell_11726 ( .C (clk), .D (signal_16613), .Q (signal_16614) ) ;
    buf_clk cell_11734 ( .C (clk), .D (signal_16621), .Q (signal_16622) ) ;
    buf_clk cell_11742 ( .C (clk), .D (signal_16629), .Q (signal_16630) ) ;
    buf_clk cell_11750 ( .C (clk), .D (signal_16637), .Q (signal_16638) ) ;
    buf_clk cell_11758 ( .C (clk), .D (signal_16645), .Q (signal_16646) ) ;
    buf_clk cell_11766 ( .C (clk), .D (signal_16653), .Q (signal_16654) ) ;
    buf_clk cell_11774 ( .C (clk), .D (signal_16661), .Q (signal_16662) ) ;
    buf_clk cell_11782 ( .C (clk), .D (signal_16669), .Q (signal_16670) ) ;
    buf_clk cell_11790 ( .C (clk), .D (signal_16677), .Q (signal_16678) ) ;
    buf_clk cell_11798 ( .C (clk), .D (signal_16685), .Q (signal_16686) ) ;
    buf_clk cell_11806 ( .C (clk), .D (signal_16693), .Q (signal_16694) ) ;
    buf_clk cell_11814 ( .C (clk), .D (signal_16701), .Q (signal_16702) ) ;
    buf_clk cell_11822 ( .C (clk), .D (signal_16709), .Q (signal_16710) ) ;
    buf_clk cell_11830 ( .C (clk), .D (signal_16717), .Q (signal_16718) ) ;
    buf_clk cell_11838 ( .C (clk), .D (signal_16725), .Q (signal_16726) ) ;
    buf_clk cell_11846 ( .C (clk), .D (signal_16733), .Q (signal_16734) ) ;
    buf_clk cell_11854 ( .C (clk), .D (signal_16741), .Q (signal_16742) ) ;
    buf_clk cell_11862 ( .C (clk), .D (signal_16749), .Q (signal_16750) ) ;
    buf_clk cell_11870 ( .C (clk), .D (signal_16757), .Q (signal_16758) ) ;
    buf_clk cell_11878 ( .C (clk), .D (signal_16765), .Q (signal_16766) ) ;
    buf_clk cell_11886 ( .C (clk), .D (signal_16773), .Q (signal_16774) ) ;
    buf_clk cell_11894 ( .C (clk), .D (signal_16781), .Q (signal_16782) ) ;
    buf_clk cell_11902 ( .C (clk), .D (signal_16789), .Q (signal_16790) ) ;
    buf_clk cell_11910 ( .C (clk), .D (signal_16797), .Q (signal_16798) ) ;
    buf_clk cell_11918 ( .C (clk), .D (signal_16805), .Q (signal_16806) ) ;
    buf_clk cell_11926 ( .C (clk), .D (signal_16813), .Q (signal_16814) ) ;
    buf_clk cell_11934 ( .C (clk), .D (signal_16821), .Q (signal_16822) ) ;
    buf_clk cell_11942 ( .C (clk), .D (signal_16829), .Q (signal_16830) ) ;
    buf_clk cell_11950 ( .C (clk), .D (signal_16837), .Q (signal_16838) ) ;
    buf_clk cell_11958 ( .C (clk), .D (signal_16845), .Q (signal_16846) ) ;
    buf_clk cell_11966 ( .C (clk), .D (signal_16853), .Q (signal_16854) ) ;
    buf_clk cell_11974 ( .C (clk), .D (signal_16861), .Q (signal_16862) ) ;
    buf_clk cell_11982 ( .C (clk), .D (signal_16869), .Q (signal_16870) ) ;
    buf_clk cell_11990 ( .C (clk), .D (signal_16877), .Q (signal_16878) ) ;
    buf_clk cell_11998 ( .C (clk), .D (signal_16885), .Q (signal_16886) ) ;
    buf_clk cell_12006 ( .C (clk), .D (signal_16893), .Q (signal_16894) ) ;
    buf_clk cell_12014 ( .C (clk), .D (signal_16901), .Q (signal_16902) ) ;
    buf_clk cell_12022 ( .C (clk), .D (signal_16909), .Q (signal_16910) ) ;
    buf_clk cell_12030 ( .C (clk), .D (signal_16917), .Q (signal_16918) ) ;
    buf_clk cell_12038 ( .C (clk), .D (signal_16925), .Q (signal_16926) ) ;
    buf_clk cell_12046 ( .C (clk), .D (signal_16933), .Q (signal_16934) ) ;
    buf_clk cell_12054 ( .C (clk), .D (signal_16941), .Q (signal_16942) ) ;
    buf_clk cell_12062 ( .C (clk), .D (signal_16949), .Q (signal_16950) ) ;
    buf_clk cell_12070 ( .C (clk), .D (signal_16957), .Q (signal_16958) ) ;
    buf_clk cell_12078 ( .C (clk), .D (signal_16965), .Q (signal_16966) ) ;
    buf_clk cell_12086 ( .C (clk), .D (signal_16973), .Q (signal_16974) ) ;
    buf_clk cell_12094 ( .C (clk), .D (signal_16981), .Q (signal_16982) ) ;
    buf_clk cell_12102 ( .C (clk), .D (signal_16989), .Q (signal_16990) ) ;
    buf_clk cell_12110 ( .C (clk), .D (signal_16997), .Q (signal_16998) ) ;
    buf_clk cell_12118 ( .C (clk), .D (signal_17005), .Q (signal_17006) ) ;
    buf_clk cell_12126 ( .C (clk), .D (signal_17013), .Q (signal_17014) ) ;
    buf_clk cell_12134 ( .C (clk), .D (signal_17021), .Q (signal_17022) ) ;
    buf_clk cell_12142 ( .C (clk), .D (signal_17029), .Q (signal_17030) ) ;
    buf_clk cell_12150 ( .C (clk), .D (signal_17037), .Q (signal_17038) ) ;
    buf_clk cell_12158 ( .C (clk), .D (signal_17045), .Q (signal_17046) ) ;
    buf_clk cell_12166 ( .C (clk), .D (signal_17053), .Q (signal_17054) ) ;
    buf_clk cell_12174 ( .C (clk), .D (signal_17061), .Q (signal_17062) ) ;
    buf_clk cell_12182 ( .C (clk), .D (signal_17069), .Q (signal_17070) ) ;
    buf_clk cell_12190 ( .C (clk), .D (signal_17077), .Q (signal_17078) ) ;
    buf_clk cell_12198 ( .C (clk), .D (signal_17085), .Q (signal_17086) ) ;
    buf_clk cell_12206 ( .C (clk), .D (signal_17093), .Q (signal_17094) ) ;
    buf_clk cell_12214 ( .C (clk), .D (signal_17101), .Q (signal_17102) ) ;
    buf_clk cell_12222 ( .C (clk), .D (signal_17109), .Q (signal_17110) ) ;
    buf_clk cell_12230 ( .C (clk), .D (signal_17117), .Q (signal_17118) ) ;
    buf_clk cell_12238 ( .C (clk), .D (signal_17125), .Q (signal_17126) ) ;
    buf_clk cell_12246 ( .C (clk), .D (signal_17133), .Q (signal_17134) ) ;
    buf_clk cell_12254 ( .C (clk), .D (signal_17141), .Q (signal_17142) ) ;
    buf_clk cell_12262 ( .C (clk), .D (signal_17149), .Q (signal_17150) ) ;
    buf_clk cell_12270 ( .C (clk), .D (signal_17157), .Q (signal_17158) ) ;
    buf_clk cell_12278 ( .C (clk), .D (signal_17165), .Q (signal_17166) ) ;
    buf_clk cell_12286 ( .C (clk), .D (signal_17173), .Q (signal_17174) ) ;
    buf_clk cell_12294 ( .C (clk), .D (signal_17181), .Q (signal_17182) ) ;
    buf_clk cell_12302 ( .C (clk), .D (signal_17189), .Q (signal_17190) ) ;
    buf_clk cell_12310 ( .C (clk), .D (signal_17197), .Q (signal_17198) ) ;
    buf_clk cell_12318 ( .C (clk), .D (signal_17205), .Q (signal_17206) ) ;
    buf_clk cell_12326 ( .C (clk), .D (signal_17213), .Q (signal_17214) ) ;
    buf_clk cell_12334 ( .C (clk), .D (signal_17221), .Q (signal_17222) ) ;
    buf_clk cell_12342 ( .C (clk), .D (signal_17229), .Q (signal_17230) ) ;
    buf_clk cell_12350 ( .C (clk), .D (signal_17237), .Q (signal_17238) ) ;
    buf_clk cell_12358 ( .C (clk), .D (signal_17245), .Q (signal_17246) ) ;
    buf_clk cell_12366 ( .C (clk), .D (signal_17253), .Q (signal_17254) ) ;
    buf_clk cell_12374 ( .C (clk), .D (signal_17261), .Q (signal_17262) ) ;
    buf_clk cell_12382 ( .C (clk), .D (signal_17269), .Q (signal_17270) ) ;
    buf_clk cell_12390 ( .C (clk), .D (signal_17277), .Q (signal_17278) ) ;
    buf_clk cell_12398 ( .C (clk), .D (signal_17285), .Q (signal_17286) ) ;
    buf_clk cell_12406 ( .C (clk), .D (signal_17293), .Q (signal_17294) ) ;
    buf_clk cell_12414 ( .C (clk), .D (signal_17301), .Q (signal_17302) ) ;
    buf_clk cell_12422 ( .C (clk), .D (signal_17309), .Q (signal_17310) ) ;
    buf_clk cell_12430 ( .C (clk), .D (signal_17317), .Q (signal_17318) ) ;
    buf_clk cell_12438 ( .C (clk), .D (signal_17325), .Q (signal_17326) ) ;
    buf_clk cell_12446 ( .C (clk), .D (signal_17333), .Q (signal_17334) ) ;
    buf_clk cell_12454 ( .C (clk), .D (signal_17341), .Q (signal_17342) ) ;
    buf_clk cell_12462 ( .C (clk), .D (signal_17349), .Q (signal_17350) ) ;
    buf_clk cell_12470 ( .C (clk), .D (signal_17357), .Q (signal_17358) ) ;
    buf_clk cell_12478 ( .C (clk), .D (signal_17365), .Q (signal_17366) ) ;
    buf_clk cell_12486 ( .C (clk), .D (signal_17373), .Q (signal_17374) ) ;
    buf_clk cell_12494 ( .C (clk), .D (signal_17381), .Q (signal_17382) ) ;
    buf_clk cell_12502 ( .C (clk), .D (signal_17389), .Q (signal_17390) ) ;
    buf_clk cell_12510 ( .C (clk), .D (signal_17397), .Q (signal_17398) ) ;
    buf_clk cell_12518 ( .C (clk), .D (signal_17405), .Q (signal_17406) ) ;
    buf_clk cell_12526 ( .C (clk), .D (signal_17413), .Q (signal_17414) ) ;
    buf_clk cell_12534 ( .C (clk), .D (signal_17421), .Q (signal_17422) ) ;
    buf_clk cell_12542 ( .C (clk), .D (signal_17429), .Q (signal_17430) ) ;
    buf_clk cell_12550 ( .C (clk), .D (signal_17437), .Q (signal_17438) ) ;
    buf_clk cell_12558 ( .C (clk), .D (signal_17445), .Q (signal_17446) ) ;
    buf_clk cell_12566 ( .C (clk), .D (signal_17453), .Q (signal_17454) ) ;
    buf_clk cell_12574 ( .C (clk), .D (signal_17461), .Q (signal_17462) ) ;
    buf_clk cell_12582 ( .C (clk), .D (signal_17469), .Q (signal_17470) ) ;
    buf_clk cell_12590 ( .C (clk), .D (signal_17477), .Q (signal_17478) ) ;
    buf_clk cell_12598 ( .C (clk), .D (signal_17485), .Q (signal_17486) ) ;
    buf_clk cell_12606 ( .C (clk), .D (signal_17493), .Q (signal_17494) ) ;
    buf_clk cell_12614 ( .C (clk), .D (signal_17501), .Q (signal_17502) ) ;
    buf_clk cell_12622 ( .C (clk), .D (signal_17509), .Q (signal_17510) ) ;
    buf_clk cell_12630 ( .C (clk), .D (signal_17517), .Q (signal_17518) ) ;
    buf_clk cell_12638 ( .C (clk), .D (signal_17525), .Q (signal_17526) ) ;
    buf_clk cell_12646 ( .C (clk), .D (signal_17533), .Q (signal_17534) ) ;
    buf_clk cell_12654 ( .C (clk), .D (signal_17541), .Q (signal_17542) ) ;
    buf_clk cell_12662 ( .C (clk), .D (signal_17549), .Q (signal_17550) ) ;
    buf_clk cell_12670 ( .C (clk), .D (signal_17557), .Q (signal_17558) ) ;
    buf_clk cell_12678 ( .C (clk), .D (signal_17565), .Q (signal_17566) ) ;
    buf_clk cell_12686 ( .C (clk), .D (signal_17573), .Q (signal_17574) ) ;
    buf_clk cell_12694 ( .C (clk), .D (signal_17581), .Q (signal_17582) ) ;
    buf_clk cell_12702 ( .C (clk), .D (signal_17589), .Q (signal_17590) ) ;
    buf_clk cell_12710 ( .C (clk), .D (signal_17597), .Q (signal_17598) ) ;
    buf_clk cell_12718 ( .C (clk), .D (signal_17605), .Q (signal_17606) ) ;
    buf_clk cell_12726 ( .C (clk), .D (signal_17613), .Q (signal_17614) ) ;
    buf_clk cell_12734 ( .C (clk), .D (signal_17621), .Q (signal_17622) ) ;
    buf_clk cell_12742 ( .C (clk), .D (signal_17629), .Q (signal_17630) ) ;
    buf_clk cell_12750 ( .C (clk), .D (signal_17637), .Q (signal_17638) ) ;
    buf_clk cell_12758 ( .C (clk), .D (signal_17645), .Q (signal_17646) ) ;
    buf_clk cell_12766 ( .C (clk), .D (signal_17653), .Q (signal_17654) ) ;
    buf_clk cell_12774 ( .C (clk), .D (signal_17661), .Q (signal_17662) ) ;
    buf_clk cell_12782 ( .C (clk), .D (signal_17669), .Q (signal_17670) ) ;
    buf_clk cell_12790 ( .C (clk), .D (signal_17677), .Q (signal_17678) ) ;
    buf_clk cell_12798 ( .C (clk), .D (signal_17685), .Q (signal_17686) ) ;
    buf_clk cell_12806 ( .C (clk), .D (signal_17693), .Q (signal_17694) ) ;
    buf_clk cell_12814 ( .C (clk), .D (signal_17701), .Q (signal_17702) ) ;
    buf_clk cell_12822 ( .C (clk), .D (signal_17709), .Q (signal_17710) ) ;
    buf_clk cell_12830 ( .C (clk), .D (signal_17717), .Q (signal_17718) ) ;
    buf_clk cell_12838 ( .C (clk), .D (signal_17725), .Q (signal_17726) ) ;
    buf_clk cell_12846 ( .C (clk), .D (signal_17733), .Q (signal_17734) ) ;
    buf_clk cell_12854 ( .C (clk), .D (signal_17741), .Q (signal_17742) ) ;
    buf_clk cell_12862 ( .C (clk), .D (signal_17749), .Q (signal_17750) ) ;
    buf_clk cell_12870 ( .C (clk), .D (signal_17757), .Q (signal_17758) ) ;
    buf_clk cell_12878 ( .C (clk), .D (signal_17765), .Q (signal_17766) ) ;
    buf_clk cell_12886 ( .C (clk), .D (signal_17773), .Q (signal_17774) ) ;
    buf_clk cell_12894 ( .C (clk), .D (signal_17781), .Q (signal_17782) ) ;
    buf_clk cell_12902 ( .C (clk), .D (signal_17789), .Q (signal_17790) ) ;
    buf_clk cell_12910 ( .C (clk), .D (signal_17797), .Q (signal_17798) ) ;
    buf_clk cell_12918 ( .C (clk), .D (signal_17805), .Q (signal_17806) ) ;
    buf_clk cell_12926 ( .C (clk), .D (signal_17813), .Q (signal_17814) ) ;
    buf_clk cell_12934 ( .C (clk), .D (signal_17821), .Q (signal_17822) ) ;
    buf_clk cell_12942 ( .C (clk), .D (signal_17829), .Q (signal_17830) ) ;
    buf_clk cell_12950 ( .C (clk), .D (signal_17837), .Q (signal_17838) ) ;
    buf_clk cell_12958 ( .C (clk), .D (signal_17845), .Q (signal_17846) ) ;
    buf_clk cell_12966 ( .C (clk), .D (signal_17853), .Q (signal_17854) ) ;
    buf_clk cell_12974 ( .C (clk), .D (signal_17861), .Q (signal_17862) ) ;
    buf_clk cell_12982 ( .C (clk), .D (signal_17869), .Q (signal_17870) ) ;
    buf_clk cell_12990 ( .C (clk), .D (signal_17877), .Q (signal_17878) ) ;
    buf_clk cell_12998 ( .C (clk), .D (signal_17885), .Q (signal_17886) ) ;
    buf_clk cell_13006 ( .C (clk), .D (signal_17893), .Q (signal_17894) ) ;
    buf_clk cell_13014 ( .C (clk), .D (signal_17901), .Q (signal_17902) ) ;
    buf_clk cell_13022 ( .C (clk), .D (signal_17909), .Q (signal_17910) ) ;
    buf_clk cell_13030 ( .C (clk), .D (signal_17917), .Q (signal_17918) ) ;
    buf_clk cell_13038 ( .C (clk), .D (signal_17925), .Q (signal_17926) ) ;
    buf_clk cell_13046 ( .C (clk), .D (signal_17933), .Q (signal_17934) ) ;
    buf_clk cell_13054 ( .C (clk), .D (signal_17941), .Q (signal_17942) ) ;
    buf_clk cell_13062 ( .C (clk), .D (signal_17949), .Q (signal_17950) ) ;
    buf_clk cell_13070 ( .C (clk), .D (signal_17957), .Q (signal_17958) ) ;
    buf_clk cell_13078 ( .C (clk), .D (signal_17965), .Q (signal_17966) ) ;
    buf_clk cell_13086 ( .C (clk), .D (signal_17973), .Q (signal_17974) ) ;
    buf_clk cell_13094 ( .C (clk), .D (signal_17981), .Q (signal_17982) ) ;
    buf_clk cell_13102 ( .C (clk), .D (signal_17989), .Q (signal_17990) ) ;
    buf_clk cell_13110 ( .C (clk), .D (signal_17997), .Q (signal_17998) ) ;
    buf_clk cell_13118 ( .C (clk), .D (signal_18005), .Q (signal_18006) ) ;
    buf_clk cell_13126 ( .C (clk), .D (signal_18013), .Q (signal_18014) ) ;
    buf_clk cell_13134 ( .C (clk), .D (signal_18021), .Q (signal_18022) ) ;
    buf_clk cell_13142 ( .C (clk), .D (signal_18029), .Q (signal_18030) ) ;
    buf_clk cell_13150 ( .C (clk), .D (signal_18037), .Q (signal_18038) ) ;
    buf_clk cell_13158 ( .C (clk), .D (signal_18045), .Q (signal_18046) ) ;
    buf_clk cell_13166 ( .C (clk), .D (signal_18053), .Q (signal_18054) ) ;
    buf_clk cell_13174 ( .C (clk), .D (signal_18061), .Q (signal_18062) ) ;
    buf_clk cell_13182 ( .C (clk), .D (signal_18069), .Q (signal_18070) ) ;
    buf_clk cell_13190 ( .C (clk), .D (signal_18077), .Q (signal_18078) ) ;
    buf_clk cell_13198 ( .C (clk), .D (signal_18085), .Q (signal_18086) ) ;
    buf_clk cell_13206 ( .C (clk), .D (signal_18093), .Q (signal_18094) ) ;
    buf_clk cell_13214 ( .C (clk), .D (signal_18101), .Q (signal_18102) ) ;
    buf_clk cell_13222 ( .C (clk), .D (signal_18109), .Q (signal_18110) ) ;
    buf_clk cell_13230 ( .C (clk), .D (signal_18117), .Q (signal_18118) ) ;
    buf_clk cell_13238 ( .C (clk), .D (signal_18125), .Q (signal_18126) ) ;
    buf_clk cell_13246 ( .C (clk), .D (signal_18133), .Q (signal_18134) ) ;
    buf_clk cell_13254 ( .C (clk), .D (signal_18141), .Q (signal_18142) ) ;
    buf_clk cell_13262 ( .C (clk), .D (signal_18149), .Q (signal_18150) ) ;
    buf_clk cell_13270 ( .C (clk), .D (signal_18157), .Q (signal_18158) ) ;
    buf_clk cell_13278 ( .C (clk), .D (signal_18165), .Q (signal_18166) ) ;
    buf_clk cell_13284 ( .C (clk), .D (signal_18171), .Q (signal_18172) ) ;
    buf_clk cell_13290 ( .C (clk), .D (signal_18177), .Q (signal_18178) ) ;
    buf_clk cell_13296 ( .C (clk), .D (signal_18183), .Q (signal_18184) ) ;
    buf_clk cell_13302 ( .C (clk), .D (signal_18189), .Q (signal_18190) ) ;
    buf_clk cell_13308 ( .C (clk), .D (signal_18195), .Q (signal_18196) ) ;
    buf_clk cell_13314 ( .C (clk), .D (signal_18201), .Q (signal_18202) ) ;
    buf_clk cell_13320 ( .C (clk), .D (signal_18207), .Q (signal_18208) ) ;
    buf_clk cell_13326 ( .C (clk), .D (signal_18213), .Q (signal_18214) ) ;
    buf_clk cell_13332 ( .C (clk), .D (signal_18219), .Q (signal_18220) ) ;
    buf_clk cell_13338 ( .C (clk), .D (signal_18225), .Q (signal_18226) ) ;
    buf_clk cell_13344 ( .C (clk), .D (signal_18231), .Q (signal_18232) ) ;
    buf_clk cell_13350 ( .C (clk), .D (signal_18237), .Q (signal_18238) ) ;
    buf_clk cell_13356 ( .C (clk), .D (signal_18243), .Q (signal_18244) ) ;
    buf_clk cell_13362 ( .C (clk), .D (signal_18249), .Q (signal_18250) ) ;
    buf_clk cell_13368 ( .C (clk), .D (signal_18255), .Q (signal_18256) ) ;
    buf_clk cell_13374 ( .C (clk), .D (signal_18261), .Q (signal_18262) ) ;
    buf_clk cell_13380 ( .C (clk), .D (signal_18267), .Q (signal_18268) ) ;
    buf_clk cell_13386 ( .C (clk), .D (signal_18273), .Q (signal_18274) ) ;
    buf_clk cell_13392 ( .C (clk), .D (signal_18279), .Q (signal_18280) ) ;
    buf_clk cell_13398 ( .C (clk), .D (signal_18285), .Q (signal_18286) ) ;
    buf_clk cell_13404 ( .C (clk), .D (signal_18291), .Q (signal_18292) ) ;
    buf_clk cell_13410 ( .C (clk), .D (signal_18297), .Q (signal_18298) ) ;
    buf_clk cell_13416 ( .C (clk), .D (signal_18303), .Q (signal_18304) ) ;
    buf_clk cell_13422 ( .C (clk), .D (signal_18309), .Q (signal_18310) ) ;
    buf_clk cell_13428 ( .C (clk), .D (signal_18315), .Q (signal_18316) ) ;
    buf_clk cell_13434 ( .C (clk), .D (signal_18321), .Q (signal_18322) ) ;
    buf_clk cell_13440 ( .C (clk), .D (signal_18327), .Q (signal_18328) ) ;
    buf_clk cell_13446 ( .C (clk), .D (signal_18333), .Q (signal_18334) ) ;
    buf_clk cell_13452 ( .C (clk), .D (signal_18339), .Q (signal_18340) ) ;
    buf_clk cell_13458 ( .C (clk), .D (signal_18345), .Q (signal_18346) ) ;
    buf_clk cell_13464 ( .C (clk), .D (signal_18351), .Q (signal_18352) ) ;
    buf_clk cell_13470 ( .C (clk), .D (signal_18357), .Q (signal_18358) ) ;
    buf_clk cell_13476 ( .C (clk), .D (signal_18363), .Q (signal_18364) ) ;
    buf_clk cell_13482 ( .C (clk), .D (signal_18369), .Q (signal_18370) ) ;
    buf_clk cell_13488 ( .C (clk), .D (signal_18375), .Q (signal_18376) ) ;
    buf_clk cell_13494 ( .C (clk), .D (signal_18381), .Q (signal_18382) ) ;
    buf_clk cell_13500 ( .C (clk), .D (signal_18387), .Q (signal_18388) ) ;
    buf_clk cell_13506 ( .C (clk), .D (signal_18393), .Q (signal_18394) ) ;
    buf_clk cell_13512 ( .C (clk), .D (signal_18399), .Q (signal_18400) ) ;
    buf_clk cell_13518 ( .C (clk), .D (signal_18405), .Q (signal_18406) ) ;
    buf_clk cell_13524 ( .C (clk), .D (signal_18411), .Q (signal_18412) ) ;
    buf_clk cell_13530 ( .C (clk), .D (signal_18417), .Q (signal_18418) ) ;
    buf_clk cell_13536 ( .C (clk), .D (signal_18423), .Q (signal_18424) ) ;
    buf_clk cell_13542 ( .C (clk), .D (signal_18429), .Q (signal_18430) ) ;
    buf_clk cell_13548 ( .C (clk), .D (signal_18435), .Q (signal_18436) ) ;
    buf_clk cell_13554 ( .C (clk), .D (signal_18441), .Q (signal_18442) ) ;
    buf_clk cell_13560 ( .C (clk), .D (signal_18447), .Q (signal_18448) ) ;
    buf_clk cell_13566 ( .C (clk), .D (signal_18453), .Q (signal_18454) ) ;
    buf_clk cell_13572 ( .C (clk), .D (signal_18459), .Q (signal_18460) ) ;
    buf_clk cell_13578 ( .C (clk), .D (signal_18465), .Q (signal_18466) ) ;
    buf_clk cell_13584 ( .C (clk), .D (signal_18471), .Q (signal_18472) ) ;
    buf_clk cell_13590 ( .C (clk), .D (signal_18477), .Q (signal_18478) ) ;
    buf_clk cell_13596 ( .C (clk), .D (signal_18483), .Q (signal_18484) ) ;
    buf_clk cell_13602 ( .C (clk), .D (signal_18489), .Q (signal_18490) ) ;
    buf_clk cell_13608 ( .C (clk), .D (signal_18495), .Q (signal_18496) ) ;
    buf_clk cell_13614 ( .C (clk), .D (signal_18501), .Q (signal_18502) ) ;
    buf_clk cell_13620 ( .C (clk), .D (signal_18507), .Q (signal_18508) ) ;
    buf_clk cell_13626 ( .C (clk), .D (signal_18513), .Q (signal_18514) ) ;
    buf_clk cell_13632 ( .C (clk), .D (signal_18519), .Q (signal_18520) ) ;
    buf_clk cell_13638 ( .C (clk), .D (signal_18525), .Q (signal_18526) ) ;
    buf_clk cell_13644 ( .C (clk), .D (signal_18531), .Q (signal_18532) ) ;
    buf_clk cell_13650 ( .C (clk), .D (signal_18537), .Q (signal_18538) ) ;
    buf_clk cell_13656 ( .C (clk), .D (signal_18543), .Q (signal_18544) ) ;
    buf_clk cell_13662 ( .C (clk), .D (signal_18549), .Q (signal_18550) ) ;
    buf_clk cell_13668 ( .C (clk), .D (signal_18555), .Q (signal_18556) ) ;
    buf_clk cell_13674 ( .C (clk), .D (signal_18561), .Q (signal_18562) ) ;
    buf_clk cell_13680 ( .C (clk), .D (signal_18567), .Q (signal_18568) ) ;
    buf_clk cell_13686 ( .C (clk), .D (signal_18573), .Q (signal_18574) ) ;
    buf_clk cell_13692 ( .C (clk), .D (signal_18579), .Q (signal_18580) ) ;
    buf_clk cell_13698 ( .C (clk), .D (signal_18585), .Q (signal_18586) ) ;
    buf_clk cell_13704 ( .C (clk), .D (signal_18591), .Q (signal_18592) ) ;
    buf_clk cell_13710 ( .C (clk), .D (signal_18597), .Q (signal_18598) ) ;
    buf_clk cell_13716 ( .C (clk), .D (signal_18603), .Q (signal_18604) ) ;
    buf_clk cell_13722 ( .C (clk), .D (signal_18609), .Q (signal_18610) ) ;
    buf_clk cell_13728 ( .C (clk), .D (signal_18615), .Q (signal_18616) ) ;
    buf_clk cell_13734 ( .C (clk), .D (signal_18621), .Q (signal_18622) ) ;
    buf_clk cell_13740 ( .C (clk), .D (signal_18627), .Q (signal_18628) ) ;
    buf_clk cell_13746 ( .C (clk), .D (signal_18633), .Q (signal_18634) ) ;
    buf_clk cell_13752 ( .C (clk), .D (signal_18639), .Q (signal_18640) ) ;
    buf_clk cell_13758 ( .C (clk), .D (signal_18645), .Q (signal_18646) ) ;
    buf_clk cell_13764 ( .C (clk), .D (signal_18651), .Q (signal_18652) ) ;
    buf_clk cell_13770 ( .C (clk), .D (signal_18657), .Q (signal_18658) ) ;
    buf_clk cell_13776 ( .C (clk), .D (signal_18663), .Q (signal_18664) ) ;
    buf_clk cell_13782 ( .C (clk), .D (signal_18669), .Q (signal_18670) ) ;
    buf_clk cell_13788 ( .C (clk), .D (signal_18675), .Q (signal_18676) ) ;
    buf_clk cell_13794 ( .C (clk), .D (signal_18681), .Q (signal_18682) ) ;
    buf_clk cell_13800 ( .C (clk), .D (signal_18687), .Q (signal_18688) ) ;
    buf_clk cell_13806 ( .C (clk), .D (signal_18693), .Q (signal_18694) ) ;
    buf_clk cell_13812 ( .C (clk), .D (signal_18699), .Q (signal_18700) ) ;
    buf_clk cell_13818 ( .C (clk), .D (signal_18705), .Q (signal_18706) ) ;
    buf_clk cell_13824 ( .C (clk), .D (signal_18711), .Q (signal_18712) ) ;
    buf_clk cell_13830 ( .C (clk), .D (signal_18717), .Q (signal_18718) ) ;
    buf_clk cell_13836 ( .C (clk), .D (signal_18723), .Q (signal_18724) ) ;
    buf_clk cell_13842 ( .C (clk), .D (signal_18729), .Q (signal_18730) ) ;
    buf_clk cell_13848 ( .C (clk), .D (signal_18735), .Q (signal_18736) ) ;
    buf_clk cell_13854 ( .C (clk), .D (signal_18741), .Q (signal_18742) ) ;
    buf_clk cell_13860 ( .C (clk), .D (signal_18747), .Q (signal_18748) ) ;
    buf_clk cell_13866 ( .C (clk), .D (signal_18753), .Q (signal_18754) ) ;
    buf_clk cell_13872 ( .C (clk), .D (signal_18759), .Q (signal_18760) ) ;
    buf_clk cell_13878 ( .C (clk), .D (signal_18765), .Q (signal_18766) ) ;
    buf_clk cell_13884 ( .C (clk), .D (signal_18771), .Q (signal_18772) ) ;
    buf_clk cell_13890 ( .C (clk), .D (signal_18777), .Q (signal_18778) ) ;
    buf_clk cell_13896 ( .C (clk), .D (signal_18783), .Q (signal_18784) ) ;
    buf_clk cell_13902 ( .C (clk), .D (signal_18789), .Q (signal_18790) ) ;
    buf_clk cell_13908 ( .C (clk), .D (signal_18795), .Q (signal_18796) ) ;
    buf_clk cell_13914 ( .C (clk), .D (signal_18801), .Q (signal_18802) ) ;
    buf_clk cell_13920 ( .C (clk), .D (signal_18807), .Q (signal_18808) ) ;
    buf_clk cell_13926 ( .C (clk), .D (signal_18813), .Q (signal_18814) ) ;
    buf_clk cell_13932 ( .C (clk), .D (signal_18819), .Q (signal_18820) ) ;
    buf_clk cell_13938 ( .C (clk), .D (signal_18825), .Q (signal_18826) ) ;
    buf_clk cell_13944 ( .C (clk), .D (signal_18831), .Q (signal_18832) ) ;
    buf_clk cell_13950 ( .C (clk), .D (signal_18837), .Q (signal_18838) ) ;
    buf_clk cell_13956 ( .C (clk), .D (signal_18843), .Q (signal_18844) ) ;
    buf_clk cell_13962 ( .C (clk), .D (signal_18849), .Q (signal_18850) ) ;
    buf_clk cell_13968 ( .C (clk), .D (signal_18855), .Q (signal_18856) ) ;
    buf_clk cell_13974 ( .C (clk), .D (signal_18861), .Q (signal_18862) ) ;
    buf_clk cell_13980 ( .C (clk), .D (signal_18867), .Q (signal_18868) ) ;
    buf_clk cell_13986 ( .C (clk), .D (signal_18873), .Q (signal_18874) ) ;
    buf_clk cell_13992 ( .C (clk), .D (signal_18879), .Q (signal_18880) ) ;
    buf_clk cell_13998 ( .C (clk), .D (signal_18885), .Q (signal_18886) ) ;
    buf_clk cell_14004 ( .C (clk), .D (signal_18891), .Q (signal_18892) ) ;
    buf_clk cell_14010 ( .C (clk), .D (signal_18897), .Q (signal_18898) ) ;
    buf_clk cell_14016 ( .C (clk), .D (signal_18903), .Q (signal_18904) ) ;
    buf_clk cell_14022 ( .C (clk), .D (signal_18909), .Q (signal_18910) ) ;
    buf_clk cell_14028 ( .C (clk), .D (signal_18915), .Q (signal_18916) ) ;
    buf_clk cell_14034 ( .C (clk), .D (signal_18921), .Q (signal_18922) ) ;
    buf_clk cell_14040 ( .C (clk), .D (signal_18927), .Q (signal_18928) ) ;
    buf_clk cell_14046 ( .C (clk), .D (signal_18933), .Q (signal_18934) ) ;
    buf_clk cell_14052 ( .C (clk), .D (signal_18939), .Q (signal_18940) ) ;
    buf_clk cell_14058 ( .C (clk), .D (signal_18945), .Q (signal_18946) ) ;
    buf_clk cell_14064 ( .C (clk), .D (signal_18951), .Q (signal_18952) ) ;
    buf_clk cell_14070 ( .C (clk), .D (signal_18957), .Q (signal_18958) ) ;
    buf_clk cell_14076 ( .C (clk), .D (signal_18963), .Q (signal_18964) ) ;
    buf_clk cell_14082 ( .C (clk), .D (signal_18969), .Q (signal_18970) ) ;
    buf_clk cell_14088 ( .C (clk), .D (signal_18975), .Q (signal_18976) ) ;
    buf_clk cell_14094 ( .C (clk), .D (signal_18981), .Q (signal_18982) ) ;
    buf_clk cell_14100 ( .C (clk), .D (signal_18987), .Q (signal_18988) ) ;
    buf_clk cell_14106 ( .C (clk), .D (signal_18993), .Q (signal_18994) ) ;
    buf_clk cell_14112 ( .C (clk), .D (signal_18999), .Q (signal_19000) ) ;
    buf_clk cell_14118 ( .C (clk), .D (signal_19005), .Q (signal_19006) ) ;
    buf_clk cell_14124 ( .C (clk), .D (signal_19011), .Q (signal_19012) ) ;
    buf_clk cell_14130 ( .C (clk), .D (signal_19017), .Q (signal_19018) ) ;
    buf_clk cell_14136 ( .C (clk), .D (signal_19023), .Q (signal_19024) ) ;
    buf_clk cell_14142 ( .C (clk), .D (signal_19029), .Q (signal_19030) ) ;
    buf_clk cell_14148 ( .C (clk), .D (signal_19035), .Q (signal_19036) ) ;
    buf_clk cell_14154 ( .C (clk), .D (signal_19041), .Q (signal_19042) ) ;
    buf_clk cell_14160 ( .C (clk), .D (signal_19047), .Q (signal_19048) ) ;
    buf_clk cell_14166 ( .C (clk), .D (signal_19053), .Q (signal_19054) ) ;
    buf_clk cell_14172 ( .C (clk), .D (signal_19059), .Q (signal_19060) ) ;
    buf_clk cell_14178 ( .C (clk), .D (signal_19065), .Q (signal_19066) ) ;
    buf_clk cell_14184 ( .C (clk), .D (signal_19071), .Q (signal_19072) ) ;
    buf_clk cell_14190 ( .C (clk), .D (signal_19077), .Q (signal_19078) ) ;
    buf_clk cell_14196 ( .C (clk), .D (signal_19083), .Q (signal_19084) ) ;
    buf_clk cell_14202 ( .C (clk), .D (signal_19089), .Q (signal_19090) ) ;
    buf_clk cell_14208 ( .C (clk), .D (signal_19095), .Q (signal_19096) ) ;
    buf_clk cell_14214 ( .C (clk), .D (signal_19101), .Q (signal_19102) ) ;
    buf_clk cell_14220 ( .C (clk), .D (signal_19107), .Q (signal_19108) ) ;
    buf_clk cell_14226 ( .C (clk), .D (signal_19113), .Q (signal_19114) ) ;
    buf_clk cell_14232 ( .C (clk), .D (signal_19119), .Q (signal_19120) ) ;
    buf_clk cell_14238 ( .C (clk), .D (signal_19125), .Q (signal_19126) ) ;
    buf_clk cell_14244 ( .C (clk), .D (signal_19131), .Q (signal_19132) ) ;
    buf_clk cell_14250 ( .C (clk), .D (signal_19137), .Q (signal_19138) ) ;
    buf_clk cell_14256 ( .C (clk), .D (signal_19143), .Q (signal_19144) ) ;
    buf_clk cell_14262 ( .C (clk), .D (signal_19149), .Q (signal_19150) ) ;
    buf_clk cell_14268 ( .C (clk), .D (signal_19155), .Q (signal_19156) ) ;
    buf_clk cell_14274 ( .C (clk), .D (signal_19161), .Q (signal_19162) ) ;
    buf_clk cell_14280 ( .C (clk), .D (signal_19167), .Q (signal_19168) ) ;
    buf_clk cell_14286 ( .C (clk), .D (signal_19173), .Q (signal_19174) ) ;
    buf_clk cell_14292 ( .C (clk), .D (signal_19179), .Q (signal_19180) ) ;
    buf_clk cell_14298 ( .C (clk), .D (signal_19185), .Q (signal_19186) ) ;
    buf_clk cell_14304 ( .C (clk), .D (signal_19191), .Q (signal_19192) ) ;
    buf_clk cell_14310 ( .C (clk), .D (signal_19197), .Q (signal_19198) ) ;
    buf_clk cell_14316 ( .C (clk), .D (signal_19203), .Q (signal_19204) ) ;
    buf_clk cell_14322 ( .C (clk), .D (signal_19209), .Q (signal_19210) ) ;
    buf_clk cell_14328 ( .C (clk), .D (signal_19215), .Q (signal_19216) ) ;
    buf_clk cell_14334 ( .C (clk), .D (signal_19221), .Q (signal_19222) ) ;
    buf_clk cell_14340 ( .C (clk), .D (signal_19227), .Q (signal_19228) ) ;
    buf_clk cell_14346 ( .C (clk), .D (signal_19233), .Q (signal_19234) ) ;
    buf_clk cell_14352 ( .C (clk), .D (signal_19239), .Q (signal_19240) ) ;
    buf_clk cell_14358 ( .C (clk), .D (signal_19245), .Q (signal_19246) ) ;
    buf_clk cell_14364 ( .C (clk), .D (signal_19251), .Q (signal_19252) ) ;
    buf_clk cell_14370 ( .C (clk), .D (signal_19257), .Q (signal_19258) ) ;
    buf_clk cell_14376 ( .C (clk), .D (signal_19263), .Q (signal_19264) ) ;
    buf_clk cell_14382 ( .C (clk), .D (signal_19269), .Q (signal_19270) ) ;
    buf_clk cell_14388 ( .C (clk), .D (signal_19275), .Q (signal_19276) ) ;
    buf_clk cell_14394 ( .C (clk), .D (signal_19281), .Q (signal_19282) ) ;
    buf_clk cell_14400 ( .C (clk), .D (signal_19287), .Q (signal_19288) ) ;
    buf_clk cell_14406 ( .C (clk), .D (signal_19293), .Q (signal_19294) ) ;
    buf_clk cell_14412 ( .C (clk), .D (signal_19299), .Q (signal_19300) ) ;
    buf_clk cell_14418 ( .C (clk), .D (signal_19305), .Q (signal_19306) ) ;
    buf_clk cell_14424 ( .C (clk), .D (signal_19311), .Q (signal_19312) ) ;
    buf_clk cell_14430 ( .C (clk), .D (signal_19317), .Q (signal_19318) ) ;
    buf_clk cell_14436 ( .C (clk), .D (signal_19323), .Q (signal_19324) ) ;
    buf_clk cell_14442 ( .C (clk), .D (signal_19329), .Q (signal_19330) ) ;
    buf_clk cell_14448 ( .C (clk), .D (signal_19335), .Q (signal_19336) ) ;
    buf_clk cell_14454 ( .C (clk), .D (signal_19341), .Q (signal_19342) ) ;
    buf_clk cell_14460 ( .C (clk), .D (signal_19347), .Q (signal_19348) ) ;
    buf_clk cell_14466 ( .C (clk), .D (signal_19353), .Q (signal_19354) ) ;
    buf_clk cell_14472 ( .C (clk), .D (signal_19359), .Q (signal_19360) ) ;
    buf_clk cell_14478 ( .C (clk), .D (signal_19365), .Q (signal_19366) ) ;
    buf_clk cell_14484 ( .C (clk), .D (signal_19371), .Q (signal_19372) ) ;
    buf_clk cell_14490 ( .C (clk), .D (signal_19377), .Q (signal_19378) ) ;
    buf_clk cell_14496 ( .C (clk), .D (signal_19383), .Q (signal_19384) ) ;
    buf_clk cell_14502 ( .C (clk), .D (signal_19389), .Q (signal_19390) ) ;
    buf_clk cell_14508 ( .C (clk), .D (signal_19395), .Q (signal_19396) ) ;
    buf_clk cell_14514 ( .C (clk), .D (signal_19401), .Q (signal_19402) ) ;
    buf_clk cell_14520 ( .C (clk), .D (signal_19407), .Q (signal_19408) ) ;
    buf_clk cell_14526 ( .C (clk), .D (signal_19413), .Q (signal_19414) ) ;
    buf_clk cell_14532 ( .C (clk), .D (signal_19419), .Q (signal_19420) ) ;
    buf_clk cell_14538 ( .C (clk), .D (signal_19425), .Q (signal_19426) ) ;
    buf_clk cell_14544 ( .C (clk), .D (signal_19431), .Q (signal_19432) ) ;
    buf_clk cell_14550 ( .C (clk), .D (signal_19437), .Q (signal_19438) ) ;
    buf_clk cell_14556 ( .C (clk), .D (signal_19443), .Q (signal_19444) ) ;
    buf_clk cell_14562 ( .C (clk), .D (signal_19449), .Q (signal_19450) ) ;
    buf_clk cell_14568 ( .C (clk), .D (signal_19455), .Q (signal_19456) ) ;
    buf_clk cell_14574 ( .C (clk), .D (signal_19461), .Q (signal_19462) ) ;
    buf_clk cell_14580 ( .C (clk), .D (signal_19467), .Q (signal_19468) ) ;
    buf_clk cell_14586 ( .C (clk), .D (signal_19473), .Q (signal_19474) ) ;
    buf_clk cell_14592 ( .C (clk), .D (signal_19479), .Q (signal_19480) ) ;
    buf_clk cell_14598 ( .C (clk), .D (signal_19485), .Q (signal_19486) ) ;
    buf_clk cell_14604 ( .C (clk), .D (signal_19491), .Q (signal_19492) ) ;
    buf_clk cell_14610 ( .C (clk), .D (signal_19497), .Q (signal_19498) ) ;
    buf_clk cell_14616 ( .C (clk), .D (signal_19503), .Q (signal_19504) ) ;
    buf_clk cell_14622 ( .C (clk), .D (signal_19509), .Q (signal_19510) ) ;
    buf_clk cell_14628 ( .C (clk), .D (signal_19515), .Q (signal_19516) ) ;
    buf_clk cell_14634 ( .C (clk), .D (signal_19521), .Q (signal_19522) ) ;
    buf_clk cell_14640 ( .C (clk), .D (signal_19527), .Q (signal_19528) ) ;
    buf_clk cell_14646 ( .C (clk), .D (signal_19533), .Q (signal_19534) ) ;
    buf_clk cell_14652 ( .C (clk), .D (signal_19539), .Q (signal_19540) ) ;
    buf_clk cell_14658 ( .C (clk), .D (signal_19545), .Q (signal_19546) ) ;
    buf_clk cell_14664 ( .C (clk), .D (signal_19551), .Q (signal_19552) ) ;
    buf_clk cell_14670 ( .C (clk), .D (signal_19557), .Q (signal_19558) ) ;
    buf_clk cell_14676 ( .C (clk), .D (signal_19563), .Q (signal_19564) ) ;
    buf_clk cell_14682 ( .C (clk), .D (signal_19569), .Q (signal_19570) ) ;
    buf_clk cell_14688 ( .C (clk), .D (signal_19575), .Q (signal_19576) ) ;
    buf_clk cell_14694 ( .C (clk), .D (signal_19581), .Q (signal_19582) ) ;
    buf_clk cell_14700 ( .C (clk), .D (signal_19587), .Q (signal_19588) ) ;
    buf_clk cell_14706 ( .C (clk), .D (signal_19593), .Q (signal_19594) ) ;
    buf_clk cell_14712 ( .C (clk), .D (signal_19599), .Q (signal_19600) ) ;
    buf_clk cell_14718 ( .C (clk), .D (signal_19605), .Q (signal_19606) ) ;
    buf_clk cell_14724 ( .C (clk), .D (signal_19611), .Q (signal_19612) ) ;
    buf_clk cell_14730 ( .C (clk), .D (signal_19617), .Q (signal_19618) ) ;
    buf_clk cell_14736 ( .C (clk), .D (signal_19623), .Q (signal_19624) ) ;
    buf_clk cell_14742 ( .C (clk), .D (signal_19629), .Q (signal_19630) ) ;
    buf_clk cell_14748 ( .C (clk), .D (signal_19635), .Q (signal_19636) ) ;
    buf_clk cell_14754 ( .C (clk), .D (signal_19641), .Q (signal_19642) ) ;
    buf_clk cell_14760 ( .C (clk), .D (signal_19647), .Q (signal_19648) ) ;
    buf_clk cell_14766 ( .C (clk), .D (signal_19653), .Q (signal_19654) ) ;
    buf_clk cell_14772 ( .C (clk), .D (signal_19659), .Q (signal_19660) ) ;
    buf_clk cell_14778 ( .C (clk), .D (signal_19665), .Q (signal_19666) ) ;
    buf_clk cell_14784 ( .C (clk), .D (signal_19671), .Q (signal_19672) ) ;
    buf_clk cell_14790 ( .C (clk), .D (signal_19677), .Q (signal_19678) ) ;
    buf_clk cell_14796 ( .C (clk), .D (signal_19683), .Q (signal_19684) ) ;
    buf_clk cell_14802 ( .C (clk), .D (signal_19689), .Q (signal_19690) ) ;
    buf_clk cell_14808 ( .C (clk), .D (signal_19695), .Q (signal_19696) ) ;
    buf_clk cell_14814 ( .C (clk), .D (signal_19701), .Q (signal_19702) ) ;
    buf_clk cell_14820 ( .C (clk), .D (signal_19707), .Q (signal_19708) ) ;
    buf_clk cell_14826 ( .C (clk), .D (signal_19713), .Q (signal_19714) ) ;
    buf_clk cell_14832 ( .C (clk), .D (signal_19719), .Q (signal_19720) ) ;
    buf_clk cell_14838 ( .C (clk), .D (signal_19725), .Q (signal_19726) ) ;
    buf_clk cell_14844 ( .C (clk), .D (signal_19731), .Q (signal_19732) ) ;
    buf_clk cell_14850 ( .C (clk), .D (signal_19737), .Q (signal_19738) ) ;
    buf_clk cell_14856 ( .C (clk), .D (signal_19743), .Q (signal_19744) ) ;
    buf_clk cell_14862 ( .C (clk), .D (signal_19749), .Q (signal_19750) ) ;
    buf_clk cell_14868 ( .C (clk), .D (signal_19755), .Q (signal_19756) ) ;
    buf_clk cell_14874 ( .C (clk), .D (signal_19761), .Q (signal_19762) ) ;
    buf_clk cell_14880 ( .C (clk), .D (signal_19767), .Q (signal_19768) ) ;
    buf_clk cell_14886 ( .C (clk), .D (signal_19773), .Q (signal_19774) ) ;
    buf_clk cell_14892 ( .C (clk), .D (signal_19779), .Q (signal_19780) ) ;
    buf_clk cell_14898 ( .C (clk), .D (signal_19785), .Q (signal_19786) ) ;
    buf_clk cell_14904 ( .C (clk), .D (signal_19791), .Q (signal_19792) ) ;
    buf_clk cell_14910 ( .C (clk), .D (signal_19797), .Q (signal_19798) ) ;
    buf_clk cell_14916 ( .C (clk), .D (signal_19803), .Q (signal_19804) ) ;
    buf_clk cell_14922 ( .C (clk), .D (signal_19809), .Q (signal_19810) ) ;
    buf_clk cell_14928 ( .C (clk), .D (signal_19815), .Q (signal_19816) ) ;
    buf_clk cell_14934 ( .C (clk), .D (signal_19821), .Q (signal_19822) ) ;
    buf_clk cell_14940 ( .C (clk), .D (signal_19827), .Q (signal_19828) ) ;
    buf_clk cell_14946 ( .C (clk), .D (signal_19833), .Q (signal_19834) ) ;
    buf_clk cell_14952 ( .C (clk), .D (signal_19839), .Q (signal_19840) ) ;
    buf_clk cell_14958 ( .C (clk), .D (signal_19845), .Q (signal_19846) ) ;
    buf_clk cell_14964 ( .C (clk), .D (signal_19851), .Q (signal_19852) ) ;
    buf_clk cell_14970 ( .C (clk), .D (signal_19857), .Q (signal_19858) ) ;
    buf_clk cell_14976 ( .C (clk), .D (signal_19863), .Q (signal_19864) ) ;
    buf_clk cell_14982 ( .C (clk), .D (signal_19869), .Q (signal_19870) ) ;
    buf_clk cell_14988 ( .C (clk), .D (signal_19875), .Q (signal_19876) ) ;
    buf_clk cell_14994 ( .C (clk), .D (signal_19881), .Q (signal_19882) ) ;
    buf_clk cell_15000 ( .C (clk), .D (signal_19887), .Q (signal_19888) ) ;
    buf_clk cell_15006 ( .C (clk), .D (signal_19893), .Q (signal_19894) ) ;
    buf_clk cell_15012 ( .C (clk), .D (signal_19899), .Q (signal_19900) ) ;
    buf_clk cell_15018 ( .C (clk), .D (signal_19905), .Q (signal_19906) ) ;
    buf_clk cell_15024 ( .C (clk), .D (signal_19911), .Q (signal_19912) ) ;
    buf_clk cell_15030 ( .C (clk), .D (signal_19917), .Q (signal_19918) ) ;
    buf_clk cell_15036 ( .C (clk), .D (signal_19923), .Q (signal_19924) ) ;
    buf_clk cell_15042 ( .C (clk), .D (signal_19929), .Q (signal_19930) ) ;
    buf_clk cell_15048 ( .C (clk), .D (signal_19935), .Q (signal_19936) ) ;
    buf_clk cell_15054 ( .C (clk), .D (signal_19941), .Q (signal_19942) ) ;
    buf_clk cell_15060 ( .C (clk), .D (signal_19947), .Q (signal_19948) ) ;
    buf_clk cell_15066 ( .C (clk), .D (signal_19953), .Q (signal_19954) ) ;
    buf_clk cell_15072 ( .C (clk), .D (signal_19959), .Q (signal_19960) ) ;
    buf_clk cell_15078 ( .C (clk), .D (signal_19965), .Q (signal_19966) ) ;
    buf_clk cell_15084 ( .C (clk), .D (signal_19971), .Q (signal_19972) ) ;
    buf_clk cell_15090 ( .C (clk), .D (signal_19977), .Q (signal_19978) ) ;
    buf_clk cell_15096 ( .C (clk), .D (signal_19983), .Q (signal_19984) ) ;
    buf_clk cell_15102 ( .C (clk), .D (signal_19989), .Q (signal_19990) ) ;
    buf_clk cell_15108 ( .C (clk), .D (signal_19995), .Q (signal_19996) ) ;
    buf_clk cell_15114 ( .C (clk), .D (signal_20001), .Q (signal_20002) ) ;
    buf_clk cell_15120 ( .C (clk), .D (signal_20007), .Q (signal_20008) ) ;
    buf_clk cell_15126 ( .C (clk), .D (signal_20013), .Q (signal_20014) ) ;
    buf_clk cell_15132 ( .C (clk), .D (signal_20019), .Q (signal_20020) ) ;
    buf_clk cell_15138 ( .C (clk), .D (signal_20025), .Q (signal_20026) ) ;
    buf_clk cell_15144 ( .C (clk), .D (signal_20031), .Q (signal_20032) ) ;
    buf_clk cell_15150 ( .C (clk), .D (signal_20037), .Q (signal_20038) ) ;
    buf_clk cell_15156 ( .C (clk), .D (signal_20043), .Q (signal_20044) ) ;
    buf_clk cell_15162 ( .C (clk), .D (signal_20049), .Q (signal_20050) ) ;
    buf_clk cell_15168 ( .C (clk), .D (signal_20055), .Q (signal_20056) ) ;
    buf_clk cell_15174 ( .C (clk), .D (signal_20061), .Q (signal_20062) ) ;
    buf_clk cell_15180 ( .C (clk), .D (signal_20067), .Q (signal_20068) ) ;
    buf_clk cell_15186 ( .C (clk), .D (signal_20073), .Q (signal_20074) ) ;
    buf_clk cell_15192 ( .C (clk), .D (signal_20079), .Q (signal_20080) ) ;
    buf_clk cell_15198 ( .C (clk), .D (signal_20085), .Q (signal_20086) ) ;
    buf_clk cell_15204 ( .C (clk), .D (signal_20091), .Q (signal_20092) ) ;
    buf_clk cell_15210 ( .C (clk), .D (signal_20097), .Q (signal_20098) ) ;
    buf_clk cell_15216 ( .C (clk), .D (signal_20103), .Q (signal_20104) ) ;
    buf_clk cell_15222 ( .C (clk), .D (signal_20109), .Q (signal_20110) ) ;
    buf_clk cell_15228 ( .C (clk), .D (signal_20115), .Q (signal_20116) ) ;
    buf_clk cell_15234 ( .C (clk), .D (signal_20121), .Q (signal_20122) ) ;
    buf_clk cell_15240 ( .C (clk), .D (signal_20127), .Q (signal_20128) ) ;
    buf_clk cell_15246 ( .C (clk), .D (signal_20133), .Q (signal_20134) ) ;
    buf_clk cell_15252 ( .C (clk), .D (signal_20139), .Q (signal_20140) ) ;
    buf_clk cell_15258 ( .C (clk), .D (signal_20145), .Q (signal_20146) ) ;
    buf_clk cell_15264 ( .C (clk), .D (signal_20151), .Q (signal_20152) ) ;
    buf_clk cell_15270 ( .C (clk), .D (signal_20157), .Q (signal_20158) ) ;
    buf_clk cell_15276 ( .C (clk), .D (signal_20163), .Q (signal_20164) ) ;
    buf_clk cell_15282 ( .C (clk), .D (signal_20169), .Q (signal_20170) ) ;
    buf_clk cell_15288 ( .C (clk), .D (signal_20175), .Q (signal_20176) ) ;
    buf_clk cell_15294 ( .C (clk), .D (signal_20181), .Q (signal_20182) ) ;
    buf_clk cell_15300 ( .C (clk), .D (signal_20187), .Q (signal_20188) ) ;
    buf_clk cell_15306 ( .C (clk), .D (signal_20193), .Q (signal_20194) ) ;
    buf_clk cell_15312 ( .C (clk), .D (signal_20199), .Q (signal_20200) ) ;
    buf_clk cell_15318 ( .C (clk), .D (signal_20205), .Q (signal_20206) ) ;
    buf_clk cell_15324 ( .C (clk), .D (signal_20211), .Q (signal_20212) ) ;
    buf_clk cell_15330 ( .C (clk), .D (signal_20217), .Q (signal_20218) ) ;
    buf_clk cell_15336 ( .C (clk), .D (signal_20223), .Q (signal_20224) ) ;
    buf_clk cell_15342 ( .C (clk), .D (signal_20229), .Q (signal_20230) ) ;
    buf_clk cell_15348 ( .C (clk), .D (signal_20235), .Q (signal_20236) ) ;
    buf_clk cell_15354 ( .C (clk), .D (signal_20241), .Q (signal_20242) ) ;
    buf_clk cell_15360 ( .C (clk), .D (signal_20247), .Q (signal_20248) ) ;
    buf_clk cell_15366 ( .C (clk), .D (signal_20253), .Q (signal_20254) ) ;
    buf_clk cell_15372 ( .C (clk), .D (signal_20259), .Q (signal_20260) ) ;
    buf_clk cell_15378 ( .C (clk), .D (signal_20265), .Q (signal_20266) ) ;
    buf_clk cell_15384 ( .C (clk), .D (signal_20271), .Q (signal_20272) ) ;
    buf_clk cell_15390 ( .C (clk), .D (signal_20277), .Q (signal_20278) ) ;
    buf_clk cell_15396 ( .C (clk), .D (signal_20283), .Q (signal_20284) ) ;
    buf_clk cell_15402 ( .C (clk), .D (signal_20289), .Q (signal_20290) ) ;
    buf_clk cell_15408 ( .C (clk), .D (signal_20295), .Q (signal_20296) ) ;
    buf_clk cell_15414 ( .C (clk), .D (signal_20301), .Q (signal_20302) ) ;
    buf_clk cell_15420 ( .C (clk), .D (signal_20307), .Q (signal_20308) ) ;
    buf_clk cell_15426 ( .C (clk), .D (signal_20313), .Q (signal_20314) ) ;
    buf_clk cell_15432 ( .C (clk), .D (signal_20319), .Q (signal_20320) ) ;
    buf_clk cell_15438 ( .C (clk), .D (signal_20325), .Q (signal_20326) ) ;
    buf_clk cell_15444 ( .C (clk), .D (signal_20331), .Q (signal_20332) ) ;
    buf_clk cell_15450 ( .C (clk), .D (signal_20337), .Q (signal_20338) ) ;
    buf_clk cell_15456 ( .C (clk), .D (signal_20343), .Q (signal_20344) ) ;
    buf_clk cell_15462 ( .C (clk), .D (signal_20349), .Q (signal_20350) ) ;
    buf_clk cell_15468 ( .C (clk), .D (signal_20355), .Q (signal_20356) ) ;
    buf_clk cell_15474 ( .C (clk), .D (signal_20361), .Q (signal_20362) ) ;
    buf_clk cell_15480 ( .C (clk), .D (signal_20367), .Q (signal_20368) ) ;
    buf_clk cell_15486 ( .C (clk), .D (signal_20373), .Q (signal_20374) ) ;
    buf_clk cell_15492 ( .C (clk), .D (signal_20379), .Q (signal_20380) ) ;
    buf_clk cell_15498 ( .C (clk), .D (signal_20385), .Q (signal_20386) ) ;
    buf_clk cell_15504 ( .C (clk), .D (signal_20391), .Q (signal_20392) ) ;
    buf_clk cell_15510 ( .C (clk), .D (signal_20397), .Q (signal_20398) ) ;
    buf_clk cell_15516 ( .C (clk), .D (signal_20403), .Q (signal_20404) ) ;
    buf_clk cell_15522 ( .C (clk), .D (signal_20409), .Q (signal_20410) ) ;
    buf_clk cell_15528 ( .C (clk), .D (signal_20415), .Q (signal_20416) ) ;
    buf_clk cell_15534 ( .C (clk), .D (signal_20421), .Q (signal_20422) ) ;
    buf_clk cell_15540 ( .C (clk), .D (signal_20427), .Q (signal_20428) ) ;
    buf_clk cell_15546 ( .C (clk), .D (signal_20433), .Q (signal_20434) ) ;
    buf_clk cell_15552 ( .C (clk), .D (signal_20439), .Q (signal_20440) ) ;
    buf_clk cell_15558 ( .C (clk), .D (signal_20445), .Q (signal_20446) ) ;
    buf_clk cell_15564 ( .C (clk), .D (signal_20451), .Q (signal_20452) ) ;
    buf_clk cell_15570 ( .C (clk), .D (signal_20457), .Q (signal_20458) ) ;
    buf_clk cell_15576 ( .C (clk), .D (signal_20463), .Q (signal_20464) ) ;
    buf_clk cell_15582 ( .C (clk), .D (signal_20469), .Q (signal_20470) ) ;
    buf_clk cell_15588 ( .C (clk), .D (signal_20475), .Q (signal_20476) ) ;
    buf_clk cell_15594 ( .C (clk), .D (signal_20481), .Q (signal_20482) ) ;
    buf_clk cell_15600 ( .C (clk), .D (signal_20487), .Q (signal_20488) ) ;
    buf_clk cell_15606 ( .C (clk), .D (signal_20493), .Q (signal_20494) ) ;
    buf_clk cell_15612 ( .C (clk), .D (signal_20499), .Q (signal_20500) ) ;
    buf_clk cell_15618 ( .C (clk), .D (signal_20505), .Q (signal_20506) ) ;
    buf_clk cell_15624 ( .C (clk), .D (signal_20511), .Q (signal_20512) ) ;
    buf_clk cell_15630 ( .C (clk), .D (signal_20517), .Q (signal_20518) ) ;
    buf_clk cell_15636 ( .C (clk), .D (signal_20523), .Q (signal_20524) ) ;
    buf_clk cell_15642 ( .C (clk), .D (signal_20529), .Q (signal_20530) ) ;
    buf_clk cell_15648 ( .C (clk), .D (signal_20535), .Q (signal_20536) ) ;
    buf_clk cell_15654 ( .C (clk), .D (signal_20541), .Q (signal_20542) ) ;
    buf_clk cell_15660 ( .C (clk), .D (signal_20547), .Q (signal_20548) ) ;
    buf_clk cell_15666 ( .C (clk), .D (signal_20553), .Q (signal_20554) ) ;
    buf_clk cell_15672 ( .C (clk), .D (signal_20559), .Q (signal_20560) ) ;
    buf_clk cell_15678 ( .C (clk), .D (signal_20565), .Q (signal_20566) ) ;
    buf_clk cell_15684 ( .C (clk), .D (signal_20571), .Q (signal_20572) ) ;
    buf_clk cell_15690 ( .C (clk), .D (signal_20577), .Q (signal_20578) ) ;
    buf_clk cell_15696 ( .C (clk), .D (signal_20583), .Q (signal_20584) ) ;
    buf_clk cell_15702 ( .C (clk), .D (signal_20589), .Q (signal_20590) ) ;
    buf_clk cell_15708 ( .C (clk), .D (signal_20595), .Q (signal_20596) ) ;
    buf_clk cell_15714 ( .C (clk), .D (signal_20601), .Q (signal_20602) ) ;
    buf_clk cell_15720 ( .C (clk), .D (signal_20607), .Q (signal_20608) ) ;
    buf_clk cell_15726 ( .C (clk), .D (signal_20613), .Q (signal_20614) ) ;
    buf_clk cell_15732 ( .C (clk), .D (signal_20619), .Q (signal_20620) ) ;
    buf_clk cell_15738 ( .C (clk), .D (signal_20625), .Q (signal_20626) ) ;
    buf_clk cell_15744 ( .C (clk), .D (signal_20631), .Q (signal_20632) ) ;
    buf_clk cell_15750 ( .C (clk), .D (signal_20637), .Q (signal_20638) ) ;
    buf_clk cell_15756 ( .C (clk), .D (signal_20643), .Q (signal_20644) ) ;
    buf_clk cell_15762 ( .C (clk), .D (signal_20649), .Q (signal_20650) ) ;
    buf_clk cell_15768 ( .C (clk), .D (signal_20655), .Q (signal_20656) ) ;
    buf_clk cell_15774 ( .C (clk), .D (signal_20661), .Q (signal_20662) ) ;
    buf_clk cell_15780 ( .C (clk), .D (signal_20667), .Q (signal_20668) ) ;
    buf_clk cell_15786 ( .C (clk), .D (signal_20673), .Q (signal_20674) ) ;
    buf_clk cell_15792 ( .C (clk), .D (signal_20679), .Q (signal_20680) ) ;
    buf_clk cell_15798 ( .C (clk), .D (signal_20685), .Q (signal_20686) ) ;
    buf_clk cell_15804 ( .C (clk), .D (signal_20691), .Q (signal_20692) ) ;
    buf_clk cell_15810 ( .C (clk), .D (signal_20697), .Q (signal_20698) ) ;
    buf_clk cell_15816 ( .C (clk), .D (signal_20703), .Q (signal_20704) ) ;
    buf_clk cell_15822 ( .C (clk), .D (signal_20709), .Q (signal_20710) ) ;
    buf_clk cell_15828 ( .C (clk), .D (signal_20715), .Q (signal_20716) ) ;
    buf_clk cell_15834 ( .C (clk), .D (signal_20721), .Q (signal_20722) ) ;
    buf_clk cell_15840 ( .C (clk), .D (signal_20727), .Q (signal_20728) ) ;
    buf_clk cell_15846 ( .C (clk), .D (signal_20733), .Q (signal_20734) ) ;
    buf_clk cell_15852 ( .C (clk), .D (signal_20739), .Q (signal_20740) ) ;
    buf_clk cell_15858 ( .C (clk), .D (signal_20745), .Q (signal_20746) ) ;
    buf_clk cell_15864 ( .C (clk), .D (signal_20751), .Q (signal_20752) ) ;
    buf_clk cell_15870 ( .C (clk), .D (signal_20757), .Q (signal_20758) ) ;
    buf_clk cell_15876 ( .C (clk), .D (signal_20763), .Q (signal_20764) ) ;
    buf_clk cell_15882 ( .C (clk), .D (signal_20769), .Q (signal_20770) ) ;
    buf_clk cell_15888 ( .C (clk), .D (signal_20775), .Q (signal_20776) ) ;
    buf_clk cell_15894 ( .C (clk), .D (signal_20781), .Q (signal_20782) ) ;
    buf_clk cell_15900 ( .C (clk), .D (signal_20787), .Q (signal_20788) ) ;
    buf_clk cell_15906 ( .C (clk), .D (signal_20793), .Q (signal_20794) ) ;
    buf_clk cell_15912 ( .C (clk), .D (signal_20799), .Q (signal_20800) ) ;
    buf_clk cell_15918 ( .C (clk), .D (signal_20805), .Q (signal_20806) ) ;
    buf_clk cell_15924 ( .C (clk), .D (signal_20811), .Q (signal_20812) ) ;
    buf_clk cell_15930 ( .C (clk), .D (signal_20817), .Q (signal_20818) ) ;
    buf_clk cell_15936 ( .C (clk), .D (signal_20823), .Q (signal_20824) ) ;
    buf_clk cell_15942 ( .C (clk), .D (signal_20829), .Q (signal_20830) ) ;
    buf_clk cell_15948 ( .C (clk), .D (signal_20835), .Q (signal_20836) ) ;
    buf_clk cell_15954 ( .C (clk), .D (signal_20841), .Q (signal_20842) ) ;
    buf_clk cell_15960 ( .C (clk), .D (signal_20847), .Q (signal_20848) ) ;
    buf_clk cell_15966 ( .C (clk), .D (signal_20853), .Q (signal_20854) ) ;
    buf_clk cell_15972 ( .C (clk), .D (signal_20859), .Q (signal_20860) ) ;
    buf_clk cell_15978 ( .C (clk), .D (signal_20865), .Q (signal_20866) ) ;
    buf_clk cell_15984 ( .C (clk), .D (signal_20871), .Q (signal_20872) ) ;
    buf_clk cell_15990 ( .C (clk), .D (signal_20877), .Q (signal_20878) ) ;
    buf_clk cell_15996 ( .C (clk), .D (signal_20883), .Q (signal_20884) ) ;
    buf_clk cell_16002 ( .C (clk), .D (signal_20889), .Q (signal_20890) ) ;
    buf_clk cell_16008 ( .C (clk), .D (signal_20895), .Q (signal_20896) ) ;
    buf_clk cell_16014 ( .C (clk), .D (signal_20901), .Q (signal_20902) ) ;
    buf_clk cell_16020 ( .C (clk), .D (signal_20907), .Q (signal_20908) ) ;
    buf_clk cell_16026 ( .C (clk), .D (signal_20913), .Q (signal_20914) ) ;
    buf_clk cell_16032 ( .C (clk), .D (signal_20919), .Q (signal_20920) ) ;
    buf_clk cell_16038 ( .C (clk), .D (signal_20925), .Q (signal_20926) ) ;
    buf_clk cell_16044 ( .C (clk), .D (signal_20931), .Q (signal_20932) ) ;
    buf_clk cell_16050 ( .C (clk), .D (signal_20937), .Q (signal_20938) ) ;
    buf_clk cell_16056 ( .C (clk), .D (signal_20943), .Q (signal_20944) ) ;
    buf_clk cell_16062 ( .C (clk), .D (signal_20949), .Q (signal_20950) ) ;
    buf_clk cell_16068 ( .C (clk), .D (signal_20955), .Q (signal_20956) ) ;
    buf_clk cell_16074 ( .C (clk), .D (signal_20961), .Q (signal_20962) ) ;
    buf_clk cell_16080 ( .C (clk), .D (signal_20967), .Q (signal_20968) ) ;
    buf_clk cell_16086 ( .C (clk), .D (signal_20973), .Q (signal_20974) ) ;
    buf_clk cell_16092 ( .C (clk), .D (signal_20979), .Q (signal_20980) ) ;
    buf_clk cell_16098 ( .C (clk), .D (signal_20985), .Q (signal_20986) ) ;
    buf_clk cell_16104 ( .C (clk), .D (signal_20991), .Q (signal_20992) ) ;
    buf_clk cell_16110 ( .C (clk), .D (signal_20997), .Q (signal_20998) ) ;
    buf_clk cell_16116 ( .C (clk), .D (signal_21003), .Q (signal_21004) ) ;
    buf_clk cell_16122 ( .C (clk), .D (signal_21009), .Q (signal_21010) ) ;
    buf_clk cell_16128 ( .C (clk), .D (signal_21015), .Q (signal_21016) ) ;
    buf_clk cell_16134 ( .C (clk), .D (signal_21021), .Q (signal_21022) ) ;
    buf_clk cell_16140 ( .C (clk), .D (signal_21027), .Q (signal_21028) ) ;
    buf_clk cell_16146 ( .C (clk), .D (signal_21033), .Q (signal_21034) ) ;
    buf_clk cell_16152 ( .C (clk), .D (signal_21039), .Q (signal_21040) ) ;
    buf_clk cell_16158 ( .C (clk), .D (signal_21045), .Q (signal_21046) ) ;
    buf_clk cell_16164 ( .C (clk), .D (signal_21051), .Q (signal_21052) ) ;
    buf_clk cell_16170 ( .C (clk), .D (signal_21057), .Q (signal_21058) ) ;
    buf_clk cell_16176 ( .C (clk), .D (signal_21063), .Q (signal_21064) ) ;
    buf_clk cell_16182 ( .C (clk), .D (signal_21069), .Q (signal_21070) ) ;
    buf_clk cell_16188 ( .C (clk), .D (signal_21075), .Q (signal_21076) ) ;
    buf_clk cell_16194 ( .C (clk), .D (signal_21081), .Q (signal_21082) ) ;
    buf_clk cell_16200 ( .C (clk), .D (signal_21087), .Q (signal_21088) ) ;
    buf_clk cell_16206 ( .C (clk), .D (signal_21093), .Q (signal_21094) ) ;
    buf_clk cell_16212 ( .C (clk), .D (signal_21099), .Q (signal_21100) ) ;
    buf_clk cell_16218 ( .C (clk), .D (signal_21105), .Q (signal_21106) ) ;
    buf_clk cell_16224 ( .C (clk), .D (signal_21111), .Q (signal_21112) ) ;
    buf_clk cell_16230 ( .C (clk), .D (signal_21117), .Q (signal_21118) ) ;
    buf_clk cell_16236 ( .C (clk), .D (signal_21123), .Q (signal_21124) ) ;
    buf_clk cell_16242 ( .C (clk), .D (signal_21129), .Q (signal_21130) ) ;
    buf_clk cell_16248 ( .C (clk), .D (signal_21135), .Q (signal_21136) ) ;
    buf_clk cell_16254 ( .C (clk), .D (signal_21141), .Q (signal_21142) ) ;
    buf_clk cell_16260 ( .C (clk), .D (signal_21147), .Q (signal_21148) ) ;
    buf_clk cell_16266 ( .C (clk), .D (signal_21153), .Q (signal_21154) ) ;
    buf_clk cell_16272 ( .C (clk), .D (signal_21159), .Q (signal_21160) ) ;
    buf_clk cell_16278 ( .C (clk), .D (signal_21165), .Q (signal_21166) ) ;
    buf_clk cell_16284 ( .C (clk), .D (signal_21171), .Q (signal_21172) ) ;
    buf_clk cell_16290 ( .C (clk), .D (signal_21177), .Q (signal_21178) ) ;
    buf_clk cell_16296 ( .C (clk), .D (signal_21183), .Q (signal_21184) ) ;
    buf_clk cell_16302 ( .C (clk), .D (signal_21189), .Q (signal_21190) ) ;
    buf_clk cell_16308 ( .C (clk), .D (signal_21195), .Q (signal_21196) ) ;
    buf_clk cell_16314 ( .C (clk), .D (signal_21201), .Q (signal_21202) ) ;
    buf_clk cell_16320 ( .C (clk), .D (signal_21207), .Q (signal_21208) ) ;
    buf_clk cell_16326 ( .C (clk), .D (signal_21213), .Q (signal_21214) ) ;
    buf_clk cell_16332 ( .C (clk), .D (signal_21219), .Q (signal_21220) ) ;
    buf_clk cell_16338 ( .C (clk), .D (signal_21225), .Q (signal_21226) ) ;
    buf_clk cell_16344 ( .C (clk), .D (signal_21231), .Q (signal_21232) ) ;
    buf_clk cell_16350 ( .C (clk), .D (signal_21237), .Q (signal_21238) ) ;
    buf_clk cell_16356 ( .C (clk), .D (signal_21243), .Q (signal_21244) ) ;
    buf_clk cell_16362 ( .C (clk), .D (signal_21249), .Q (signal_21250) ) ;
    buf_clk cell_16368 ( .C (clk), .D (signal_21255), .Q (signal_21256) ) ;
    buf_clk cell_16374 ( .C (clk), .D (signal_21261), .Q (signal_21262) ) ;
    buf_clk cell_16380 ( .C (clk), .D (signal_21267), .Q (signal_21268) ) ;
    buf_clk cell_16386 ( .C (clk), .D (signal_21273), .Q (signal_21274) ) ;
    buf_clk cell_16392 ( .C (clk), .D (signal_21279), .Q (signal_21280) ) ;
    buf_clk cell_16398 ( .C (clk), .D (signal_21285), .Q (signal_21286) ) ;
    buf_clk cell_16404 ( .C (clk), .D (signal_21291), .Q (signal_21292) ) ;
    buf_clk cell_16410 ( .C (clk), .D (signal_21297), .Q (signal_21298) ) ;
    buf_clk cell_16416 ( .C (clk), .D (signal_21303), .Q (signal_21304) ) ;
    buf_clk cell_16422 ( .C (clk), .D (signal_21309), .Q (signal_21310) ) ;
    buf_clk cell_16428 ( .C (clk), .D (signal_21315), .Q (signal_21316) ) ;
    buf_clk cell_16434 ( .C (clk), .D (signal_21321), .Q (signal_21322) ) ;
    buf_clk cell_16440 ( .C (clk), .D (signal_21327), .Q (signal_21328) ) ;
    buf_clk cell_16446 ( .C (clk), .D (signal_21333), .Q (signal_21334) ) ;
    buf_clk cell_16452 ( .C (clk), .D (signal_21339), .Q (signal_21340) ) ;
    buf_clk cell_16458 ( .C (clk), .D (signal_21345), .Q (signal_21346) ) ;
    buf_clk cell_16464 ( .C (clk), .D (signal_21351), .Q (signal_21352) ) ;
    buf_clk cell_16470 ( .C (clk), .D (signal_21357), .Q (signal_21358) ) ;
    buf_clk cell_16476 ( .C (clk), .D (signal_21363), .Q (signal_21364) ) ;
    buf_clk cell_16482 ( .C (clk), .D (signal_21369), .Q (signal_21370) ) ;
    buf_clk cell_16488 ( .C (clk), .D (signal_21375), .Q (signal_21376) ) ;
    buf_clk cell_16494 ( .C (clk), .D (signal_21381), .Q (signal_21382) ) ;
    buf_clk cell_16500 ( .C (clk), .D (signal_21387), .Q (signal_21388) ) ;
    buf_clk cell_16506 ( .C (clk), .D (signal_21393), .Q (signal_21394) ) ;
    buf_clk cell_16512 ( .C (clk), .D (signal_21399), .Q (signal_21400) ) ;
    buf_clk cell_16518 ( .C (clk), .D (signal_21405), .Q (signal_21406) ) ;
    buf_clk cell_16524 ( .C (clk), .D (signal_21411), .Q (signal_21412) ) ;
    buf_clk cell_16530 ( .C (clk), .D (signal_21417), .Q (signal_21418) ) ;
    buf_clk cell_16536 ( .C (clk), .D (signal_21423), .Q (signal_21424) ) ;
    buf_clk cell_16542 ( .C (clk), .D (signal_21429), .Q (signal_21430) ) ;
    buf_clk cell_16548 ( .C (clk), .D (signal_21435), .Q (signal_21436) ) ;
    buf_clk cell_16554 ( .C (clk), .D (signal_21441), .Q (signal_21442) ) ;
    buf_clk cell_16560 ( .C (clk), .D (signal_21447), .Q (signal_21448) ) ;
    buf_clk cell_16566 ( .C (clk), .D (signal_21453), .Q (signal_21454) ) ;
    buf_clk cell_16572 ( .C (clk), .D (signal_21459), .Q (signal_21460) ) ;
    buf_clk cell_16578 ( .C (clk), .D (signal_21465), .Q (signal_21466) ) ;
    buf_clk cell_16584 ( .C (clk), .D (signal_21471), .Q (signal_21472) ) ;
    buf_clk cell_16590 ( .C (clk), .D (signal_21477), .Q (signal_21478) ) ;
    buf_clk cell_16596 ( .C (clk), .D (signal_21483), .Q (signal_21484) ) ;
    buf_clk cell_16602 ( .C (clk), .D (signal_21489), .Q (signal_21490) ) ;
    buf_clk cell_16608 ( .C (clk), .D (signal_21495), .Q (signal_21496) ) ;
    buf_clk cell_16614 ( .C (clk), .D (signal_21501), .Q (signal_21502) ) ;
    buf_clk cell_16620 ( .C (clk), .D (signal_21507), .Q (signal_21508) ) ;
    buf_clk cell_16626 ( .C (clk), .D (signal_21513), .Q (signal_21514) ) ;
    buf_clk cell_16632 ( .C (clk), .D (signal_21519), .Q (signal_21520) ) ;
    buf_clk cell_16638 ( .C (clk), .D (signal_21525), .Q (signal_21526) ) ;
    buf_clk cell_16644 ( .C (clk), .D (signal_21531), .Q (signal_21532) ) ;
    buf_clk cell_16650 ( .C (clk), .D (signal_21537), .Q (signal_21538) ) ;
    buf_clk cell_16656 ( .C (clk), .D (signal_21543), .Q (signal_21544) ) ;
    buf_clk cell_16662 ( .C (clk), .D (signal_21549), .Q (signal_21550) ) ;
    buf_clk cell_16668 ( .C (clk), .D (signal_21555), .Q (signal_21556) ) ;
    buf_clk cell_16674 ( .C (clk), .D (signal_21561), .Q (signal_21562) ) ;
    buf_clk cell_16680 ( .C (clk), .D (signal_21567), .Q (signal_21568) ) ;
    buf_clk cell_16686 ( .C (clk), .D (signal_21573), .Q (signal_21574) ) ;
    buf_clk cell_16692 ( .C (clk), .D (signal_21579), .Q (signal_21580) ) ;
    buf_clk cell_16698 ( .C (clk), .D (signal_21585), .Q (signal_21586) ) ;
    buf_clk cell_16704 ( .C (clk), .D (signal_21591), .Q (signal_21592) ) ;
    buf_clk cell_16710 ( .C (clk), .D (signal_21597), .Q (signal_21598) ) ;
    buf_clk cell_16716 ( .C (clk), .D (signal_21603), .Q (signal_21604) ) ;
    buf_clk cell_16722 ( .C (clk), .D (signal_21609), .Q (signal_21610) ) ;
    buf_clk cell_16728 ( .C (clk), .D (signal_21615), .Q (signal_21616) ) ;
    buf_clk cell_16734 ( .C (clk), .D (signal_21621), .Q (signal_21622) ) ;
    buf_clk cell_16740 ( .C (clk), .D (signal_21627), .Q (signal_21628) ) ;
    buf_clk cell_16746 ( .C (clk), .D (signal_21633), .Q (signal_21634) ) ;
    buf_clk cell_16752 ( .C (clk), .D (signal_21639), .Q (signal_21640) ) ;
    buf_clk cell_16758 ( .C (clk), .D (signal_21645), .Q (signal_21646) ) ;
    buf_clk cell_16764 ( .C (clk), .D (signal_21651), .Q (signal_21652) ) ;
    buf_clk cell_16770 ( .C (clk), .D (signal_21657), .Q (signal_21658) ) ;
    buf_clk cell_16776 ( .C (clk), .D (signal_21663), .Q (signal_21664) ) ;
    buf_clk cell_16782 ( .C (clk), .D (signal_21669), .Q (signal_21670) ) ;
    buf_clk cell_16788 ( .C (clk), .D (signal_21675), .Q (signal_21676) ) ;
    buf_clk cell_16794 ( .C (clk), .D (signal_21681), .Q (signal_21682) ) ;
    buf_clk cell_16800 ( .C (clk), .D (signal_21687), .Q (signal_21688) ) ;
    buf_clk cell_16806 ( .C (clk), .D (signal_21693), .Q (signal_21694) ) ;
    buf_clk cell_16812 ( .C (clk), .D (signal_21699), .Q (signal_21700) ) ;
    buf_clk cell_16818 ( .C (clk), .D (signal_21705), .Q (signal_21706) ) ;
    buf_clk cell_16824 ( .C (clk), .D (signal_21711), .Q (signal_21712) ) ;
    buf_clk cell_16830 ( .C (clk), .D (signal_21717), .Q (signal_21718) ) ;
    buf_clk cell_16836 ( .C (clk), .D (signal_21723), .Q (signal_21724) ) ;
    buf_clk cell_16842 ( .C (clk), .D (signal_21729), .Q (signal_21730) ) ;
    buf_clk cell_16848 ( .C (clk), .D (signal_21735), .Q (signal_21736) ) ;
    buf_clk cell_16854 ( .C (clk), .D (signal_21741), .Q (signal_21742) ) ;
    buf_clk cell_16860 ( .C (clk), .D (signal_21747), .Q (signal_21748) ) ;
    buf_clk cell_16866 ( .C (clk), .D (signal_21753), .Q (signal_21754) ) ;
    buf_clk cell_16872 ( .C (clk), .D (signal_21759), .Q (signal_21760) ) ;
    buf_clk cell_16878 ( .C (clk), .D (signal_21765), .Q (signal_21766) ) ;
    buf_clk cell_16884 ( .C (clk), .D (signal_21771), .Q (signal_21772) ) ;
    buf_clk cell_16890 ( .C (clk), .D (signal_21777), .Q (signal_21778) ) ;
    buf_clk cell_16896 ( .C (clk), .D (signal_21783), .Q (signal_21784) ) ;
    buf_clk cell_16902 ( .C (clk), .D (signal_21789), .Q (signal_21790) ) ;
    buf_clk cell_16908 ( .C (clk), .D (signal_21795), .Q (signal_21796) ) ;
    buf_clk cell_16914 ( .C (clk), .D (signal_21801), .Q (signal_21802) ) ;
    buf_clk cell_16920 ( .C (clk), .D (signal_21807), .Q (signal_21808) ) ;
    buf_clk cell_16926 ( .C (clk), .D (signal_21813), .Q (signal_21814) ) ;
    buf_clk cell_16932 ( .C (clk), .D (signal_21819), .Q (signal_21820) ) ;
    buf_clk cell_16938 ( .C (clk), .D (signal_21825), .Q (signal_21826) ) ;
    buf_clk cell_16944 ( .C (clk), .D (signal_21831), .Q (signal_21832) ) ;
    buf_clk cell_16950 ( .C (clk), .D (signal_21837), .Q (signal_21838) ) ;
    buf_clk cell_16956 ( .C (clk), .D (signal_21843), .Q (signal_21844) ) ;
    buf_clk cell_16962 ( .C (clk), .D (signal_21849), .Q (signal_21850) ) ;
    buf_clk cell_16968 ( .C (clk), .D (signal_21855), .Q (signal_21856) ) ;
    buf_clk cell_16974 ( .C (clk), .D (signal_21861), .Q (signal_21862) ) ;
    buf_clk cell_16980 ( .C (clk), .D (signal_21867), .Q (signal_21868) ) ;
    buf_clk cell_16986 ( .C (clk), .D (signal_21873), .Q (signal_21874) ) ;
    buf_clk cell_16992 ( .C (clk), .D (signal_21879), .Q (signal_21880) ) ;
    buf_clk cell_16998 ( .C (clk), .D (signal_21885), .Q (signal_21886) ) ;
    buf_clk cell_17004 ( .C (clk), .D (signal_21891), .Q (signal_21892) ) ;
    buf_clk cell_17010 ( .C (clk), .D (signal_21897), .Q (signal_21898) ) ;
    buf_clk cell_17016 ( .C (clk), .D (signal_21903), .Q (signal_21904) ) ;
    buf_clk cell_17022 ( .C (clk), .D (signal_21909), .Q (signal_21910) ) ;
    buf_clk cell_17028 ( .C (clk), .D (signal_21915), .Q (signal_21916) ) ;
    buf_clk cell_17034 ( .C (clk), .D (signal_21921), .Q (signal_21922) ) ;
    buf_clk cell_17040 ( .C (clk), .D (signal_21927), .Q (signal_21928) ) ;
    buf_clk cell_17046 ( .C (clk), .D (signal_21933), .Q (signal_21934) ) ;
    buf_clk cell_17052 ( .C (clk), .D (signal_21939), .Q (signal_21940) ) ;
    buf_clk cell_17058 ( .C (clk), .D (signal_21945), .Q (signal_21946) ) ;
    buf_clk cell_17064 ( .C (clk), .D (signal_21951), .Q (signal_21952) ) ;
    buf_clk cell_17070 ( .C (clk), .D (signal_21957), .Q (signal_21958) ) ;
    buf_clk cell_17076 ( .C (clk), .D (signal_21963), .Q (signal_21964) ) ;
    buf_clk cell_17082 ( .C (clk), .D (signal_21969), .Q (signal_21970) ) ;
    buf_clk cell_17088 ( .C (clk), .D (signal_21975), .Q (signal_21976) ) ;
    buf_clk cell_17094 ( .C (clk), .D (signal_21981), .Q (signal_21982) ) ;
    buf_clk cell_17100 ( .C (clk), .D (signal_21987), .Q (signal_21988) ) ;
    buf_clk cell_17106 ( .C (clk), .D (signal_21993), .Q (signal_21994) ) ;
    buf_clk cell_17112 ( .C (clk), .D (signal_21999), .Q (signal_22000) ) ;
    buf_clk cell_17118 ( .C (clk), .D (signal_22005), .Q (signal_22006) ) ;
    buf_clk cell_17124 ( .C (clk), .D (signal_22011), .Q (signal_22012) ) ;
    buf_clk cell_17130 ( .C (clk), .D (signal_22017), .Q (signal_22018) ) ;
    buf_clk cell_17136 ( .C (clk), .D (signal_22023), .Q (signal_22024) ) ;
    buf_clk cell_17142 ( .C (clk), .D (signal_22029), .Q (signal_22030) ) ;
    buf_clk cell_17148 ( .C (clk), .D (signal_22035), .Q (signal_22036) ) ;
    buf_clk cell_17154 ( .C (clk), .D (signal_22041), .Q (signal_22042) ) ;
    buf_clk cell_17160 ( .C (clk), .D (signal_22047), .Q (signal_22048) ) ;
    buf_clk cell_17166 ( .C (clk), .D (signal_22053), .Q (signal_22054) ) ;
    buf_clk cell_17172 ( .C (clk), .D (signal_22059), .Q (signal_22060) ) ;
    buf_clk cell_17178 ( .C (clk), .D (signal_22065), .Q (signal_22066) ) ;
    buf_clk cell_17184 ( .C (clk), .D (signal_22071), .Q (signal_22072) ) ;
    buf_clk cell_17190 ( .C (clk), .D (signal_22077), .Q (signal_22078) ) ;
    buf_clk cell_17196 ( .C (clk), .D (signal_22083), .Q (signal_22084) ) ;
    buf_clk cell_17202 ( .C (clk), .D (signal_22089), .Q (signal_22090) ) ;
    buf_clk cell_17208 ( .C (clk), .D (signal_22095), .Q (signal_22096) ) ;
    buf_clk cell_17214 ( .C (clk), .D (signal_22101), .Q (signal_22102) ) ;
    buf_clk cell_17220 ( .C (clk), .D (signal_22107), .Q (signal_22108) ) ;
    buf_clk cell_17226 ( .C (clk), .D (signal_22113), .Q (signal_22114) ) ;
    buf_clk cell_17232 ( .C (clk), .D (signal_22119), .Q (signal_22120) ) ;
    buf_clk cell_17238 ( .C (clk), .D (signal_22125), .Q (signal_22126) ) ;
    buf_clk cell_17244 ( .C (clk), .D (signal_22131), .Q (signal_22132) ) ;
    buf_clk cell_17250 ( .C (clk), .D (signal_22137), .Q (signal_22138) ) ;
    buf_clk cell_17256 ( .C (clk), .D (signal_22143), .Q (signal_22144) ) ;
    buf_clk cell_17262 ( .C (clk), .D (signal_22149), .Q (signal_22150) ) ;
    buf_clk cell_17268 ( .C (clk), .D (signal_22155), .Q (signal_22156) ) ;
    buf_clk cell_17274 ( .C (clk), .D (signal_22161), .Q (signal_22162) ) ;
    buf_clk cell_17280 ( .C (clk), .D (signal_22167), .Q (signal_22168) ) ;
    buf_clk cell_17286 ( .C (clk), .D (signal_22173), .Q (signal_22174) ) ;
    buf_clk cell_17292 ( .C (clk), .D (signal_22179), .Q (signal_22180) ) ;
    buf_clk cell_17298 ( .C (clk), .D (signal_22185), .Q (signal_22186) ) ;
    buf_clk cell_17304 ( .C (clk), .D (signal_22191), .Q (signal_22192) ) ;
    buf_clk cell_17310 ( .C (clk), .D (signal_22197), .Q (signal_22198) ) ;
    buf_clk cell_17316 ( .C (clk), .D (signal_22203), .Q (signal_22204) ) ;
    buf_clk cell_17322 ( .C (clk), .D (signal_22209), .Q (signal_22210) ) ;
    buf_clk cell_17328 ( .C (clk), .D (signal_22215), .Q (signal_22216) ) ;
    buf_clk cell_17334 ( .C (clk), .D (signal_22221), .Q (signal_22222) ) ;
    buf_clk cell_17340 ( .C (clk), .D (signal_22227), .Q (signal_22228) ) ;
    buf_clk cell_17346 ( .C (clk), .D (signal_22233), .Q (signal_22234) ) ;
    buf_clk cell_17352 ( .C (clk), .D (signal_22239), .Q (signal_22240) ) ;
    buf_clk cell_17358 ( .C (clk), .D (signal_22245), .Q (signal_22246) ) ;
    buf_clk cell_17364 ( .C (clk), .D (signal_22251), .Q (signal_22252) ) ;
    buf_clk cell_17370 ( .C (clk), .D (signal_22257), .Q (signal_22258) ) ;
    buf_clk cell_17376 ( .C (clk), .D (signal_22263), .Q (signal_22264) ) ;
    buf_clk cell_17382 ( .C (clk), .D (signal_22269), .Q (signal_22270) ) ;
    buf_clk cell_17388 ( .C (clk), .D (signal_22275), .Q (signal_22276) ) ;
    buf_clk cell_17394 ( .C (clk), .D (signal_22281), .Q (signal_22282) ) ;
    buf_clk cell_17400 ( .C (clk), .D (signal_22287), .Q (signal_22288) ) ;
    buf_clk cell_17406 ( .C (clk), .D (signal_22293), .Q (signal_22294) ) ;
    buf_clk cell_17412 ( .C (clk), .D (signal_22299), .Q (signal_22300) ) ;
    buf_clk cell_17418 ( .C (clk), .D (signal_22305), .Q (signal_22306) ) ;
    buf_clk cell_17424 ( .C (clk), .D (signal_22311), .Q (signal_22312) ) ;
    buf_clk cell_17430 ( .C (clk), .D (signal_22317), .Q (signal_22318) ) ;
    buf_clk cell_17436 ( .C (clk), .D (signal_22323), .Q (signal_22324) ) ;
    buf_clk cell_17442 ( .C (clk), .D (signal_22329), .Q (signal_22330) ) ;
    buf_clk cell_17448 ( .C (clk), .D (signal_22335), .Q (signal_22336) ) ;
    buf_clk cell_17454 ( .C (clk), .D (signal_22341), .Q (signal_22342) ) ;
    buf_clk cell_17460 ( .C (clk), .D (signal_22347), .Q (signal_22348) ) ;
    buf_clk cell_17466 ( .C (clk), .D (signal_22353), .Q (signal_22354) ) ;
    buf_clk cell_17472 ( .C (clk), .D (signal_22359), .Q (signal_22360) ) ;
    buf_clk cell_17478 ( .C (clk), .D (signal_22365), .Q (signal_22366) ) ;
    buf_clk cell_17484 ( .C (clk), .D (signal_22371), .Q (signal_22372) ) ;
    buf_clk cell_17490 ( .C (clk), .D (signal_22377), .Q (signal_22378) ) ;
    buf_clk cell_17496 ( .C (clk), .D (signal_22383), .Q (signal_22384) ) ;
    buf_clk cell_17502 ( .C (clk), .D (signal_22389), .Q (signal_22390) ) ;
    buf_clk cell_17508 ( .C (clk), .D (signal_22395), .Q (signal_22396) ) ;
    buf_clk cell_17514 ( .C (clk), .D (signal_22401), .Q (signal_22402) ) ;
    buf_clk cell_17520 ( .C (clk), .D (signal_22407), .Q (signal_22408) ) ;
    buf_clk cell_17526 ( .C (clk), .D (signal_22413), .Q (signal_22414) ) ;
    buf_clk cell_17532 ( .C (clk), .D (signal_22419), .Q (signal_22420) ) ;
    buf_clk cell_17538 ( .C (clk), .D (signal_22425), .Q (signal_22426) ) ;
    buf_clk cell_17544 ( .C (clk), .D (signal_22431), .Q (signal_22432) ) ;
    buf_clk cell_17550 ( .C (clk), .D (signal_22437), .Q (signal_22438) ) ;
    buf_clk cell_17556 ( .C (clk), .D (signal_22443), .Q (signal_22444) ) ;
    buf_clk cell_17562 ( .C (clk), .D (signal_22449), .Q (signal_22450) ) ;
    buf_clk cell_17568 ( .C (clk), .D (signal_22455), .Q (signal_22456) ) ;
    buf_clk cell_17574 ( .C (clk), .D (signal_22461), .Q (signal_22462) ) ;
    buf_clk cell_17580 ( .C (clk), .D (signal_22467), .Q (signal_22468) ) ;
    buf_clk cell_17586 ( .C (clk), .D (signal_22473), .Q (signal_22474) ) ;
    buf_clk cell_17594 ( .C (clk), .D (signal_22481), .Q (signal_22482) ) ;
    buf_clk cell_17602 ( .C (clk), .D (signal_22489), .Q (signal_22490) ) ;
    buf_clk cell_17610 ( .C (clk), .D (signal_22497), .Q (signal_22498) ) ;
    buf_clk cell_17618 ( .C (clk), .D (signal_22505), .Q (signal_22506) ) ;
    buf_clk cell_17626 ( .C (clk), .D (signal_22513), .Q (signal_22514) ) ;
    buf_clk cell_17634 ( .C (clk), .D (signal_22521), .Q (signal_22522) ) ;
    buf_clk cell_17642 ( .C (clk), .D (signal_22529), .Q (signal_22530) ) ;
    buf_clk cell_17650 ( .C (clk), .D (signal_22537), .Q (signal_22538) ) ;
    buf_clk cell_17658 ( .C (clk), .D (signal_22545), .Q (signal_22546) ) ;
    buf_clk cell_17666 ( .C (clk), .D (signal_22553), .Q (signal_22554) ) ;
    buf_clk cell_17674 ( .C (clk), .D (signal_22561), .Q (signal_22562) ) ;
    buf_clk cell_17682 ( .C (clk), .D (signal_22569), .Q (signal_22570) ) ;
    buf_clk cell_17690 ( .C (clk), .D (signal_22577), .Q (signal_22578) ) ;
    buf_clk cell_17698 ( .C (clk), .D (signal_22585), .Q (signal_22586) ) ;
    buf_clk cell_17706 ( .C (clk), .D (signal_22593), .Q (signal_22594) ) ;
    buf_clk cell_17714 ( .C (clk), .D (signal_22601), .Q (signal_22602) ) ;
    buf_clk cell_17722 ( .C (clk), .D (signal_22609), .Q (signal_22610) ) ;
    buf_clk cell_17730 ( .C (clk), .D (signal_22617), .Q (signal_22618) ) ;
    buf_clk cell_17738 ( .C (clk), .D (signal_22625), .Q (signal_22626) ) ;
    buf_clk cell_17746 ( .C (clk), .D (signal_22633), .Q (signal_22634) ) ;
    buf_clk cell_17754 ( .C (clk), .D (signal_22641), .Q (signal_22642) ) ;
    buf_clk cell_17762 ( .C (clk), .D (signal_22649), .Q (signal_22650) ) ;
    buf_clk cell_17770 ( .C (clk), .D (signal_22657), .Q (signal_22658) ) ;
    buf_clk cell_17778 ( .C (clk), .D (signal_22665), .Q (signal_22666) ) ;
    buf_clk cell_17786 ( .C (clk), .D (signal_22673), .Q (signal_22674) ) ;
    buf_clk cell_17794 ( .C (clk), .D (signal_22681), .Q (signal_22682) ) ;
    buf_clk cell_17802 ( .C (clk), .D (signal_22689), .Q (signal_22690) ) ;
    buf_clk cell_17810 ( .C (clk), .D (signal_22697), .Q (signal_22698) ) ;
    buf_clk cell_17818 ( .C (clk), .D (signal_22705), .Q (signal_22706) ) ;
    buf_clk cell_17826 ( .C (clk), .D (signal_22713), .Q (signal_22714) ) ;
    buf_clk cell_17834 ( .C (clk), .D (signal_22721), .Q (signal_22722) ) ;
    buf_clk cell_17842 ( .C (clk), .D (signal_22729), .Q (signal_22730) ) ;
    buf_clk cell_17850 ( .C (clk), .D (signal_22737), .Q (signal_22738) ) ;
    buf_clk cell_17858 ( .C (clk), .D (signal_22745), .Q (signal_22746) ) ;
    buf_clk cell_17866 ( .C (clk), .D (signal_22753), .Q (signal_22754) ) ;
    buf_clk cell_17874 ( .C (clk), .D (signal_22761), .Q (signal_22762) ) ;
    buf_clk cell_17882 ( .C (clk), .D (signal_22769), .Q (signal_22770) ) ;
    buf_clk cell_17890 ( .C (clk), .D (signal_22777), .Q (signal_22778) ) ;
    buf_clk cell_17898 ( .C (clk), .D (signal_22785), .Q (signal_22786) ) ;
    buf_clk cell_17906 ( .C (clk), .D (signal_22793), .Q (signal_22794) ) ;
    buf_clk cell_17914 ( .C (clk), .D (signal_22801), .Q (signal_22802) ) ;
    buf_clk cell_17922 ( .C (clk), .D (signal_22809), .Q (signal_22810) ) ;
    buf_clk cell_17930 ( .C (clk), .D (signal_22817), .Q (signal_22818) ) ;
    buf_clk cell_17938 ( .C (clk), .D (signal_22825), .Q (signal_22826) ) ;
    buf_clk cell_17946 ( .C (clk), .D (signal_22833), .Q (signal_22834) ) ;
    buf_clk cell_17954 ( .C (clk), .D (signal_22841), .Q (signal_22842) ) ;
    buf_clk cell_17962 ( .C (clk), .D (signal_22849), .Q (signal_22850) ) ;
    buf_clk cell_17970 ( .C (clk), .D (signal_22857), .Q (signal_22858) ) ;
    buf_clk cell_17978 ( .C (clk), .D (signal_22865), .Q (signal_22866) ) ;
    buf_clk cell_17986 ( .C (clk), .D (signal_22873), .Q (signal_22874) ) ;
    buf_clk cell_17994 ( .C (clk), .D (signal_22881), .Q (signal_22882) ) ;
    buf_clk cell_18002 ( .C (clk), .D (signal_22889), .Q (signal_22890) ) ;
    buf_clk cell_18010 ( .C (clk), .D (signal_22897), .Q (signal_22898) ) ;
    buf_clk cell_18018 ( .C (clk), .D (signal_22905), .Q (signal_22906) ) ;
    buf_clk cell_18026 ( .C (clk), .D (signal_22913), .Q (signal_22914) ) ;
    buf_clk cell_18034 ( .C (clk), .D (signal_22921), .Q (signal_22922) ) ;
    buf_clk cell_18042 ( .C (clk), .D (signal_22929), .Q (signal_22930) ) ;
    buf_clk cell_18050 ( .C (clk), .D (signal_22937), .Q (signal_22938) ) ;
    buf_clk cell_18058 ( .C (clk), .D (signal_22945), .Q (signal_22946) ) ;
    buf_clk cell_18066 ( .C (clk), .D (signal_22953), .Q (signal_22954) ) ;
    buf_clk cell_18074 ( .C (clk), .D (signal_22961), .Q (signal_22962) ) ;
    buf_clk cell_18082 ( .C (clk), .D (signal_22969), .Q (signal_22970) ) ;
    buf_clk cell_18090 ( .C (clk), .D (signal_22977), .Q (signal_22978) ) ;
    buf_clk cell_18098 ( .C (clk), .D (signal_22985), .Q (signal_22986) ) ;
    buf_clk cell_18106 ( .C (clk), .D (signal_22993), .Q (signal_22994) ) ;
    buf_clk cell_18114 ( .C (clk), .D (signal_23001), .Q (signal_23002) ) ;
    buf_clk cell_18122 ( .C (clk), .D (signal_23009), .Q (signal_23010) ) ;
    buf_clk cell_18130 ( .C (clk), .D (signal_23017), .Q (signal_23018) ) ;
    buf_clk cell_18138 ( .C (clk), .D (signal_23025), .Q (signal_23026) ) ;
    buf_clk cell_18146 ( .C (clk), .D (signal_23033), .Q (signal_23034) ) ;
    buf_clk cell_18154 ( .C (clk), .D (signal_23041), .Q (signal_23042) ) ;
    buf_clk cell_18162 ( .C (clk), .D (signal_23049), .Q (signal_23050) ) ;
    buf_clk cell_18170 ( .C (clk), .D (signal_23057), .Q (signal_23058) ) ;
    buf_clk cell_18178 ( .C (clk), .D (signal_23065), .Q (signal_23066) ) ;
    buf_clk cell_18186 ( .C (clk), .D (signal_23073), .Q (signal_23074) ) ;
    buf_clk cell_18194 ( .C (clk), .D (signal_23081), .Q (signal_23082) ) ;
    buf_clk cell_18202 ( .C (clk), .D (signal_23089), .Q (signal_23090) ) ;
    buf_clk cell_18210 ( .C (clk), .D (signal_23097), .Q (signal_23098) ) ;
    buf_clk cell_18218 ( .C (clk), .D (signal_23105), .Q (signal_23106) ) ;
    buf_clk cell_18226 ( .C (clk), .D (signal_23113), .Q (signal_23114) ) ;
    buf_clk cell_18234 ( .C (clk), .D (signal_23121), .Q (signal_23122) ) ;
    buf_clk cell_18242 ( .C (clk), .D (signal_23129), .Q (signal_23130) ) ;
    buf_clk cell_18250 ( .C (clk), .D (signal_23137), .Q (signal_23138) ) ;
    buf_clk cell_18258 ( .C (clk), .D (signal_23145), .Q (signal_23146) ) ;
    buf_clk cell_18266 ( .C (clk), .D (signal_23153), .Q (signal_23154) ) ;
    buf_clk cell_18274 ( .C (clk), .D (signal_23161), .Q (signal_23162) ) ;
    buf_clk cell_18282 ( .C (clk), .D (signal_23169), .Q (signal_23170) ) ;
    buf_clk cell_18290 ( .C (clk), .D (signal_23177), .Q (signal_23178) ) ;
    buf_clk cell_18298 ( .C (clk), .D (signal_23185), .Q (signal_23186) ) ;
    buf_clk cell_18306 ( .C (clk), .D (signal_23193), .Q (signal_23194) ) ;
    buf_clk cell_18314 ( .C (clk), .D (signal_23201), .Q (signal_23202) ) ;
    buf_clk cell_18322 ( .C (clk), .D (signal_23209), .Q (signal_23210) ) ;
    buf_clk cell_18330 ( .C (clk), .D (signal_23217), .Q (signal_23218) ) ;
    buf_clk cell_18338 ( .C (clk), .D (signal_23225), .Q (signal_23226) ) ;
    buf_clk cell_18346 ( .C (clk), .D (signal_23233), .Q (signal_23234) ) ;
    buf_clk cell_18354 ( .C (clk), .D (signal_23241), .Q (signal_23242) ) ;
    buf_clk cell_18362 ( .C (clk), .D (signal_23249), .Q (signal_23250) ) ;
    buf_clk cell_18370 ( .C (clk), .D (signal_23257), .Q (signal_23258) ) ;
    buf_clk cell_18378 ( .C (clk), .D (signal_23265), .Q (signal_23266) ) ;
    buf_clk cell_18386 ( .C (clk), .D (signal_23273), .Q (signal_23274) ) ;
    buf_clk cell_18394 ( .C (clk), .D (signal_23281), .Q (signal_23282) ) ;
    buf_clk cell_18406 ( .C (clk), .D (signal_23293), .Q (signal_23294) ) ;
    buf_clk cell_18414 ( .C (clk), .D (signal_23301), .Q (signal_23302) ) ;
    buf_clk cell_18422 ( .C (clk), .D (signal_23309), .Q (signal_23310) ) ;
    buf_clk cell_18430 ( .C (clk), .D (signal_23317), .Q (signal_23318) ) ;
    buf_clk cell_18438 ( .C (clk), .D (signal_23325), .Q (signal_23326) ) ;
    buf_clk cell_18446 ( .C (clk), .D (signal_23333), .Q (signal_23334) ) ;
    buf_clk cell_18454 ( .C (clk), .D (signal_23341), .Q (signal_23342) ) ;
    buf_clk cell_18462 ( .C (clk), .D (signal_23349), .Q (signal_23350) ) ;
    buf_clk cell_18470 ( .C (clk), .D (signal_23357), .Q (signal_23358) ) ;
    buf_clk cell_18478 ( .C (clk), .D (signal_23365), .Q (signal_23366) ) ;
    buf_clk cell_18486 ( .C (clk), .D (signal_23373), .Q (signal_23374) ) ;
    buf_clk cell_18494 ( .C (clk), .D (signal_23381), .Q (signal_23382) ) ;
    buf_clk cell_18502 ( .C (clk), .D (signal_23389), .Q (signal_23390) ) ;
    buf_clk cell_18510 ( .C (clk), .D (signal_23397), .Q (signal_23398) ) ;
    buf_clk cell_18518 ( .C (clk), .D (signal_23405), .Q (signal_23406) ) ;
    buf_clk cell_18526 ( .C (clk), .D (signal_23413), .Q (signal_23414) ) ;
    buf_clk cell_18534 ( .C (clk), .D (signal_23421), .Q (signal_23422) ) ;
    buf_clk cell_18542 ( .C (clk), .D (signal_23429), .Q (signal_23430) ) ;
    buf_clk cell_18550 ( .C (clk), .D (signal_23437), .Q (signal_23438) ) ;
    buf_clk cell_18558 ( .C (clk), .D (signal_23445), .Q (signal_23446) ) ;
    buf_clk cell_18566 ( .C (clk), .D (signal_23453), .Q (signal_23454) ) ;
    buf_clk cell_18574 ( .C (clk), .D (signal_23461), .Q (signal_23462) ) ;
    buf_clk cell_18582 ( .C (clk), .D (signal_23469), .Q (signal_23470) ) ;
    buf_clk cell_18590 ( .C (clk), .D (signal_23477), .Q (signal_23478) ) ;
    buf_clk cell_18598 ( .C (clk), .D (signal_23485), .Q (signal_23486) ) ;
    buf_clk cell_18606 ( .C (clk), .D (signal_23493), .Q (signal_23494) ) ;
    buf_clk cell_18614 ( .C (clk), .D (signal_23501), .Q (signal_23502) ) ;
    buf_clk cell_18622 ( .C (clk), .D (signal_23509), .Q (signal_23510) ) ;
    buf_clk cell_18630 ( .C (clk), .D (signal_23517), .Q (signal_23518) ) ;
    buf_clk cell_18638 ( .C (clk), .D (signal_23525), .Q (signal_23526) ) ;
    buf_clk cell_18650 ( .C (clk), .D (signal_23537), .Q (signal_23538) ) ;
    buf_clk cell_18658 ( .C (clk), .D (signal_23545), .Q (signal_23546) ) ;
    buf_clk cell_18666 ( .C (clk), .D (signal_23553), .Q (signal_23554) ) ;
    buf_clk cell_18674 ( .C (clk), .D (signal_23561), .Q (signal_23562) ) ;
    buf_clk cell_18682 ( .C (clk), .D (signal_23569), .Q (signal_23570) ) ;
    buf_clk cell_18690 ( .C (clk), .D (signal_23577), .Q (signal_23578) ) ;
    buf_clk cell_18698 ( .C (clk), .D (signal_23585), .Q (signal_23586) ) ;
    buf_clk cell_18706 ( .C (clk), .D (signal_23593), .Q (signal_23594) ) ;
    buf_clk cell_18714 ( .C (clk), .D (signal_23601), .Q (signal_23602) ) ;
    buf_clk cell_18722 ( .C (clk), .D (signal_23609), .Q (signal_23610) ) ;
    buf_clk cell_18730 ( .C (clk), .D (signal_23617), .Q (signal_23618) ) ;
    buf_clk cell_18738 ( .C (clk), .D (signal_23625), .Q (signal_23626) ) ;
    buf_clk cell_18750 ( .C (clk), .D (signal_23637), .Q (signal_23638) ) ;
    buf_clk cell_18758 ( .C (clk), .D (signal_23645), .Q (signal_23646) ) ;
    buf_clk cell_18766 ( .C (clk), .D (signal_23653), .Q (signal_23654) ) ;
    buf_clk cell_18774 ( .C (clk), .D (signal_23661), .Q (signal_23662) ) ;
    buf_clk cell_18782 ( .C (clk), .D (signal_23669), .Q (signal_23670) ) ;
    buf_clk cell_18790 ( .C (clk), .D (signal_23677), .Q (signal_23678) ) ;
    buf_clk cell_18798 ( .C (clk), .D (signal_23685), .Q (signal_23686) ) ;
    buf_clk cell_18806 ( .C (clk), .D (signal_23693), .Q (signal_23694) ) ;
    buf_clk cell_18814 ( .C (clk), .D (signal_23701), .Q (signal_23702) ) ;
    buf_clk cell_18822 ( .C (clk), .D (signal_23709), .Q (signal_23710) ) ;
    buf_clk cell_18830 ( .C (clk), .D (signal_23717), .Q (signal_23718) ) ;
    buf_clk cell_18838 ( .C (clk), .D (signal_23725), .Q (signal_23726) ) ;
    buf_clk cell_18846 ( .C (clk), .D (signal_23733), .Q (signal_23734) ) ;
    buf_clk cell_18854 ( .C (clk), .D (signal_23741), .Q (signal_23742) ) ;
    buf_clk cell_18862 ( .C (clk), .D (signal_23749), .Q (signal_23750) ) ;
    buf_clk cell_18870 ( .C (clk), .D (signal_23757), .Q (signal_23758) ) ;
    buf_clk cell_18878 ( .C (clk), .D (signal_23765), .Q (signal_23766) ) ;
    buf_clk cell_18886 ( .C (clk), .D (signal_23773), .Q (signal_23774) ) ;
    buf_clk cell_18894 ( .C (clk), .D (signal_23781), .Q (signal_23782) ) ;
    buf_clk cell_18902 ( .C (clk), .D (signal_23789), .Q (signal_23790) ) ;
    buf_clk cell_18910 ( .C (clk), .D (signal_23797), .Q (signal_23798) ) ;
    buf_clk cell_18918 ( .C (clk), .D (signal_23805), .Q (signal_23806) ) ;
    buf_clk cell_18926 ( .C (clk), .D (signal_23813), .Q (signal_23814) ) ;
    buf_clk cell_18934 ( .C (clk), .D (signal_23821), .Q (signal_23822) ) ;
    buf_clk cell_18942 ( .C (clk), .D (signal_23829), .Q (signal_23830) ) ;
    buf_clk cell_18950 ( .C (clk), .D (signal_23837), .Q (signal_23838) ) ;
    buf_clk cell_18958 ( .C (clk), .D (signal_23845), .Q (signal_23846) ) ;
    buf_clk cell_18966 ( .C (clk), .D (signal_23853), .Q (signal_23854) ) ;
    buf_clk cell_18974 ( .C (clk), .D (signal_23861), .Q (signal_23862) ) ;
    buf_clk cell_18982 ( .C (clk), .D (signal_23869), .Q (signal_23870) ) ;
    buf_clk cell_18990 ( .C (clk), .D (signal_23877), .Q (signal_23878) ) ;
    buf_clk cell_18998 ( .C (clk), .D (signal_23885), .Q (signal_23886) ) ;
    buf_clk cell_19006 ( .C (clk), .D (signal_23893), .Q (signal_23894) ) ;
    buf_clk cell_19014 ( .C (clk), .D (signal_23901), .Q (signal_23902) ) ;
    buf_clk cell_19022 ( .C (clk), .D (signal_23909), .Q (signal_23910) ) ;
    buf_clk cell_19030 ( .C (clk), .D (signal_23917), .Q (signal_23918) ) ;
    buf_clk cell_19038 ( .C (clk), .D (signal_23925), .Q (signal_23926) ) ;
    buf_clk cell_19046 ( .C (clk), .D (signal_23933), .Q (signal_23934) ) ;
    buf_clk cell_19054 ( .C (clk), .D (signal_23941), .Q (signal_23942) ) ;
    buf_clk cell_19062 ( .C (clk), .D (signal_23949), .Q (signal_23950) ) ;
    buf_clk cell_19070 ( .C (clk), .D (signal_23957), .Q (signal_23958) ) ;
    buf_clk cell_19078 ( .C (clk), .D (signal_23965), .Q (signal_23966) ) ;
    buf_clk cell_19086 ( .C (clk), .D (signal_23973), .Q (signal_23974) ) ;
    buf_clk cell_19094 ( .C (clk), .D (signal_23981), .Q (signal_23982) ) ;
    buf_clk cell_19102 ( .C (clk), .D (signal_23989), .Q (signal_23990) ) ;
    buf_clk cell_19110 ( .C (clk), .D (signal_23997), .Q (signal_23998) ) ;

    /* cells in depth 3 */
    buf_clk cell_7901 ( .C (clk), .D (signal_5421), .Q (signal_12789) ) ;
    buf_clk cell_7903 ( .C (clk), .D (signal_8759), .Q (signal_12791) ) ;
    buf_clk cell_7905 ( .C (clk), .D (signal_5519), .Q (signal_12793) ) ;
    buf_clk cell_7907 ( .C (clk), .D (signal_8843), .Q (signal_12795) ) ;
    buf_clk cell_7909 ( .C (clk), .D (signal_5520), .Q (signal_12797) ) ;
    buf_clk cell_7911 ( .C (clk), .D (signal_8844), .Q (signal_12799) ) ;
    buf_clk cell_7913 ( .C (clk), .D (signal_5440), .Q (signal_12801) ) ;
    buf_clk cell_7915 ( .C (clk), .D (signal_8763), .Q (signal_12803) ) ;
    buf_clk cell_7917 ( .C (clk), .D (signal_5533), .Q (signal_12805) ) ;
    buf_clk cell_7919 ( .C (clk), .D (signal_8845), .Q (signal_12807) ) ;
    buf_clk cell_7921 ( .C (clk), .D (signal_5534), .Q (signal_12809) ) ;
    buf_clk cell_7923 ( .C (clk), .D (signal_8846), .Q (signal_12811) ) ;
    buf_clk cell_7925 ( .C (clk), .D (signal_5459), .Q (signal_12813) ) ;
    buf_clk cell_7927 ( .C (clk), .D (signal_8767), .Q (signal_12815) ) ;
    buf_clk cell_7929 ( .C (clk), .D (signal_5547), .Q (signal_12817) ) ;
    buf_clk cell_7931 ( .C (clk), .D (signal_8847), .Q (signal_12819) ) ;
    buf_clk cell_7933 ( .C (clk), .D (signal_5548), .Q (signal_12821) ) ;
    buf_clk cell_7935 ( .C (clk), .D (signal_8848), .Q (signal_12823) ) ;
    buf_clk cell_7937 ( .C (clk), .D (signal_5463), .Q (signal_12825) ) ;
    buf_clk cell_7939 ( .C (clk), .D (signal_8743), .Q (signal_12827) ) ;
    buf_clk cell_7941 ( .C (clk), .D (signal_5549), .Q (signal_12829) ) ;
    buf_clk cell_7943 ( .C (clk), .D (signal_8829), .Q (signal_12831) ) ;
    buf_clk cell_7945 ( .C (clk), .D (signal_5550), .Q (signal_12833) ) ;
    buf_clk cell_7947 ( .C (clk), .D (signal_8830), .Q (signal_12835) ) ;
    buf_clk cell_7949 ( .C (clk), .D (signal_5467), .Q (signal_12837) ) ;
    buf_clk cell_7951 ( .C (clk), .D (signal_8747), .Q (signal_12839) ) ;
    buf_clk cell_7953 ( .C (clk), .D (signal_5551), .Q (signal_12841) ) ;
    buf_clk cell_7955 ( .C (clk), .D (signal_8831), .Q (signal_12843) ) ;
    buf_clk cell_7957 ( .C (clk), .D (signal_5552), .Q (signal_12845) ) ;
    buf_clk cell_7959 ( .C (clk), .D (signal_8832), .Q (signal_12847) ) ;
    buf_clk cell_7961 ( .C (clk), .D (signal_5471), .Q (signal_12849) ) ;
    buf_clk cell_7963 ( .C (clk), .D (signal_8751), .Q (signal_12851) ) ;
    buf_clk cell_7965 ( .C (clk), .D (signal_5553), .Q (signal_12853) ) ;
    buf_clk cell_7967 ( .C (clk), .D (signal_8833), .Q (signal_12855) ) ;
    buf_clk cell_7969 ( .C (clk), .D (signal_5554), .Q (signal_12857) ) ;
    buf_clk cell_7971 ( .C (clk), .D (signal_8834), .Q (signal_12859) ) ;
    buf_clk cell_7973 ( .C (clk), .D (signal_5475), .Q (signal_12861) ) ;
    buf_clk cell_7975 ( .C (clk), .D (signal_8755), .Q (signal_12863) ) ;
    buf_clk cell_7977 ( .C (clk), .D (signal_5555), .Q (signal_12865) ) ;
    buf_clk cell_7979 ( .C (clk), .D (signal_8835), .Q (signal_12867) ) ;
    buf_clk cell_7981 ( .C (clk), .D (signal_5556), .Q (signal_12869) ) ;
    buf_clk cell_7983 ( .C (clk), .D (signal_8836), .Q (signal_12871) ) ;
    buf_clk cell_7985 ( .C (clk), .D (signal_5493), .Q (signal_12873) ) ;
    buf_clk cell_7987 ( .C (clk), .D (signal_8779), .Q (signal_12875) ) ;
    buf_clk cell_7989 ( .C (clk), .D (signal_5590), .Q (signal_12877) ) ;
    buf_clk cell_7991 ( .C (clk), .D (signal_8879), .Q (signal_12879) ) ;
    buf_clk cell_7993 ( .C (clk), .D (signal_5591), .Q (signal_12881) ) ;
    buf_clk cell_7995 ( .C (clk), .D (signal_8880), .Q (signal_12883) ) ;
    buf_clk cell_7997 ( .C (clk), .D (signal_5497), .Q (signal_12885) ) ;
    buf_clk cell_7999 ( .C (clk), .D (signal_8783), .Q (signal_12887) ) ;
    buf_clk cell_8001 ( .C (clk), .D (signal_5592), .Q (signal_12889) ) ;
    buf_clk cell_8003 ( .C (clk), .D (signal_8881), .Q (signal_12891) ) ;
    buf_clk cell_8005 ( .C (clk), .D (signal_5593), .Q (signal_12893) ) ;
    buf_clk cell_8007 ( .C (clk), .D (signal_8882), .Q (signal_12895) ) ;
    buf_clk cell_8009 ( .C (clk), .D (signal_5501), .Q (signal_12897) ) ;
    buf_clk cell_8011 ( .C (clk), .D (signal_8787), .Q (signal_12899) ) ;
    buf_clk cell_8013 ( .C (clk), .D (signal_5594), .Q (signal_12901) ) ;
    buf_clk cell_8015 ( .C (clk), .D (signal_8883), .Q (signal_12903) ) ;
    buf_clk cell_8017 ( .C (clk), .D (signal_5595), .Q (signal_12905) ) ;
    buf_clk cell_8019 ( .C (clk), .D (signal_8884), .Q (signal_12907) ) ;
    buf_clk cell_8021 ( .C (clk), .D (signal_5505), .Q (signal_12909) ) ;
    buf_clk cell_8023 ( .C (clk), .D (signal_8791), .Q (signal_12911) ) ;
    buf_clk cell_8025 ( .C (clk), .D (signal_5596), .Q (signal_12913) ) ;
    buf_clk cell_8027 ( .C (clk), .D (signal_8885), .Q (signal_12915) ) ;
    buf_clk cell_8029 ( .C (clk), .D (signal_5597), .Q (signal_12917) ) ;
    buf_clk cell_8031 ( .C (clk), .D (signal_8886), .Q (signal_12919) ) ;
    buf_clk cell_8033 ( .C (clk), .D (signal_5509), .Q (signal_12921) ) ;
    buf_clk cell_8035 ( .C (clk), .D (signal_8795), .Q (signal_12923) ) ;
    buf_clk cell_8037 ( .C (clk), .D (signal_5598), .Q (signal_12925) ) ;
    buf_clk cell_8039 ( .C (clk), .D (signal_8887), .Q (signal_12927) ) ;
    buf_clk cell_8041 ( .C (clk), .D (signal_5599), .Q (signal_12929) ) ;
    buf_clk cell_8043 ( .C (clk), .D (signal_8888), .Q (signal_12931) ) ;
    buf_clk cell_8045 ( .C (clk), .D (signal_5513), .Q (signal_12933) ) ;
    buf_clk cell_8047 ( .C (clk), .D (signal_8799), .Q (signal_12935) ) ;
    buf_clk cell_8049 ( .C (clk), .D (signal_5600), .Q (signal_12937) ) ;
    buf_clk cell_8051 ( .C (clk), .D (signal_8889), .Q (signal_12939) ) ;
    buf_clk cell_8053 ( .C (clk), .D (signal_5601), .Q (signal_12941) ) ;
    buf_clk cell_8055 ( .C (clk), .D (signal_8890), .Q (signal_12943) ) ;
    buf_clk cell_8057 ( .C (clk), .D (signal_5517), .Q (signal_12945) ) ;
    buf_clk cell_8059 ( .C (clk), .D (signal_8803), .Q (signal_12947) ) ;
    buf_clk cell_8061 ( .C (clk), .D (signal_5602), .Q (signal_12949) ) ;
    buf_clk cell_8063 ( .C (clk), .D (signal_8891), .Q (signal_12951) ) ;
    buf_clk cell_8065 ( .C (clk), .D (signal_5603), .Q (signal_12953) ) ;
    buf_clk cell_8067 ( .C (clk), .D (signal_8892), .Q (signal_12955) ) ;
    buf_clk cell_8069 ( .C (clk), .D (signal_5604), .Q (signal_12957) ) ;
    buf_clk cell_8071 ( .C (clk), .D (signal_8924), .Q (signal_12959) ) ;
    buf_clk cell_8073 ( .C (clk), .D (signal_5523), .Q (signal_12961) ) ;
    buf_clk cell_8075 ( .C (clk), .D (signal_8807), .Q (signal_12963) ) ;
    buf_clk cell_8077 ( .C (clk), .D (signal_5608), .Q (signal_12965) ) ;
    buf_clk cell_8079 ( .C (clk), .D (signal_8893), .Q (signal_12967) ) ;
    buf_clk cell_8081 ( .C (clk), .D (signal_5609), .Q (signal_12969) ) ;
    buf_clk cell_8083 ( .C (clk), .D (signal_8894), .Q (signal_12971) ) ;
    buf_clk cell_8085 ( .C (clk), .D (signal_5527), .Q (signal_12973) ) ;
    buf_clk cell_8087 ( .C (clk), .D (signal_8811), .Q (signal_12975) ) ;
    buf_clk cell_8089 ( .C (clk), .D (signal_5610), .Q (signal_12977) ) ;
    buf_clk cell_8091 ( .C (clk), .D (signal_8895), .Q (signal_12979) ) ;
    buf_clk cell_8093 ( .C (clk), .D (signal_5611), .Q (signal_12981) ) ;
    buf_clk cell_8095 ( .C (clk), .D (signal_8896), .Q (signal_12983) ) ;
    buf_clk cell_8097 ( .C (clk), .D (signal_5531), .Q (signal_12985) ) ;
    buf_clk cell_8099 ( .C (clk), .D (signal_8815), .Q (signal_12987) ) ;
    buf_clk cell_8101 ( .C (clk), .D (signal_5612), .Q (signal_12989) ) ;
    buf_clk cell_8103 ( .C (clk), .D (signal_8897), .Q (signal_12991) ) ;
    buf_clk cell_8105 ( .C (clk), .D (signal_5613), .Q (signal_12993) ) ;
    buf_clk cell_8107 ( .C (clk), .D (signal_8898), .Q (signal_12995) ) ;
    buf_clk cell_8109 ( .C (clk), .D (signal_5614), .Q (signal_12997) ) ;
    buf_clk cell_8111 ( .C (clk), .D (signal_8928), .Q (signal_12999) ) ;
    buf_clk cell_8113 ( .C (clk), .D (signal_5537), .Q (signal_13001) ) ;
    buf_clk cell_8115 ( .C (clk), .D (signal_8819), .Q (signal_13003) ) ;
    buf_clk cell_8117 ( .C (clk), .D (signal_5618), .Q (signal_13005) ) ;
    buf_clk cell_8119 ( .C (clk), .D (signal_8899), .Q (signal_13007) ) ;
    buf_clk cell_8121 ( .C (clk), .D (signal_5619), .Q (signal_13009) ) ;
    buf_clk cell_8123 ( .C (clk), .D (signal_8900), .Q (signal_13011) ) ;
    buf_clk cell_8125 ( .C (clk), .D (signal_5541), .Q (signal_13013) ) ;
    buf_clk cell_8127 ( .C (clk), .D (signal_8823), .Q (signal_13015) ) ;
    buf_clk cell_8129 ( .C (clk), .D (signal_5620), .Q (signal_13017) ) ;
    buf_clk cell_8131 ( .C (clk), .D (signal_8901), .Q (signal_13019) ) ;
    buf_clk cell_8133 ( .C (clk), .D (signal_5621), .Q (signal_13021) ) ;
    buf_clk cell_8135 ( .C (clk), .D (signal_8902), .Q (signal_13023) ) ;
    buf_clk cell_8137 ( .C (clk), .D (signal_5545), .Q (signal_13025) ) ;
    buf_clk cell_8139 ( .C (clk), .D (signal_8827), .Q (signal_13027) ) ;
    buf_clk cell_8141 ( .C (clk), .D (signal_5622), .Q (signal_13029) ) ;
    buf_clk cell_8143 ( .C (clk), .D (signal_8903), .Q (signal_13031) ) ;
    buf_clk cell_8145 ( .C (clk), .D (signal_5623), .Q (signal_13033) ) ;
    buf_clk cell_8147 ( .C (clk), .D (signal_8904), .Q (signal_13035) ) ;
    buf_clk cell_8149 ( .C (clk), .D (signal_5624), .Q (signal_13037) ) ;
    buf_clk cell_8151 ( .C (clk), .D (signal_8932), .Q (signal_13039) ) ;
    buf_clk cell_8153 ( .C (clk), .D (signal_5628), .Q (signal_13041) ) ;
    buf_clk cell_8155 ( .C (clk), .D (signal_8905), .Q (signal_13043) ) ;
    buf_clk cell_8157 ( .C (clk), .D (signal_5632), .Q (signal_13045) ) ;
    buf_clk cell_8159 ( .C (clk), .D (signal_8909), .Q (signal_13047) ) ;
    buf_clk cell_8161 ( .C (clk), .D (signal_5636), .Q (signal_13049) ) ;
    buf_clk cell_8163 ( .C (clk), .D (signal_8913), .Q (signal_13051) ) ;
    buf_clk cell_8165 ( .C (clk), .D (signal_5640), .Q (signal_13053) ) ;
    buf_clk cell_8167 ( .C (clk), .D (signal_8917), .Q (signal_13055) ) ;
    buf_clk cell_8169 ( .C (clk), .D (signal_5685), .Q (signal_13057) ) ;
    buf_clk cell_8171 ( .C (clk), .D (signal_8965), .Q (signal_13059) ) ;
    buf_clk cell_8173 ( .C (clk), .D (signal_5689), .Q (signal_13061) ) ;
    buf_clk cell_8175 ( .C (clk), .D (signal_8969), .Q (signal_13063) ) ;
    buf_clk cell_8177 ( .C (clk), .D (signal_5693), .Q (signal_13065) ) ;
    buf_clk cell_8179 ( .C (clk), .D (signal_8973), .Q (signal_13067) ) ;
    buf_clk cell_8181 ( .C (clk), .D (signal_5697), .Q (signal_13069) ) ;
    buf_clk cell_8183 ( .C (clk), .D (signal_8977), .Q (signal_13071) ) ;
    buf_clk cell_8185 ( .C (clk), .D (signal_5701), .Q (signal_13073) ) ;
    buf_clk cell_8187 ( .C (clk), .D (signal_8981), .Q (signal_13075) ) ;
    buf_clk cell_8189 ( .C (clk), .D (signal_5705), .Q (signal_13077) ) ;
    buf_clk cell_8191 ( .C (clk), .D (signal_8985), .Q (signal_13079) ) ;
    buf_clk cell_8193 ( .C (clk), .D (signal_5709), .Q (signal_13081) ) ;
    buf_clk cell_8195 ( .C (clk), .D (signal_8989), .Q (signal_13083) ) ;
    buf_clk cell_8197 ( .C (clk), .D (signal_5714), .Q (signal_13085) ) ;
    buf_clk cell_8199 ( .C (clk), .D (signal_8993), .Q (signal_13087) ) ;
    buf_clk cell_8201 ( .C (clk), .D (signal_5718), .Q (signal_13089) ) ;
    buf_clk cell_8203 ( .C (clk), .D (signal_8997), .Q (signal_13091) ) ;
    buf_clk cell_8205 ( .C (clk), .D (signal_5722), .Q (signal_13093) ) ;
    buf_clk cell_8207 ( .C (clk), .D (signal_9001), .Q (signal_13095) ) ;
    buf_clk cell_8209 ( .C (clk), .D (signal_5727), .Q (signal_13097) ) ;
    buf_clk cell_8211 ( .C (clk), .D (signal_9005), .Q (signal_13099) ) ;
    buf_clk cell_8213 ( .C (clk), .D (signal_5731), .Q (signal_13101) ) ;
    buf_clk cell_8215 ( .C (clk), .D (signal_9009), .Q (signal_13103) ) ;
    buf_clk cell_8217 ( .C (clk), .D (signal_5735), .Q (signal_13105) ) ;
    buf_clk cell_8219 ( .C (clk), .D (signal_9013), .Q (signal_13107) ) ;
    buf_clk cell_8543 ( .C (clk), .D (signal_13430), .Q (signal_13431) ) ;
    buf_clk cell_8551 ( .C (clk), .D (signal_13438), .Q (signal_13439) ) ;
    buf_clk cell_8559 ( .C (clk), .D (signal_13446), .Q (signal_13447) ) ;
    buf_clk cell_8567 ( .C (clk), .D (signal_13454), .Q (signal_13455) ) ;
    buf_clk cell_8575 ( .C (clk), .D (signal_13462), .Q (signal_13463) ) ;
    buf_clk cell_8583 ( .C (clk), .D (signal_13470), .Q (signal_13471) ) ;
    buf_clk cell_8591 ( .C (clk), .D (signal_13478), .Q (signal_13479) ) ;
    buf_clk cell_8599 ( .C (clk), .D (signal_13486), .Q (signal_13487) ) ;
    buf_clk cell_8607 ( .C (clk), .D (signal_13494), .Q (signal_13495) ) ;
    buf_clk cell_8615 ( .C (clk), .D (signal_13502), .Q (signal_13503) ) ;
    buf_clk cell_8623 ( .C (clk), .D (signal_13510), .Q (signal_13511) ) ;
    buf_clk cell_8631 ( .C (clk), .D (signal_13518), .Q (signal_13519) ) ;
    buf_clk cell_8639 ( .C (clk), .D (signal_13526), .Q (signal_13527) ) ;
    buf_clk cell_8647 ( .C (clk), .D (signal_13534), .Q (signal_13535) ) ;
    buf_clk cell_8655 ( .C (clk), .D (signal_13542), .Q (signal_13543) ) ;
    buf_clk cell_8663 ( .C (clk), .D (signal_13550), .Q (signal_13551) ) ;
    buf_clk cell_8671 ( .C (clk), .D (signal_13558), .Q (signal_13559) ) ;
    buf_clk cell_8679 ( .C (clk), .D (signal_13566), .Q (signal_13567) ) ;
    buf_clk cell_8687 ( .C (clk), .D (signal_13574), .Q (signal_13575) ) ;
    buf_clk cell_8695 ( .C (clk), .D (signal_13582), .Q (signal_13583) ) ;
    buf_clk cell_8703 ( .C (clk), .D (signal_13590), .Q (signal_13591) ) ;
    buf_clk cell_8711 ( .C (clk), .D (signal_13598), .Q (signal_13599) ) ;
    buf_clk cell_8719 ( .C (clk), .D (signal_13606), .Q (signal_13607) ) ;
    buf_clk cell_8727 ( .C (clk), .D (signal_13614), .Q (signal_13615) ) ;
    buf_clk cell_8735 ( .C (clk), .D (signal_13622), .Q (signal_13623) ) ;
    buf_clk cell_8743 ( .C (clk), .D (signal_13630), .Q (signal_13631) ) ;
    buf_clk cell_8751 ( .C (clk), .D (signal_13638), .Q (signal_13639) ) ;
    buf_clk cell_8759 ( .C (clk), .D (signal_13646), .Q (signal_13647) ) ;
    buf_clk cell_8767 ( .C (clk), .D (signal_13654), .Q (signal_13655) ) ;
    buf_clk cell_8775 ( .C (clk), .D (signal_13662), .Q (signal_13663) ) ;
    buf_clk cell_8783 ( .C (clk), .D (signal_13670), .Q (signal_13671) ) ;
    buf_clk cell_8791 ( .C (clk), .D (signal_13678), .Q (signal_13679) ) ;
    buf_clk cell_8799 ( .C (clk), .D (signal_13686), .Q (signal_13687) ) ;
    buf_clk cell_8807 ( .C (clk), .D (signal_13694), .Q (signal_13695) ) ;
    buf_clk cell_8815 ( .C (clk), .D (signal_13702), .Q (signal_13703) ) ;
    buf_clk cell_8823 ( .C (clk), .D (signal_13710), .Q (signal_13711) ) ;
    buf_clk cell_8831 ( .C (clk), .D (signal_13718), .Q (signal_13719) ) ;
    buf_clk cell_8839 ( .C (clk), .D (signal_13726), .Q (signal_13727) ) ;
    buf_clk cell_8847 ( .C (clk), .D (signal_13734), .Q (signal_13735) ) ;
    buf_clk cell_8855 ( .C (clk), .D (signal_13742), .Q (signal_13743) ) ;
    buf_clk cell_8863 ( .C (clk), .D (signal_13750), .Q (signal_13751) ) ;
    buf_clk cell_8871 ( .C (clk), .D (signal_13758), .Q (signal_13759) ) ;
    buf_clk cell_8879 ( .C (clk), .D (signal_13766), .Q (signal_13767) ) ;
    buf_clk cell_8887 ( .C (clk), .D (signal_13774), .Q (signal_13775) ) ;
    buf_clk cell_8895 ( .C (clk), .D (signal_13782), .Q (signal_13783) ) ;
    buf_clk cell_8903 ( .C (clk), .D (signal_13790), .Q (signal_13791) ) ;
    buf_clk cell_8911 ( .C (clk), .D (signal_13798), .Q (signal_13799) ) ;
    buf_clk cell_8919 ( .C (clk), .D (signal_13806), .Q (signal_13807) ) ;
    buf_clk cell_8927 ( .C (clk), .D (signal_13814), .Q (signal_13815) ) ;
    buf_clk cell_8935 ( .C (clk), .D (signal_13822), .Q (signal_13823) ) ;
    buf_clk cell_8943 ( .C (clk), .D (signal_13830), .Q (signal_13831) ) ;
    buf_clk cell_8951 ( .C (clk), .D (signal_13838), .Q (signal_13839) ) ;
    buf_clk cell_8959 ( .C (clk), .D (signal_13846), .Q (signal_13847) ) ;
    buf_clk cell_8967 ( .C (clk), .D (signal_13854), .Q (signal_13855) ) ;
    buf_clk cell_8975 ( .C (clk), .D (signal_13862), .Q (signal_13863) ) ;
    buf_clk cell_8983 ( .C (clk), .D (signal_13870), .Q (signal_13871) ) ;
    buf_clk cell_8991 ( .C (clk), .D (signal_13878), .Q (signal_13879) ) ;
    buf_clk cell_8999 ( .C (clk), .D (signal_13886), .Q (signal_13887) ) ;
    buf_clk cell_9007 ( .C (clk), .D (signal_13894), .Q (signal_13895) ) ;
    buf_clk cell_9015 ( .C (clk), .D (signal_13902), .Q (signal_13903) ) ;
    buf_clk cell_9023 ( .C (clk), .D (signal_13910), .Q (signal_13911) ) ;
    buf_clk cell_9031 ( .C (clk), .D (signal_13918), .Q (signal_13919) ) ;
    buf_clk cell_9039 ( .C (clk), .D (signal_13926), .Q (signal_13927) ) ;
    buf_clk cell_9047 ( .C (clk), .D (signal_13934), .Q (signal_13935) ) ;
    buf_clk cell_9055 ( .C (clk), .D (signal_13942), .Q (signal_13943) ) ;
    buf_clk cell_9063 ( .C (clk), .D (signal_13950), .Q (signal_13951) ) ;
    buf_clk cell_9071 ( .C (clk), .D (signal_13958), .Q (signal_13959) ) ;
    buf_clk cell_9079 ( .C (clk), .D (signal_13966), .Q (signal_13967) ) ;
    buf_clk cell_9087 ( .C (clk), .D (signal_13974), .Q (signal_13975) ) ;
    buf_clk cell_9095 ( .C (clk), .D (signal_13982), .Q (signal_13983) ) ;
    buf_clk cell_9103 ( .C (clk), .D (signal_13990), .Q (signal_13991) ) ;
    buf_clk cell_9111 ( .C (clk), .D (signal_13998), .Q (signal_13999) ) ;
    buf_clk cell_9119 ( .C (clk), .D (signal_14006), .Q (signal_14007) ) ;
    buf_clk cell_9127 ( .C (clk), .D (signal_14014), .Q (signal_14015) ) ;
    buf_clk cell_9135 ( .C (clk), .D (signal_14022), .Q (signal_14023) ) ;
    buf_clk cell_9143 ( .C (clk), .D (signal_14030), .Q (signal_14031) ) ;
    buf_clk cell_9151 ( .C (clk), .D (signal_14038), .Q (signal_14039) ) ;
    buf_clk cell_9159 ( .C (clk), .D (signal_14046), .Q (signal_14047) ) ;
    buf_clk cell_9167 ( .C (clk), .D (signal_14054), .Q (signal_14055) ) ;
    buf_clk cell_9175 ( .C (clk), .D (signal_14062), .Q (signal_14063) ) ;
    buf_clk cell_9183 ( .C (clk), .D (signal_14070), .Q (signal_14071) ) ;
    buf_clk cell_9191 ( .C (clk), .D (signal_14078), .Q (signal_14079) ) ;
    buf_clk cell_9199 ( .C (clk), .D (signal_14086), .Q (signal_14087) ) ;
    buf_clk cell_9207 ( .C (clk), .D (signal_14094), .Q (signal_14095) ) ;
    buf_clk cell_9215 ( .C (clk), .D (signal_14102), .Q (signal_14103) ) ;
    buf_clk cell_9223 ( .C (clk), .D (signal_14110), .Q (signal_14111) ) ;
    buf_clk cell_9231 ( .C (clk), .D (signal_14118), .Q (signal_14119) ) ;
    buf_clk cell_9239 ( .C (clk), .D (signal_14126), .Q (signal_14127) ) ;
    buf_clk cell_9247 ( .C (clk), .D (signal_14134), .Q (signal_14135) ) ;
    buf_clk cell_9255 ( .C (clk), .D (signal_14142), .Q (signal_14143) ) ;
    buf_clk cell_9263 ( .C (clk), .D (signal_14150), .Q (signal_14151) ) ;
    buf_clk cell_9271 ( .C (clk), .D (signal_14158), .Q (signal_14159) ) ;
    buf_clk cell_9279 ( .C (clk), .D (signal_14166), .Q (signal_14167) ) ;
    buf_clk cell_9287 ( .C (clk), .D (signal_14174), .Q (signal_14175) ) ;
    buf_clk cell_9295 ( .C (clk), .D (signal_14182), .Q (signal_14183) ) ;
    buf_clk cell_9303 ( .C (clk), .D (signal_14190), .Q (signal_14191) ) ;
    buf_clk cell_9311 ( .C (clk), .D (signal_14198), .Q (signal_14199) ) ;
    buf_clk cell_9319 ( .C (clk), .D (signal_14206), .Q (signal_14207) ) ;
    buf_clk cell_9327 ( .C (clk), .D (signal_14214), .Q (signal_14215) ) ;
    buf_clk cell_9335 ( .C (clk), .D (signal_14222), .Q (signal_14223) ) ;
    buf_clk cell_9343 ( .C (clk), .D (signal_14230), .Q (signal_14231) ) ;
    buf_clk cell_9351 ( .C (clk), .D (signal_14238), .Q (signal_14239) ) ;
    buf_clk cell_9359 ( .C (clk), .D (signal_14246), .Q (signal_14247) ) ;
    buf_clk cell_9367 ( .C (clk), .D (signal_14254), .Q (signal_14255) ) ;
    buf_clk cell_9375 ( .C (clk), .D (signal_14262), .Q (signal_14263) ) ;
    buf_clk cell_9383 ( .C (clk), .D (signal_14270), .Q (signal_14271) ) ;
    buf_clk cell_9391 ( .C (clk), .D (signal_14278), .Q (signal_14279) ) ;
    buf_clk cell_9399 ( .C (clk), .D (signal_14286), .Q (signal_14287) ) ;
    buf_clk cell_9407 ( .C (clk), .D (signal_14294), .Q (signal_14295) ) ;
    buf_clk cell_9415 ( .C (clk), .D (signal_14302), .Q (signal_14303) ) ;
    buf_clk cell_9423 ( .C (clk), .D (signal_14310), .Q (signal_14311) ) ;
    buf_clk cell_9431 ( .C (clk), .D (signal_14318), .Q (signal_14319) ) ;
    buf_clk cell_9439 ( .C (clk), .D (signal_14326), .Q (signal_14327) ) ;
    buf_clk cell_9447 ( .C (clk), .D (signal_14334), .Q (signal_14335) ) ;
    buf_clk cell_9455 ( .C (clk), .D (signal_14342), .Q (signal_14343) ) ;
    buf_clk cell_9463 ( .C (clk), .D (signal_14350), .Q (signal_14351) ) ;
    buf_clk cell_9471 ( .C (clk), .D (signal_14358), .Q (signal_14359) ) ;
    buf_clk cell_9479 ( .C (clk), .D (signal_14366), .Q (signal_14367) ) ;
    buf_clk cell_9487 ( .C (clk), .D (signal_14374), .Q (signal_14375) ) ;
    buf_clk cell_9495 ( .C (clk), .D (signal_14382), .Q (signal_14383) ) ;
    buf_clk cell_9503 ( .C (clk), .D (signal_14390), .Q (signal_14391) ) ;
    buf_clk cell_9511 ( .C (clk), .D (signal_14398), .Q (signal_14399) ) ;
    buf_clk cell_9519 ( .C (clk), .D (signal_14406), .Q (signal_14407) ) ;
    buf_clk cell_9527 ( .C (clk), .D (signal_14414), .Q (signal_14415) ) ;
    buf_clk cell_9535 ( .C (clk), .D (signal_14422), .Q (signal_14423) ) ;
    buf_clk cell_9543 ( .C (clk), .D (signal_14430), .Q (signal_14431) ) ;
    buf_clk cell_9551 ( .C (clk), .D (signal_14438), .Q (signal_14439) ) ;
    buf_clk cell_9559 ( .C (clk), .D (signal_14446), .Q (signal_14447) ) ;
    buf_clk cell_9567 ( .C (clk), .D (signal_14454), .Q (signal_14455) ) ;
    buf_clk cell_9575 ( .C (clk), .D (signal_14462), .Q (signal_14463) ) ;
    buf_clk cell_9583 ( .C (clk), .D (signal_14470), .Q (signal_14471) ) ;
    buf_clk cell_9591 ( .C (clk), .D (signal_14478), .Q (signal_14479) ) ;
    buf_clk cell_9599 ( .C (clk), .D (signal_14486), .Q (signal_14487) ) ;
    buf_clk cell_9607 ( .C (clk), .D (signal_14494), .Q (signal_14495) ) ;
    buf_clk cell_9615 ( .C (clk), .D (signal_14502), .Q (signal_14503) ) ;
    buf_clk cell_9623 ( .C (clk), .D (signal_14510), .Q (signal_14511) ) ;
    buf_clk cell_9631 ( .C (clk), .D (signal_14518), .Q (signal_14519) ) ;
    buf_clk cell_9639 ( .C (clk), .D (signal_14526), .Q (signal_14527) ) ;
    buf_clk cell_9647 ( .C (clk), .D (signal_14534), .Q (signal_14535) ) ;
    buf_clk cell_9655 ( .C (clk), .D (signal_14542), .Q (signal_14543) ) ;
    buf_clk cell_9663 ( .C (clk), .D (signal_14550), .Q (signal_14551) ) ;
    buf_clk cell_9671 ( .C (clk), .D (signal_14558), .Q (signal_14559) ) ;
    buf_clk cell_9679 ( .C (clk), .D (signal_14566), .Q (signal_14567) ) ;
    buf_clk cell_9687 ( .C (clk), .D (signal_14574), .Q (signal_14575) ) ;
    buf_clk cell_9695 ( .C (clk), .D (signal_14582), .Q (signal_14583) ) ;
    buf_clk cell_9703 ( .C (clk), .D (signal_14590), .Q (signal_14591) ) ;
    buf_clk cell_9711 ( .C (clk), .D (signal_14598), .Q (signal_14599) ) ;
    buf_clk cell_9719 ( .C (clk), .D (signal_14606), .Q (signal_14607) ) ;
    buf_clk cell_9727 ( .C (clk), .D (signal_14614), .Q (signal_14615) ) ;
    buf_clk cell_9735 ( .C (clk), .D (signal_14622), .Q (signal_14623) ) ;
    buf_clk cell_9743 ( .C (clk), .D (signal_14630), .Q (signal_14631) ) ;
    buf_clk cell_9751 ( .C (clk), .D (signal_14638), .Q (signal_14639) ) ;
    buf_clk cell_9759 ( .C (clk), .D (signal_14646), .Q (signal_14647) ) ;
    buf_clk cell_9767 ( .C (clk), .D (signal_14654), .Q (signal_14655) ) ;
    buf_clk cell_9775 ( .C (clk), .D (signal_14662), .Q (signal_14663) ) ;
    buf_clk cell_9783 ( .C (clk), .D (signal_14670), .Q (signal_14671) ) ;
    buf_clk cell_9791 ( .C (clk), .D (signal_14678), .Q (signal_14679) ) ;
    buf_clk cell_9799 ( .C (clk), .D (signal_14686), .Q (signal_14687) ) ;
    buf_clk cell_9807 ( .C (clk), .D (signal_14694), .Q (signal_14695) ) ;
    buf_clk cell_9815 ( .C (clk), .D (signal_14702), .Q (signal_14703) ) ;
    buf_clk cell_9823 ( .C (clk), .D (signal_14710), .Q (signal_14711) ) ;
    buf_clk cell_9831 ( .C (clk), .D (signal_14718), .Q (signal_14719) ) ;
    buf_clk cell_9839 ( .C (clk), .D (signal_14726), .Q (signal_14727) ) ;
    buf_clk cell_9847 ( .C (clk), .D (signal_14734), .Q (signal_14735) ) ;
    buf_clk cell_9855 ( .C (clk), .D (signal_14742), .Q (signal_14743) ) ;
    buf_clk cell_9863 ( .C (clk), .D (signal_14750), .Q (signal_14751) ) ;
    buf_clk cell_9871 ( .C (clk), .D (signal_14758), .Q (signal_14759) ) ;
    buf_clk cell_9879 ( .C (clk), .D (signal_14766), .Q (signal_14767) ) ;
    buf_clk cell_9887 ( .C (clk), .D (signal_14774), .Q (signal_14775) ) ;
    buf_clk cell_9895 ( .C (clk), .D (signal_14782), .Q (signal_14783) ) ;
    buf_clk cell_9903 ( .C (clk), .D (signal_14790), .Q (signal_14791) ) ;
    buf_clk cell_9911 ( .C (clk), .D (signal_14798), .Q (signal_14799) ) ;
    buf_clk cell_9919 ( .C (clk), .D (signal_14806), .Q (signal_14807) ) ;
    buf_clk cell_9927 ( .C (clk), .D (signal_14814), .Q (signal_14815) ) ;
    buf_clk cell_9935 ( .C (clk), .D (signal_14822), .Q (signal_14823) ) ;
    buf_clk cell_9943 ( .C (clk), .D (signal_14830), .Q (signal_14831) ) ;
    buf_clk cell_9951 ( .C (clk), .D (signal_14838), .Q (signal_14839) ) ;
    buf_clk cell_9959 ( .C (clk), .D (signal_14846), .Q (signal_14847) ) ;
    buf_clk cell_9967 ( .C (clk), .D (signal_14854), .Q (signal_14855) ) ;
    buf_clk cell_9975 ( .C (clk), .D (signal_14862), .Q (signal_14863) ) ;
    buf_clk cell_9983 ( .C (clk), .D (signal_14870), .Q (signal_14871) ) ;
    buf_clk cell_9991 ( .C (clk), .D (signal_14878), .Q (signal_14879) ) ;
    buf_clk cell_9999 ( .C (clk), .D (signal_14886), .Q (signal_14887) ) ;
    buf_clk cell_10007 ( .C (clk), .D (signal_14894), .Q (signal_14895) ) ;
    buf_clk cell_10015 ( .C (clk), .D (signal_14902), .Q (signal_14903) ) ;
    buf_clk cell_10023 ( .C (clk), .D (signal_14910), .Q (signal_14911) ) ;
    buf_clk cell_10031 ( .C (clk), .D (signal_14918), .Q (signal_14919) ) ;
    buf_clk cell_10039 ( .C (clk), .D (signal_14926), .Q (signal_14927) ) ;
    buf_clk cell_10047 ( .C (clk), .D (signal_14934), .Q (signal_14935) ) ;
    buf_clk cell_10055 ( .C (clk), .D (signal_14942), .Q (signal_14943) ) ;
    buf_clk cell_10063 ( .C (clk), .D (signal_14950), .Q (signal_14951) ) ;
    buf_clk cell_10071 ( .C (clk), .D (signal_14958), .Q (signal_14959) ) ;
    buf_clk cell_10079 ( .C (clk), .D (signal_14966), .Q (signal_14967) ) ;
    buf_clk cell_10087 ( .C (clk), .D (signal_14974), .Q (signal_14975) ) ;
    buf_clk cell_10095 ( .C (clk), .D (signal_14982), .Q (signal_14983) ) ;
    buf_clk cell_10103 ( .C (clk), .D (signal_14990), .Q (signal_14991) ) ;
    buf_clk cell_10111 ( .C (clk), .D (signal_14998), .Q (signal_14999) ) ;
    buf_clk cell_10119 ( .C (clk), .D (signal_15006), .Q (signal_15007) ) ;
    buf_clk cell_10127 ( .C (clk), .D (signal_15014), .Q (signal_15015) ) ;
    buf_clk cell_10135 ( .C (clk), .D (signal_15022), .Q (signal_15023) ) ;
    buf_clk cell_10143 ( .C (clk), .D (signal_15030), .Q (signal_15031) ) ;
    buf_clk cell_10151 ( .C (clk), .D (signal_15038), .Q (signal_15039) ) ;
    buf_clk cell_10159 ( .C (clk), .D (signal_15046), .Q (signal_15047) ) ;
    buf_clk cell_10167 ( .C (clk), .D (signal_15054), .Q (signal_15055) ) ;
    buf_clk cell_10175 ( .C (clk), .D (signal_15062), .Q (signal_15063) ) ;
    buf_clk cell_10183 ( .C (clk), .D (signal_15070), .Q (signal_15071) ) ;
    buf_clk cell_10191 ( .C (clk), .D (signal_15078), .Q (signal_15079) ) ;
    buf_clk cell_10199 ( .C (clk), .D (signal_15086), .Q (signal_15087) ) ;
    buf_clk cell_10207 ( .C (clk), .D (signal_15094), .Q (signal_15095) ) ;
    buf_clk cell_10215 ( .C (clk), .D (signal_15102), .Q (signal_15103) ) ;
    buf_clk cell_10223 ( .C (clk), .D (signal_15110), .Q (signal_15111) ) ;
    buf_clk cell_10231 ( .C (clk), .D (signal_15118), .Q (signal_15119) ) ;
    buf_clk cell_10239 ( .C (clk), .D (signal_15126), .Q (signal_15127) ) ;
    buf_clk cell_10247 ( .C (clk), .D (signal_15134), .Q (signal_15135) ) ;
    buf_clk cell_10255 ( .C (clk), .D (signal_15142), .Q (signal_15143) ) ;
    buf_clk cell_10263 ( .C (clk), .D (signal_15150), .Q (signal_15151) ) ;
    buf_clk cell_10271 ( .C (clk), .D (signal_15158), .Q (signal_15159) ) ;
    buf_clk cell_10279 ( .C (clk), .D (signal_15166), .Q (signal_15167) ) ;
    buf_clk cell_10287 ( .C (clk), .D (signal_15174), .Q (signal_15175) ) ;
    buf_clk cell_10295 ( .C (clk), .D (signal_15182), .Q (signal_15183) ) ;
    buf_clk cell_10303 ( .C (clk), .D (signal_15190), .Q (signal_15191) ) ;
    buf_clk cell_10311 ( .C (clk), .D (signal_15198), .Q (signal_15199) ) ;
    buf_clk cell_10319 ( .C (clk), .D (signal_15206), .Q (signal_15207) ) ;
    buf_clk cell_10327 ( .C (clk), .D (signal_15214), .Q (signal_15215) ) ;
    buf_clk cell_10335 ( .C (clk), .D (signal_15222), .Q (signal_15223) ) ;
    buf_clk cell_10343 ( .C (clk), .D (signal_15230), .Q (signal_15231) ) ;
    buf_clk cell_10351 ( .C (clk), .D (signal_15238), .Q (signal_15239) ) ;
    buf_clk cell_10359 ( .C (clk), .D (signal_15246), .Q (signal_15247) ) ;
    buf_clk cell_10367 ( .C (clk), .D (signal_15254), .Q (signal_15255) ) ;
    buf_clk cell_10375 ( .C (clk), .D (signal_15262), .Q (signal_15263) ) ;
    buf_clk cell_10383 ( .C (clk), .D (signal_15270), .Q (signal_15271) ) ;
    buf_clk cell_10391 ( .C (clk), .D (signal_15278), .Q (signal_15279) ) ;
    buf_clk cell_10399 ( .C (clk), .D (signal_15286), .Q (signal_15287) ) ;
    buf_clk cell_10407 ( .C (clk), .D (signal_15294), .Q (signal_15295) ) ;
    buf_clk cell_10415 ( .C (clk), .D (signal_15302), .Q (signal_15303) ) ;
    buf_clk cell_10423 ( .C (clk), .D (signal_15310), .Q (signal_15311) ) ;
    buf_clk cell_10431 ( .C (clk), .D (signal_15318), .Q (signal_15319) ) ;
    buf_clk cell_10439 ( .C (clk), .D (signal_15326), .Q (signal_15327) ) ;
    buf_clk cell_10447 ( .C (clk), .D (signal_15334), .Q (signal_15335) ) ;
    buf_clk cell_10455 ( .C (clk), .D (signal_15342), .Q (signal_15343) ) ;
    buf_clk cell_10463 ( .C (clk), .D (signal_15350), .Q (signal_15351) ) ;
    buf_clk cell_10471 ( .C (clk), .D (signal_15358), .Q (signal_15359) ) ;
    buf_clk cell_10479 ( .C (clk), .D (signal_15366), .Q (signal_15367) ) ;
    buf_clk cell_10487 ( .C (clk), .D (signal_15374), .Q (signal_15375) ) ;
    buf_clk cell_10495 ( .C (clk), .D (signal_15382), .Q (signal_15383) ) ;
    buf_clk cell_10503 ( .C (clk), .D (signal_15390), .Q (signal_15391) ) ;
    buf_clk cell_10511 ( .C (clk), .D (signal_15398), .Q (signal_15399) ) ;
    buf_clk cell_10519 ( .C (clk), .D (signal_15406), .Q (signal_15407) ) ;
    buf_clk cell_10527 ( .C (clk), .D (signal_15414), .Q (signal_15415) ) ;
    buf_clk cell_10535 ( .C (clk), .D (signal_15422), .Q (signal_15423) ) ;
    buf_clk cell_10543 ( .C (clk), .D (signal_15430), .Q (signal_15431) ) ;
    buf_clk cell_10551 ( .C (clk), .D (signal_15438), .Q (signal_15439) ) ;
    buf_clk cell_10559 ( .C (clk), .D (signal_15446), .Q (signal_15447) ) ;
    buf_clk cell_10567 ( .C (clk), .D (signal_15454), .Q (signal_15455) ) ;
    buf_clk cell_10575 ( .C (clk), .D (signal_15462), .Q (signal_15463) ) ;
    buf_clk cell_10583 ( .C (clk), .D (signal_15470), .Q (signal_15471) ) ;
    buf_clk cell_10591 ( .C (clk), .D (signal_15478), .Q (signal_15479) ) ;
    buf_clk cell_10599 ( .C (clk), .D (signal_15486), .Q (signal_15487) ) ;
    buf_clk cell_10607 ( .C (clk), .D (signal_15494), .Q (signal_15495) ) ;
    buf_clk cell_10615 ( .C (clk), .D (signal_15502), .Q (signal_15503) ) ;
    buf_clk cell_10623 ( .C (clk), .D (signal_15510), .Q (signal_15511) ) ;
    buf_clk cell_10631 ( .C (clk), .D (signal_15518), .Q (signal_15519) ) ;
    buf_clk cell_10639 ( .C (clk), .D (signal_15526), .Q (signal_15527) ) ;
    buf_clk cell_10647 ( .C (clk), .D (signal_15534), .Q (signal_15535) ) ;
    buf_clk cell_10655 ( .C (clk), .D (signal_15542), .Q (signal_15543) ) ;
    buf_clk cell_10663 ( .C (clk), .D (signal_15550), .Q (signal_15551) ) ;
    buf_clk cell_10671 ( .C (clk), .D (signal_15558), .Q (signal_15559) ) ;
    buf_clk cell_10679 ( .C (clk), .D (signal_15566), .Q (signal_15567) ) ;
    buf_clk cell_10687 ( .C (clk), .D (signal_15574), .Q (signal_15575) ) ;
    buf_clk cell_10695 ( .C (clk), .D (signal_15582), .Q (signal_15583) ) ;
    buf_clk cell_10703 ( .C (clk), .D (signal_15590), .Q (signal_15591) ) ;
    buf_clk cell_10711 ( .C (clk), .D (signal_15598), .Q (signal_15599) ) ;
    buf_clk cell_10719 ( .C (clk), .D (signal_15606), .Q (signal_15607) ) ;
    buf_clk cell_10727 ( .C (clk), .D (signal_15614), .Q (signal_15615) ) ;
    buf_clk cell_10735 ( .C (clk), .D (signal_15622), .Q (signal_15623) ) ;
    buf_clk cell_10743 ( .C (clk), .D (signal_15630), .Q (signal_15631) ) ;
    buf_clk cell_10751 ( .C (clk), .D (signal_15638), .Q (signal_15639) ) ;
    buf_clk cell_10759 ( .C (clk), .D (signal_15646), .Q (signal_15647) ) ;
    buf_clk cell_10767 ( .C (clk), .D (signal_15654), .Q (signal_15655) ) ;
    buf_clk cell_10775 ( .C (clk), .D (signal_15662), .Q (signal_15663) ) ;
    buf_clk cell_10783 ( .C (clk), .D (signal_15670), .Q (signal_15671) ) ;
    buf_clk cell_10791 ( .C (clk), .D (signal_15678), .Q (signal_15679) ) ;
    buf_clk cell_10799 ( .C (clk), .D (signal_15686), .Q (signal_15687) ) ;
    buf_clk cell_10807 ( .C (clk), .D (signal_15694), .Q (signal_15695) ) ;
    buf_clk cell_10815 ( .C (clk), .D (signal_15702), .Q (signal_15703) ) ;
    buf_clk cell_10823 ( .C (clk), .D (signal_15710), .Q (signal_15711) ) ;
    buf_clk cell_10831 ( .C (clk), .D (signal_15718), .Q (signal_15719) ) ;
    buf_clk cell_10839 ( .C (clk), .D (signal_15726), .Q (signal_15727) ) ;
    buf_clk cell_10847 ( .C (clk), .D (signal_15734), .Q (signal_15735) ) ;
    buf_clk cell_10855 ( .C (clk), .D (signal_15742), .Q (signal_15743) ) ;
    buf_clk cell_10863 ( .C (clk), .D (signal_15750), .Q (signal_15751) ) ;
    buf_clk cell_10871 ( .C (clk), .D (signal_15758), .Q (signal_15759) ) ;
    buf_clk cell_10879 ( .C (clk), .D (signal_15766), .Q (signal_15767) ) ;
    buf_clk cell_10887 ( .C (clk), .D (signal_15774), .Q (signal_15775) ) ;
    buf_clk cell_10895 ( .C (clk), .D (signal_15782), .Q (signal_15783) ) ;
    buf_clk cell_10903 ( .C (clk), .D (signal_15790), .Q (signal_15791) ) ;
    buf_clk cell_10911 ( .C (clk), .D (signal_15798), .Q (signal_15799) ) ;
    buf_clk cell_10919 ( .C (clk), .D (signal_15806), .Q (signal_15807) ) ;
    buf_clk cell_10927 ( .C (clk), .D (signal_15814), .Q (signal_15815) ) ;
    buf_clk cell_10935 ( .C (clk), .D (signal_15822), .Q (signal_15823) ) ;
    buf_clk cell_10943 ( .C (clk), .D (signal_15830), .Q (signal_15831) ) ;
    buf_clk cell_10951 ( .C (clk), .D (signal_15838), .Q (signal_15839) ) ;
    buf_clk cell_10959 ( .C (clk), .D (signal_15846), .Q (signal_15847) ) ;
    buf_clk cell_10967 ( .C (clk), .D (signal_15854), .Q (signal_15855) ) ;
    buf_clk cell_10975 ( .C (clk), .D (signal_15862), .Q (signal_15863) ) ;
    buf_clk cell_10983 ( .C (clk), .D (signal_15870), .Q (signal_15871) ) ;
    buf_clk cell_10991 ( .C (clk), .D (signal_15878), .Q (signal_15879) ) ;
    buf_clk cell_10999 ( .C (clk), .D (signal_15886), .Q (signal_15887) ) ;
    buf_clk cell_11007 ( .C (clk), .D (signal_15894), .Q (signal_15895) ) ;
    buf_clk cell_11015 ( .C (clk), .D (signal_15902), .Q (signal_15903) ) ;
    buf_clk cell_11023 ( .C (clk), .D (signal_15910), .Q (signal_15911) ) ;
    buf_clk cell_11031 ( .C (clk), .D (signal_15918), .Q (signal_15919) ) ;
    buf_clk cell_11039 ( .C (clk), .D (signal_15926), .Q (signal_15927) ) ;
    buf_clk cell_11047 ( .C (clk), .D (signal_15934), .Q (signal_15935) ) ;
    buf_clk cell_11055 ( .C (clk), .D (signal_15942), .Q (signal_15943) ) ;
    buf_clk cell_11063 ( .C (clk), .D (signal_15950), .Q (signal_15951) ) ;
    buf_clk cell_11071 ( .C (clk), .D (signal_15958), .Q (signal_15959) ) ;
    buf_clk cell_11079 ( .C (clk), .D (signal_15966), .Q (signal_15967) ) ;
    buf_clk cell_11087 ( .C (clk), .D (signal_15974), .Q (signal_15975) ) ;
    buf_clk cell_11095 ( .C (clk), .D (signal_15982), .Q (signal_15983) ) ;
    buf_clk cell_11103 ( .C (clk), .D (signal_15990), .Q (signal_15991) ) ;
    buf_clk cell_11111 ( .C (clk), .D (signal_15998), .Q (signal_15999) ) ;
    buf_clk cell_11119 ( .C (clk), .D (signal_16006), .Q (signal_16007) ) ;
    buf_clk cell_11127 ( .C (clk), .D (signal_16014), .Q (signal_16015) ) ;
    buf_clk cell_11135 ( .C (clk), .D (signal_16022), .Q (signal_16023) ) ;
    buf_clk cell_11143 ( .C (clk), .D (signal_16030), .Q (signal_16031) ) ;
    buf_clk cell_11151 ( .C (clk), .D (signal_16038), .Q (signal_16039) ) ;
    buf_clk cell_11159 ( .C (clk), .D (signal_16046), .Q (signal_16047) ) ;
    buf_clk cell_11167 ( .C (clk), .D (signal_16054), .Q (signal_16055) ) ;
    buf_clk cell_11175 ( .C (clk), .D (signal_16062), .Q (signal_16063) ) ;
    buf_clk cell_11183 ( .C (clk), .D (signal_16070), .Q (signal_16071) ) ;
    buf_clk cell_11191 ( .C (clk), .D (signal_16078), .Q (signal_16079) ) ;
    buf_clk cell_11199 ( .C (clk), .D (signal_16086), .Q (signal_16087) ) ;
    buf_clk cell_11207 ( .C (clk), .D (signal_16094), .Q (signal_16095) ) ;
    buf_clk cell_11215 ( .C (clk), .D (signal_16102), .Q (signal_16103) ) ;
    buf_clk cell_11223 ( .C (clk), .D (signal_16110), .Q (signal_16111) ) ;
    buf_clk cell_11231 ( .C (clk), .D (signal_16118), .Q (signal_16119) ) ;
    buf_clk cell_11239 ( .C (clk), .D (signal_16126), .Q (signal_16127) ) ;
    buf_clk cell_11247 ( .C (clk), .D (signal_16134), .Q (signal_16135) ) ;
    buf_clk cell_11255 ( .C (clk), .D (signal_16142), .Q (signal_16143) ) ;
    buf_clk cell_11263 ( .C (clk), .D (signal_16150), .Q (signal_16151) ) ;
    buf_clk cell_11271 ( .C (clk), .D (signal_16158), .Q (signal_16159) ) ;
    buf_clk cell_11279 ( .C (clk), .D (signal_16166), .Q (signal_16167) ) ;
    buf_clk cell_11287 ( .C (clk), .D (signal_16174), .Q (signal_16175) ) ;
    buf_clk cell_11295 ( .C (clk), .D (signal_16182), .Q (signal_16183) ) ;
    buf_clk cell_11303 ( .C (clk), .D (signal_16190), .Q (signal_16191) ) ;
    buf_clk cell_11311 ( .C (clk), .D (signal_16198), .Q (signal_16199) ) ;
    buf_clk cell_11319 ( .C (clk), .D (signal_16206), .Q (signal_16207) ) ;
    buf_clk cell_11327 ( .C (clk), .D (signal_16214), .Q (signal_16215) ) ;
    buf_clk cell_11335 ( .C (clk), .D (signal_16222), .Q (signal_16223) ) ;
    buf_clk cell_11343 ( .C (clk), .D (signal_16230), .Q (signal_16231) ) ;
    buf_clk cell_11351 ( .C (clk), .D (signal_16238), .Q (signal_16239) ) ;
    buf_clk cell_11359 ( .C (clk), .D (signal_16246), .Q (signal_16247) ) ;
    buf_clk cell_11367 ( .C (clk), .D (signal_16254), .Q (signal_16255) ) ;
    buf_clk cell_11375 ( .C (clk), .D (signal_16262), .Q (signal_16263) ) ;
    buf_clk cell_11383 ( .C (clk), .D (signal_16270), .Q (signal_16271) ) ;
    buf_clk cell_11391 ( .C (clk), .D (signal_16278), .Q (signal_16279) ) ;
    buf_clk cell_11399 ( .C (clk), .D (signal_16286), .Q (signal_16287) ) ;
    buf_clk cell_11407 ( .C (clk), .D (signal_16294), .Q (signal_16295) ) ;
    buf_clk cell_11415 ( .C (clk), .D (signal_16302), .Q (signal_16303) ) ;
    buf_clk cell_11423 ( .C (clk), .D (signal_16310), .Q (signal_16311) ) ;
    buf_clk cell_11431 ( .C (clk), .D (signal_16318), .Q (signal_16319) ) ;
    buf_clk cell_11439 ( .C (clk), .D (signal_16326), .Q (signal_16327) ) ;
    buf_clk cell_11447 ( .C (clk), .D (signal_16334), .Q (signal_16335) ) ;
    buf_clk cell_11455 ( .C (clk), .D (signal_16342), .Q (signal_16343) ) ;
    buf_clk cell_11463 ( .C (clk), .D (signal_16350), .Q (signal_16351) ) ;
    buf_clk cell_11471 ( .C (clk), .D (signal_16358), .Q (signal_16359) ) ;
    buf_clk cell_11479 ( .C (clk), .D (signal_16366), .Q (signal_16367) ) ;
    buf_clk cell_11487 ( .C (clk), .D (signal_16374), .Q (signal_16375) ) ;
    buf_clk cell_11495 ( .C (clk), .D (signal_16382), .Q (signal_16383) ) ;
    buf_clk cell_11503 ( .C (clk), .D (signal_16390), .Q (signal_16391) ) ;
    buf_clk cell_11511 ( .C (clk), .D (signal_16398), .Q (signal_16399) ) ;
    buf_clk cell_11519 ( .C (clk), .D (signal_16406), .Q (signal_16407) ) ;
    buf_clk cell_11527 ( .C (clk), .D (signal_16414), .Q (signal_16415) ) ;
    buf_clk cell_11535 ( .C (clk), .D (signal_16422), .Q (signal_16423) ) ;
    buf_clk cell_11543 ( .C (clk), .D (signal_16430), .Q (signal_16431) ) ;
    buf_clk cell_11551 ( .C (clk), .D (signal_16438), .Q (signal_16439) ) ;
    buf_clk cell_11559 ( .C (clk), .D (signal_16446), .Q (signal_16447) ) ;
    buf_clk cell_11567 ( .C (clk), .D (signal_16454), .Q (signal_16455) ) ;
    buf_clk cell_11575 ( .C (clk), .D (signal_16462), .Q (signal_16463) ) ;
    buf_clk cell_11583 ( .C (clk), .D (signal_16470), .Q (signal_16471) ) ;
    buf_clk cell_11591 ( .C (clk), .D (signal_16478), .Q (signal_16479) ) ;
    buf_clk cell_11599 ( .C (clk), .D (signal_16486), .Q (signal_16487) ) ;
    buf_clk cell_11607 ( .C (clk), .D (signal_16494), .Q (signal_16495) ) ;
    buf_clk cell_11615 ( .C (clk), .D (signal_16502), .Q (signal_16503) ) ;
    buf_clk cell_11623 ( .C (clk), .D (signal_16510), .Q (signal_16511) ) ;
    buf_clk cell_11631 ( .C (clk), .D (signal_16518), .Q (signal_16519) ) ;
    buf_clk cell_11639 ( .C (clk), .D (signal_16526), .Q (signal_16527) ) ;
    buf_clk cell_11647 ( .C (clk), .D (signal_16534), .Q (signal_16535) ) ;
    buf_clk cell_11655 ( .C (clk), .D (signal_16542), .Q (signal_16543) ) ;
    buf_clk cell_11663 ( .C (clk), .D (signal_16550), .Q (signal_16551) ) ;
    buf_clk cell_11671 ( .C (clk), .D (signal_16558), .Q (signal_16559) ) ;
    buf_clk cell_11679 ( .C (clk), .D (signal_16566), .Q (signal_16567) ) ;
    buf_clk cell_11687 ( .C (clk), .D (signal_16574), .Q (signal_16575) ) ;
    buf_clk cell_11695 ( .C (clk), .D (signal_16582), .Q (signal_16583) ) ;
    buf_clk cell_11703 ( .C (clk), .D (signal_16590), .Q (signal_16591) ) ;
    buf_clk cell_11711 ( .C (clk), .D (signal_16598), .Q (signal_16599) ) ;
    buf_clk cell_11719 ( .C (clk), .D (signal_16606), .Q (signal_16607) ) ;
    buf_clk cell_11727 ( .C (clk), .D (signal_16614), .Q (signal_16615) ) ;
    buf_clk cell_11735 ( .C (clk), .D (signal_16622), .Q (signal_16623) ) ;
    buf_clk cell_11743 ( .C (clk), .D (signal_16630), .Q (signal_16631) ) ;
    buf_clk cell_11751 ( .C (clk), .D (signal_16638), .Q (signal_16639) ) ;
    buf_clk cell_11759 ( .C (clk), .D (signal_16646), .Q (signal_16647) ) ;
    buf_clk cell_11767 ( .C (clk), .D (signal_16654), .Q (signal_16655) ) ;
    buf_clk cell_11775 ( .C (clk), .D (signal_16662), .Q (signal_16663) ) ;
    buf_clk cell_11783 ( .C (clk), .D (signal_16670), .Q (signal_16671) ) ;
    buf_clk cell_11791 ( .C (clk), .D (signal_16678), .Q (signal_16679) ) ;
    buf_clk cell_11799 ( .C (clk), .D (signal_16686), .Q (signal_16687) ) ;
    buf_clk cell_11807 ( .C (clk), .D (signal_16694), .Q (signal_16695) ) ;
    buf_clk cell_11815 ( .C (clk), .D (signal_16702), .Q (signal_16703) ) ;
    buf_clk cell_11823 ( .C (clk), .D (signal_16710), .Q (signal_16711) ) ;
    buf_clk cell_11831 ( .C (clk), .D (signal_16718), .Q (signal_16719) ) ;
    buf_clk cell_11839 ( .C (clk), .D (signal_16726), .Q (signal_16727) ) ;
    buf_clk cell_11847 ( .C (clk), .D (signal_16734), .Q (signal_16735) ) ;
    buf_clk cell_11855 ( .C (clk), .D (signal_16742), .Q (signal_16743) ) ;
    buf_clk cell_11863 ( .C (clk), .D (signal_16750), .Q (signal_16751) ) ;
    buf_clk cell_11871 ( .C (clk), .D (signal_16758), .Q (signal_16759) ) ;
    buf_clk cell_11879 ( .C (clk), .D (signal_16766), .Q (signal_16767) ) ;
    buf_clk cell_11887 ( .C (clk), .D (signal_16774), .Q (signal_16775) ) ;
    buf_clk cell_11895 ( .C (clk), .D (signal_16782), .Q (signal_16783) ) ;
    buf_clk cell_11903 ( .C (clk), .D (signal_16790), .Q (signal_16791) ) ;
    buf_clk cell_11911 ( .C (clk), .D (signal_16798), .Q (signal_16799) ) ;
    buf_clk cell_11919 ( .C (clk), .D (signal_16806), .Q (signal_16807) ) ;
    buf_clk cell_11927 ( .C (clk), .D (signal_16814), .Q (signal_16815) ) ;
    buf_clk cell_11935 ( .C (clk), .D (signal_16822), .Q (signal_16823) ) ;
    buf_clk cell_11943 ( .C (clk), .D (signal_16830), .Q (signal_16831) ) ;
    buf_clk cell_11951 ( .C (clk), .D (signal_16838), .Q (signal_16839) ) ;
    buf_clk cell_11959 ( .C (clk), .D (signal_16846), .Q (signal_16847) ) ;
    buf_clk cell_11967 ( .C (clk), .D (signal_16854), .Q (signal_16855) ) ;
    buf_clk cell_11975 ( .C (clk), .D (signal_16862), .Q (signal_16863) ) ;
    buf_clk cell_11983 ( .C (clk), .D (signal_16870), .Q (signal_16871) ) ;
    buf_clk cell_11991 ( .C (clk), .D (signal_16878), .Q (signal_16879) ) ;
    buf_clk cell_11999 ( .C (clk), .D (signal_16886), .Q (signal_16887) ) ;
    buf_clk cell_12007 ( .C (clk), .D (signal_16894), .Q (signal_16895) ) ;
    buf_clk cell_12015 ( .C (clk), .D (signal_16902), .Q (signal_16903) ) ;
    buf_clk cell_12023 ( .C (clk), .D (signal_16910), .Q (signal_16911) ) ;
    buf_clk cell_12031 ( .C (clk), .D (signal_16918), .Q (signal_16919) ) ;
    buf_clk cell_12039 ( .C (clk), .D (signal_16926), .Q (signal_16927) ) ;
    buf_clk cell_12047 ( .C (clk), .D (signal_16934), .Q (signal_16935) ) ;
    buf_clk cell_12055 ( .C (clk), .D (signal_16942), .Q (signal_16943) ) ;
    buf_clk cell_12063 ( .C (clk), .D (signal_16950), .Q (signal_16951) ) ;
    buf_clk cell_12071 ( .C (clk), .D (signal_16958), .Q (signal_16959) ) ;
    buf_clk cell_12079 ( .C (clk), .D (signal_16966), .Q (signal_16967) ) ;
    buf_clk cell_12087 ( .C (clk), .D (signal_16974), .Q (signal_16975) ) ;
    buf_clk cell_12095 ( .C (clk), .D (signal_16982), .Q (signal_16983) ) ;
    buf_clk cell_12103 ( .C (clk), .D (signal_16990), .Q (signal_16991) ) ;
    buf_clk cell_12111 ( .C (clk), .D (signal_16998), .Q (signal_16999) ) ;
    buf_clk cell_12119 ( .C (clk), .D (signal_17006), .Q (signal_17007) ) ;
    buf_clk cell_12127 ( .C (clk), .D (signal_17014), .Q (signal_17015) ) ;
    buf_clk cell_12135 ( .C (clk), .D (signal_17022), .Q (signal_17023) ) ;
    buf_clk cell_12143 ( .C (clk), .D (signal_17030), .Q (signal_17031) ) ;
    buf_clk cell_12151 ( .C (clk), .D (signal_17038), .Q (signal_17039) ) ;
    buf_clk cell_12159 ( .C (clk), .D (signal_17046), .Q (signal_17047) ) ;
    buf_clk cell_12167 ( .C (clk), .D (signal_17054), .Q (signal_17055) ) ;
    buf_clk cell_12175 ( .C (clk), .D (signal_17062), .Q (signal_17063) ) ;
    buf_clk cell_12183 ( .C (clk), .D (signal_17070), .Q (signal_17071) ) ;
    buf_clk cell_12191 ( .C (clk), .D (signal_17078), .Q (signal_17079) ) ;
    buf_clk cell_12199 ( .C (clk), .D (signal_17086), .Q (signal_17087) ) ;
    buf_clk cell_12207 ( .C (clk), .D (signal_17094), .Q (signal_17095) ) ;
    buf_clk cell_12215 ( .C (clk), .D (signal_17102), .Q (signal_17103) ) ;
    buf_clk cell_12223 ( .C (clk), .D (signal_17110), .Q (signal_17111) ) ;
    buf_clk cell_12231 ( .C (clk), .D (signal_17118), .Q (signal_17119) ) ;
    buf_clk cell_12239 ( .C (clk), .D (signal_17126), .Q (signal_17127) ) ;
    buf_clk cell_12247 ( .C (clk), .D (signal_17134), .Q (signal_17135) ) ;
    buf_clk cell_12255 ( .C (clk), .D (signal_17142), .Q (signal_17143) ) ;
    buf_clk cell_12263 ( .C (clk), .D (signal_17150), .Q (signal_17151) ) ;
    buf_clk cell_12271 ( .C (clk), .D (signal_17158), .Q (signal_17159) ) ;
    buf_clk cell_12279 ( .C (clk), .D (signal_17166), .Q (signal_17167) ) ;
    buf_clk cell_12287 ( .C (clk), .D (signal_17174), .Q (signal_17175) ) ;
    buf_clk cell_12295 ( .C (clk), .D (signal_17182), .Q (signal_17183) ) ;
    buf_clk cell_12303 ( .C (clk), .D (signal_17190), .Q (signal_17191) ) ;
    buf_clk cell_12311 ( .C (clk), .D (signal_17198), .Q (signal_17199) ) ;
    buf_clk cell_12319 ( .C (clk), .D (signal_17206), .Q (signal_17207) ) ;
    buf_clk cell_12327 ( .C (clk), .D (signal_17214), .Q (signal_17215) ) ;
    buf_clk cell_12335 ( .C (clk), .D (signal_17222), .Q (signal_17223) ) ;
    buf_clk cell_12343 ( .C (clk), .D (signal_17230), .Q (signal_17231) ) ;
    buf_clk cell_12351 ( .C (clk), .D (signal_17238), .Q (signal_17239) ) ;
    buf_clk cell_12359 ( .C (clk), .D (signal_17246), .Q (signal_17247) ) ;
    buf_clk cell_12367 ( .C (clk), .D (signal_17254), .Q (signal_17255) ) ;
    buf_clk cell_12375 ( .C (clk), .D (signal_17262), .Q (signal_17263) ) ;
    buf_clk cell_12383 ( .C (clk), .D (signal_17270), .Q (signal_17271) ) ;
    buf_clk cell_12391 ( .C (clk), .D (signal_17278), .Q (signal_17279) ) ;
    buf_clk cell_12399 ( .C (clk), .D (signal_17286), .Q (signal_17287) ) ;
    buf_clk cell_12407 ( .C (clk), .D (signal_17294), .Q (signal_17295) ) ;
    buf_clk cell_12415 ( .C (clk), .D (signal_17302), .Q (signal_17303) ) ;
    buf_clk cell_12423 ( .C (clk), .D (signal_17310), .Q (signal_17311) ) ;
    buf_clk cell_12431 ( .C (clk), .D (signal_17318), .Q (signal_17319) ) ;
    buf_clk cell_12439 ( .C (clk), .D (signal_17326), .Q (signal_17327) ) ;
    buf_clk cell_12447 ( .C (clk), .D (signal_17334), .Q (signal_17335) ) ;
    buf_clk cell_12455 ( .C (clk), .D (signal_17342), .Q (signal_17343) ) ;
    buf_clk cell_12463 ( .C (clk), .D (signal_17350), .Q (signal_17351) ) ;
    buf_clk cell_12471 ( .C (clk), .D (signal_17358), .Q (signal_17359) ) ;
    buf_clk cell_12479 ( .C (clk), .D (signal_17366), .Q (signal_17367) ) ;
    buf_clk cell_12487 ( .C (clk), .D (signal_17374), .Q (signal_17375) ) ;
    buf_clk cell_12495 ( .C (clk), .D (signal_17382), .Q (signal_17383) ) ;
    buf_clk cell_12503 ( .C (clk), .D (signal_17390), .Q (signal_17391) ) ;
    buf_clk cell_12511 ( .C (clk), .D (signal_17398), .Q (signal_17399) ) ;
    buf_clk cell_12519 ( .C (clk), .D (signal_17406), .Q (signal_17407) ) ;
    buf_clk cell_12527 ( .C (clk), .D (signal_17414), .Q (signal_17415) ) ;
    buf_clk cell_12535 ( .C (clk), .D (signal_17422), .Q (signal_17423) ) ;
    buf_clk cell_12543 ( .C (clk), .D (signal_17430), .Q (signal_17431) ) ;
    buf_clk cell_12551 ( .C (clk), .D (signal_17438), .Q (signal_17439) ) ;
    buf_clk cell_12559 ( .C (clk), .D (signal_17446), .Q (signal_17447) ) ;
    buf_clk cell_12567 ( .C (clk), .D (signal_17454), .Q (signal_17455) ) ;
    buf_clk cell_12575 ( .C (clk), .D (signal_17462), .Q (signal_17463) ) ;
    buf_clk cell_12583 ( .C (clk), .D (signal_17470), .Q (signal_17471) ) ;
    buf_clk cell_12591 ( .C (clk), .D (signal_17478), .Q (signal_17479) ) ;
    buf_clk cell_12599 ( .C (clk), .D (signal_17486), .Q (signal_17487) ) ;
    buf_clk cell_12607 ( .C (clk), .D (signal_17494), .Q (signal_17495) ) ;
    buf_clk cell_12615 ( .C (clk), .D (signal_17502), .Q (signal_17503) ) ;
    buf_clk cell_12623 ( .C (clk), .D (signal_17510), .Q (signal_17511) ) ;
    buf_clk cell_12631 ( .C (clk), .D (signal_17518), .Q (signal_17519) ) ;
    buf_clk cell_12639 ( .C (clk), .D (signal_17526), .Q (signal_17527) ) ;
    buf_clk cell_12647 ( .C (clk), .D (signal_17534), .Q (signal_17535) ) ;
    buf_clk cell_12655 ( .C (clk), .D (signal_17542), .Q (signal_17543) ) ;
    buf_clk cell_12663 ( .C (clk), .D (signal_17550), .Q (signal_17551) ) ;
    buf_clk cell_12671 ( .C (clk), .D (signal_17558), .Q (signal_17559) ) ;
    buf_clk cell_12679 ( .C (clk), .D (signal_17566), .Q (signal_17567) ) ;
    buf_clk cell_12687 ( .C (clk), .D (signal_17574), .Q (signal_17575) ) ;
    buf_clk cell_12695 ( .C (clk), .D (signal_17582), .Q (signal_17583) ) ;
    buf_clk cell_12703 ( .C (clk), .D (signal_17590), .Q (signal_17591) ) ;
    buf_clk cell_12711 ( .C (clk), .D (signal_17598), .Q (signal_17599) ) ;
    buf_clk cell_12719 ( .C (clk), .D (signal_17606), .Q (signal_17607) ) ;
    buf_clk cell_12727 ( .C (clk), .D (signal_17614), .Q (signal_17615) ) ;
    buf_clk cell_12735 ( .C (clk), .D (signal_17622), .Q (signal_17623) ) ;
    buf_clk cell_12743 ( .C (clk), .D (signal_17630), .Q (signal_17631) ) ;
    buf_clk cell_12751 ( .C (clk), .D (signal_17638), .Q (signal_17639) ) ;
    buf_clk cell_12759 ( .C (clk), .D (signal_17646), .Q (signal_17647) ) ;
    buf_clk cell_12767 ( .C (clk), .D (signal_17654), .Q (signal_17655) ) ;
    buf_clk cell_12775 ( .C (clk), .D (signal_17662), .Q (signal_17663) ) ;
    buf_clk cell_12783 ( .C (clk), .D (signal_17670), .Q (signal_17671) ) ;
    buf_clk cell_12791 ( .C (clk), .D (signal_17678), .Q (signal_17679) ) ;
    buf_clk cell_12799 ( .C (clk), .D (signal_17686), .Q (signal_17687) ) ;
    buf_clk cell_12807 ( .C (clk), .D (signal_17694), .Q (signal_17695) ) ;
    buf_clk cell_12815 ( .C (clk), .D (signal_17702), .Q (signal_17703) ) ;
    buf_clk cell_12823 ( .C (clk), .D (signal_17710), .Q (signal_17711) ) ;
    buf_clk cell_12831 ( .C (clk), .D (signal_17718), .Q (signal_17719) ) ;
    buf_clk cell_12839 ( .C (clk), .D (signal_17726), .Q (signal_17727) ) ;
    buf_clk cell_12847 ( .C (clk), .D (signal_17734), .Q (signal_17735) ) ;
    buf_clk cell_12855 ( .C (clk), .D (signal_17742), .Q (signal_17743) ) ;
    buf_clk cell_12863 ( .C (clk), .D (signal_17750), .Q (signal_17751) ) ;
    buf_clk cell_12871 ( .C (clk), .D (signal_17758), .Q (signal_17759) ) ;
    buf_clk cell_12879 ( .C (clk), .D (signal_17766), .Q (signal_17767) ) ;
    buf_clk cell_12887 ( .C (clk), .D (signal_17774), .Q (signal_17775) ) ;
    buf_clk cell_12895 ( .C (clk), .D (signal_17782), .Q (signal_17783) ) ;
    buf_clk cell_12903 ( .C (clk), .D (signal_17790), .Q (signal_17791) ) ;
    buf_clk cell_12911 ( .C (clk), .D (signal_17798), .Q (signal_17799) ) ;
    buf_clk cell_12919 ( .C (clk), .D (signal_17806), .Q (signal_17807) ) ;
    buf_clk cell_12927 ( .C (clk), .D (signal_17814), .Q (signal_17815) ) ;
    buf_clk cell_12935 ( .C (clk), .D (signal_17822), .Q (signal_17823) ) ;
    buf_clk cell_12943 ( .C (clk), .D (signal_17830), .Q (signal_17831) ) ;
    buf_clk cell_12951 ( .C (clk), .D (signal_17838), .Q (signal_17839) ) ;
    buf_clk cell_12959 ( .C (clk), .D (signal_17846), .Q (signal_17847) ) ;
    buf_clk cell_12967 ( .C (clk), .D (signal_17854), .Q (signal_17855) ) ;
    buf_clk cell_12975 ( .C (clk), .D (signal_17862), .Q (signal_17863) ) ;
    buf_clk cell_12983 ( .C (clk), .D (signal_17870), .Q (signal_17871) ) ;
    buf_clk cell_12991 ( .C (clk), .D (signal_17878), .Q (signal_17879) ) ;
    buf_clk cell_12999 ( .C (clk), .D (signal_17886), .Q (signal_17887) ) ;
    buf_clk cell_13007 ( .C (clk), .D (signal_17894), .Q (signal_17895) ) ;
    buf_clk cell_13015 ( .C (clk), .D (signal_17902), .Q (signal_17903) ) ;
    buf_clk cell_13023 ( .C (clk), .D (signal_17910), .Q (signal_17911) ) ;
    buf_clk cell_13031 ( .C (clk), .D (signal_17918), .Q (signal_17919) ) ;
    buf_clk cell_13039 ( .C (clk), .D (signal_17926), .Q (signal_17927) ) ;
    buf_clk cell_13047 ( .C (clk), .D (signal_17934), .Q (signal_17935) ) ;
    buf_clk cell_13055 ( .C (clk), .D (signal_17942), .Q (signal_17943) ) ;
    buf_clk cell_13063 ( .C (clk), .D (signal_17950), .Q (signal_17951) ) ;
    buf_clk cell_13071 ( .C (clk), .D (signal_17958), .Q (signal_17959) ) ;
    buf_clk cell_13079 ( .C (clk), .D (signal_17966), .Q (signal_17967) ) ;
    buf_clk cell_13087 ( .C (clk), .D (signal_17974), .Q (signal_17975) ) ;
    buf_clk cell_13095 ( .C (clk), .D (signal_17982), .Q (signal_17983) ) ;
    buf_clk cell_13103 ( .C (clk), .D (signal_17990), .Q (signal_17991) ) ;
    buf_clk cell_13111 ( .C (clk), .D (signal_17998), .Q (signal_17999) ) ;
    buf_clk cell_13119 ( .C (clk), .D (signal_18006), .Q (signal_18007) ) ;
    buf_clk cell_13127 ( .C (clk), .D (signal_18014), .Q (signal_18015) ) ;
    buf_clk cell_13135 ( .C (clk), .D (signal_18022), .Q (signal_18023) ) ;
    buf_clk cell_13143 ( .C (clk), .D (signal_18030), .Q (signal_18031) ) ;
    buf_clk cell_13151 ( .C (clk), .D (signal_18038), .Q (signal_18039) ) ;
    buf_clk cell_13159 ( .C (clk), .D (signal_18046), .Q (signal_18047) ) ;
    buf_clk cell_13167 ( .C (clk), .D (signal_18054), .Q (signal_18055) ) ;
    buf_clk cell_13175 ( .C (clk), .D (signal_18062), .Q (signal_18063) ) ;
    buf_clk cell_13183 ( .C (clk), .D (signal_18070), .Q (signal_18071) ) ;
    buf_clk cell_13191 ( .C (clk), .D (signal_18078), .Q (signal_18079) ) ;
    buf_clk cell_13199 ( .C (clk), .D (signal_18086), .Q (signal_18087) ) ;
    buf_clk cell_13207 ( .C (clk), .D (signal_18094), .Q (signal_18095) ) ;
    buf_clk cell_13215 ( .C (clk), .D (signal_18102), .Q (signal_18103) ) ;
    buf_clk cell_13223 ( .C (clk), .D (signal_18110), .Q (signal_18111) ) ;
    buf_clk cell_13231 ( .C (clk), .D (signal_18118), .Q (signal_18119) ) ;
    buf_clk cell_13239 ( .C (clk), .D (signal_18126), .Q (signal_18127) ) ;
    buf_clk cell_13247 ( .C (clk), .D (signal_18134), .Q (signal_18135) ) ;
    buf_clk cell_13255 ( .C (clk), .D (signal_18142), .Q (signal_18143) ) ;
    buf_clk cell_13263 ( .C (clk), .D (signal_18150), .Q (signal_18151) ) ;
    buf_clk cell_13271 ( .C (clk), .D (signal_18158), .Q (signal_18159) ) ;
    buf_clk cell_13279 ( .C (clk), .D (signal_18166), .Q (signal_18167) ) ;
    buf_clk cell_13285 ( .C (clk), .D (signal_18172), .Q (signal_18173) ) ;
    buf_clk cell_13291 ( .C (clk), .D (signal_18178), .Q (signal_18179) ) ;
    buf_clk cell_13297 ( .C (clk), .D (signal_18184), .Q (signal_18185) ) ;
    buf_clk cell_13303 ( .C (clk), .D (signal_18190), .Q (signal_18191) ) ;
    buf_clk cell_13309 ( .C (clk), .D (signal_18196), .Q (signal_18197) ) ;
    buf_clk cell_13315 ( .C (clk), .D (signal_18202), .Q (signal_18203) ) ;
    buf_clk cell_13321 ( .C (clk), .D (signal_18208), .Q (signal_18209) ) ;
    buf_clk cell_13327 ( .C (clk), .D (signal_18214), .Q (signal_18215) ) ;
    buf_clk cell_13333 ( .C (clk), .D (signal_18220), .Q (signal_18221) ) ;
    buf_clk cell_13339 ( .C (clk), .D (signal_18226), .Q (signal_18227) ) ;
    buf_clk cell_13345 ( .C (clk), .D (signal_18232), .Q (signal_18233) ) ;
    buf_clk cell_13351 ( .C (clk), .D (signal_18238), .Q (signal_18239) ) ;
    buf_clk cell_13357 ( .C (clk), .D (signal_18244), .Q (signal_18245) ) ;
    buf_clk cell_13363 ( .C (clk), .D (signal_18250), .Q (signal_18251) ) ;
    buf_clk cell_13369 ( .C (clk), .D (signal_18256), .Q (signal_18257) ) ;
    buf_clk cell_13375 ( .C (clk), .D (signal_18262), .Q (signal_18263) ) ;
    buf_clk cell_13381 ( .C (clk), .D (signal_18268), .Q (signal_18269) ) ;
    buf_clk cell_13387 ( .C (clk), .D (signal_18274), .Q (signal_18275) ) ;
    buf_clk cell_13393 ( .C (clk), .D (signal_18280), .Q (signal_18281) ) ;
    buf_clk cell_13399 ( .C (clk), .D (signal_18286), .Q (signal_18287) ) ;
    buf_clk cell_13405 ( .C (clk), .D (signal_18292), .Q (signal_18293) ) ;
    buf_clk cell_13411 ( .C (clk), .D (signal_18298), .Q (signal_18299) ) ;
    buf_clk cell_13417 ( .C (clk), .D (signal_18304), .Q (signal_18305) ) ;
    buf_clk cell_13423 ( .C (clk), .D (signal_18310), .Q (signal_18311) ) ;
    buf_clk cell_13429 ( .C (clk), .D (signal_18316), .Q (signal_18317) ) ;
    buf_clk cell_13435 ( .C (clk), .D (signal_18322), .Q (signal_18323) ) ;
    buf_clk cell_13441 ( .C (clk), .D (signal_18328), .Q (signal_18329) ) ;
    buf_clk cell_13447 ( .C (clk), .D (signal_18334), .Q (signal_18335) ) ;
    buf_clk cell_13453 ( .C (clk), .D (signal_18340), .Q (signal_18341) ) ;
    buf_clk cell_13459 ( .C (clk), .D (signal_18346), .Q (signal_18347) ) ;
    buf_clk cell_13465 ( .C (clk), .D (signal_18352), .Q (signal_18353) ) ;
    buf_clk cell_13471 ( .C (clk), .D (signal_18358), .Q (signal_18359) ) ;
    buf_clk cell_13477 ( .C (clk), .D (signal_18364), .Q (signal_18365) ) ;
    buf_clk cell_13483 ( .C (clk), .D (signal_18370), .Q (signal_18371) ) ;
    buf_clk cell_13489 ( .C (clk), .D (signal_18376), .Q (signal_18377) ) ;
    buf_clk cell_13495 ( .C (clk), .D (signal_18382), .Q (signal_18383) ) ;
    buf_clk cell_13501 ( .C (clk), .D (signal_18388), .Q (signal_18389) ) ;
    buf_clk cell_13507 ( .C (clk), .D (signal_18394), .Q (signal_18395) ) ;
    buf_clk cell_13513 ( .C (clk), .D (signal_18400), .Q (signal_18401) ) ;
    buf_clk cell_13519 ( .C (clk), .D (signal_18406), .Q (signal_18407) ) ;
    buf_clk cell_13525 ( .C (clk), .D (signal_18412), .Q (signal_18413) ) ;
    buf_clk cell_13531 ( .C (clk), .D (signal_18418), .Q (signal_18419) ) ;
    buf_clk cell_13537 ( .C (clk), .D (signal_18424), .Q (signal_18425) ) ;
    buf_clk cell_13543 ( .C (clk), .D (signal_18430), .Q (signal_18431) ) ;
    buf_clk cell_13549 ( .C (clk), .D (signal_18436), .Q (signal_18437) ) ;
    buf_clk cell_13555 ( .C (clk), .D (signal_18442), .Q (signal_18443) ) ;
    buf_clk cell_13561 ( .C (clk), .D (signal_18448), .Q (signal_18449) ) ;
    buf_clk cell_13567 ( .C (clk), .D (signal_18454), .Q (signal_18455) ) ;
    buf_clk cell_13573 ( .C (clk), .D (signal_18460), .Q (signal_18461) ) ;
    buf_clk cell_13579 ( .C (clk), .D (signal_18466), .Q (signal_18467) ) ;
    buf_clk cell_13585 ( .C (clk), .D (signal_18472), .Q (signal_18473) ) ;
    buf_clk cell_13591 ( .C (clk), .D (signal_18478), .Q (signal_18479) ) ;
    buf_clk cell_13597 ( .C (clk), .D (signal_18484), .Q (signal_18485) ) ;
    buf_clk cell_13603 ( .C (clk), .D (signal_18490), .Q (signal_18491) ) ;
    buf_clk cell_13609 ( .C (clk), .D (signal_18496), .Q (signal_18497) ) ;
    buf_clk cell_13615 ( .C (clk), .D (signal_18502), .Q (signal_18503) ) ;
    buf_clk cell_13621 ( .C (clk), .D (signal_18508), .Q (signal_18509) ) ;
    buf_clk cell_13627 ( .C (clk), .D (signal_18514), .Q (signal_18515) ) ;
    buf_clk cell_13633 ( .C (clk), .D (signal_18520), .Q (signal_18521) ) ;
    buf_clk cell_13639 ( .C (clk), .D (signal_18526), .Q (signal_18527) ) ;
    buf_clk cell_13645 ( .C (clk), .D (signal_18532), .Q (signal_18533) ) ;
    buf_clk cell_13651 ( .C (clk), .D (signal_18538), .Q (signal_18539) ) ;
    buf_clk cell_13657 ( .C (clk), .D (signal_18544), .Q (signal_18545) ) ;
    buf_clk cell_13663 ( .C (clk), .D (signal_18550), .Q (signal_18551) ) ;
    buf_clk cell_13669 ( .C (clk), .D (signal_18556), .Q (signal_18557) ) ;
    buf_clk cell_13675 ( .C (clk), .D (signal_18562), .Q (signal_18563) ) ;
    buf_clk cell_13681 ( .C (clk), .D (signal_18568), .Q (signal_18569) ) ;
    buf_clk cell_13687 ( .C (clk), .D (signal_18574), .Q (signal_18575) ) ;
    buf_clk cell_13693 ( .C (clk), .D (signal_18580), .Q (signal_18581) ) ;
    buf_clk cell_13699 ( .C (clk), .D (signal_18586), .Q (signal_18587) ) ;
    buf_clk cell_13705 ( .C (clk), .D (signal_18592), .Q (signal_18593) ) ;
    buf_clk cell_13711 ( .C (clk), .D (signal_18598), .Q (signal_18599) ) ;
    buf_clk cell_13717 ( .C (clk), .D (signal_18604), .Q (signal_18605) ) ;
    buf_clk cell_13723 ( .C (clk), .D (signal_18610), .Q (signal_18611) ) ;
    buf_clk cell_13729 ( .C (clk), .D (signal_18616), .Q (signal_18617) ) ;
    buf_clk cell_13735 ( .C (clk), .D (signal_18622), .Q (signal_18623) ) ;
    buf_clk cell_13741 ( .C (clk), .D (signal_18628), .Q (signal_18629) ) ;
    buf_clk cell_13747 ( .C (clk), .D (signal_18634), .Q (signal_18635) ) ;
    buf_clk cell_13753 ( .C (clk), .D (signal_18640), .Q (signal_18641) ) ;
    buf_clk cell_13759 ( .C (clk), .D (signal_18646), .Q (signal_18647) ) ;
    buf_clk cell_13765 ( .C (clk), .D (signal_18652), .Q (signal_18653) ) ;
    buf_clk cell_13771 ( .C (clk), .D (signal_18658), .Q (signal_18659) ) ;
    buf_clk cell_13777 ( .C (clk), .D (signal_18664), .Q (signal_18665) ) ;
    buf_clk cell_13783 ( .C (clk), .D (signal_18670), .Q (signal_18671) ) ;
    buf_clk cell_13789 ( .C (clk), .D (signal_18676), .Q (signal_18677) ) ;
    buf_clk cell_13795 ( .C (clk), .D (signal_18682), .Q (signal_18683) ) ;
    buf_clk cell_13801 ( .C (clk), .D (signal_18688), .Q (signal_18689) ) ;
    buf_clk cell_13807 ( .C (clk), .D (signal_18694), .Q (signal_18695) ) ;
    buf_clk cell_13813 ( .C (clk), .D (signal_18700), .Q (signal_18701) ) ;
    buf_clk cell_13819 ( .C (clk), .D (signal_18706), .Q (signal_18707) ) ;
    buf_clk cell_13825 ( .C (clk), .D (signal_18712), .Q (signal_18713) ) ;
    buf_clk cell_13831 ( .C (clk), .D (signal_18718), .Q (signal_18719) ) ;
    buf_clk cell_13837 ( .C (clk), .D (signal_18724), .Q (signal_18725) ) ;
    buf_clk cell_13843 ( .C (clk), .D (signal_18730), .Q (signal_18731) ) ;
    buf_clk cell_13849 ( .C (clk), .D (signal_18736), .Q (signal_18737) ) ;
    buf_clk cell_13855 ( .C (clk), .D (signal_18742), .Q (signal_18743) ) ;
    buf_clk cell_13861 ( .C (clk), .D (signal_18748), .Q (signal_18749) ) ;
    buf_clk cell_13867 ( .C (clk), .D (signal_18754), .Q (signal_18755) ) ;
    buf_clk cell_13873 ( .C (clk), .D (signal_18760), .Q (signal_18761) ) ;
    buf_clk cell_13879 ( .C (clk), .D (signal_18766), .Q (signal_18767) ) ;
    buf_clk cell_13885 ( .C (clk), .D (signal_18772), .Q (signal_18773) ) ;
    buf_clk cell_13891 ( .C (clk), .D (signal_18778), .Q (signal_18779) ) ;
    buf_clk cell_13897 ( .C (clk), .D (signal_18784), .Q (signal_18785) ) ;
    buf_clk cell_13903 ( .C (clk), .D (signal_18790), .Q (signal_18791) ) ;
    buf_clk cell_13909 ( .C (clk), .D (signal_18796), .Q (signal_18797) ) ;
    buf_clk cell_13915 ( .C (clk), .D (signal_18802), .Q (signal_18803) ) ;
    buf_clk cell_13921 ( .C (clk), .D (signal_18808), .Q (signal_18809) ) ;
    buf_clk cell_13927 ( .C (clk), .D (signal_18814), .Q (signal_18815) ) ;
    buf_clk cell_13933 ( .C (clk), .D (signal_18820), .Q (signal_18821) ) ;
    buf_clk cell_13939 ( .C (clk), .D (signal_18826), .Q (signal_18827) ) ;
    buf_clk cell_13945 ( .C (clk), .D (signal_18832), .Q (signal_18833) ) ;
    buf_clk cell_13951 ( .C (clk), .D (signal_18838), .Q (signal_18839) ) ;
    buf_clk cell_13957 ( .C (clk), .D (signal_18844), .Q (signal_18845) ) ;
    buf_clk cell_13963 ( .C (clk), .D (signal_18850), .Q (signal_18851) ) ;
    buf_clk cell_13969 ( .C (clk), .D (signal_18856), .Q (signal_18857) ) ;
    buf_clk cell_13975 ( .C (clk), .D (signal_18862), .Q (signal_18863) ) ;
    buf_clk cell_13981 ( .C (clk), .D (signal_18868), .Q (signal_18869) ) ;
    buf_clk cell_13987 ( .C (clk), .D (signal_18874), .Q (signal_18875) ) ;
    buf_clk cell_13993 ( .C (clk), .D (signal_18880), .Q (signal_18881) ) ;
    buf_clk cell_13999 ( .C (clk), .D (signal_18886), .Q (signal_18887) ) ;
    buf_clk cell_14005 ( .C (clk), .D (signal_18892), .Q (signal_18893) ) ;
    buf_clk cell_14011 ( .C (clk), .D (signal_18898), .Q (signal_18899) ) ;
    buf_clk cell_14017 ( .C (clk), .D (signal_18904), .Q (signal_18905) ) ;
    buf_clk cell_14023 ( .C (clk), .D (signal_18910), .Q (signal_18911) ) ;
    buf_clk cell_14029 ( .C (clk), .D (signal_18916), .Q (signal_18917) ) ;
    buf_clk cell_14035 ( .C (clk), .D (signal_18922), .Q (signal_18923) ) ;
    buf_clk cell_14041 ( .C (clk), .D (signal_18928), .Q (signal_18929) ) ;
    buf_clk cell_14047 ( .C (clk), .D (signal_18934), .Q (signal_18935) ) ;
    buf_clk cell_14053 ( .C (clk), .D (signal_18940), .Q (signal_18941) ) ;
    buf_clk cell_14059 ( .C (clk), .D (signal_18946), .Q (signal_18947) ) ;
    buf_clk cell_14065 ( .C (clk), .D (signal_18952), .Q (signal_18953) ) ;
    buf_clk cell_14071 ( .C (clk), .D (signal_18958), .Q (signal_18959) ) ;
    buf_clk cell_14077 ( .C (clk), .D (signal_18964), .Q (signal_18965) ) ;
    buf_clk cell_14083 ( .C (clk), .D (signal_18970), .Q (signal_18971) ) ;
    buf_clk cell_14089 ( .C (clk), .D (signal_18976), .Q (signal_18977) ) ;
    buf_clk cell_14095 ( .C (clk), .D (signal_18982), .Q (signal_18983) ) ;
    buf_clk cell_14101 ( .C (clk), .D (signal_18988), .Q (signal_18989) ) ;
    buf_clk cell_14107 ( .C (clk), .D (signal_18994), .Q (signal_18995) ) ;
    buf_clk cell_14113 ( .C (clk), .D (signal_19000), .Q (signal_19001) ) ;
    buf_clk cell_14119 ( .C (clk), .D (signal_19006), .Q (signal_19007) ) ;
    buf_clk cell_14125 ( .C (clk), .D (signal_19012), .Q (signal_19013) ) ;
    buf_clk cell_14131 ( .C (clk), .D (signal_19018), .Q (signal_19019) ) ;
    buf_clk cell_14137 ( .C (clk), .D (signal_19024), .Q (signal_19025) ) ;
    buf_clk cell_14143 ( .C (clk), .D (signal_19030), .Q (signal_19031) ) ;
    buf_clk cell_14149 ( .C (clk), .D (signal_19036), .Q (signal_19037) ) ;
    buf_clk cell_14155 ( .C (clk), .D (signal_19042), .Q (signal_19043) ) ;
    buf_clk cell_14161 ( .C (clk), .D (signal_19048), .Q (signal_19049) ) ;
    buf_clk cell_14167 ( .C (clk), .D (signal_19054), .Q (signal_19055) ) ;
    buf_clk cell_14173 ( .C (clk), .D (signal_19060), .Q (signal_19061) ) ;
    buf_clk cell_14179 ( .C (clk), .D (signal_19066), .Q (signal_19067) ) ;
    buf_clk cell_14185 ( .C (clk), .D (signal_19072), .Q (signal_19073) ) ;
    buf_clk cell_14191 ( .C (clk), .D (signal_19078), .Q (signal_19079) ) ;
    buf_clk cell_14197 ( .C (clk), .D (signal_19084), .Q (signal_19085) ) ;
    buf_clk cell_14203 ( .C (clk), .D (signal_19090), .Q (signal_19091) ) ;
    buf_clk cell_14209 ( .C (clk), .D (signal_19096), .Q (signal_19097) ) ;
    buf_clk cell_14215 ( .C (clk), .D (signal_19102), .Q (signal_19103) ) ;
    buf_clk cell_14221 ( .C (clk), .D (signal_19108), .Q (signal_19109) ) ;
    buf_clk cell_14227 ( .C (clk), .D (signal_19114), .Q (signal_19115) ) ;
    buf_clk cell_14233 ( .C (clk), .D (signal_19120), .Q (signal_19121) ) ;
    buf_clk cell_14239 ( .C (clk), .D (signal_19126), .Q (signal_19127) ) ;
    buf_clk cell_14245 ( .C (clk), .D (signal_19132), .Q (signal_19133) ) ;
    buf_clk cell_14251 ( .C (clk), .D (signal_19138), .Q (signal_19139) ) ;
    buf_clk cell_14257 ( .C (clk), .D (signal_19144), .Q (signal_19145) ) ;
    buf_clk cell_14263 ( .C (clk), .D (signal_19150), .Q (signal_19151) ) ;
    buf_clk cell_14269 ( .C (clk), .D (signal_19156), .Q (signal_19157) ) ;
    buf_clk cell_14275 ( .C (clk), .D (signal_19162), .Q (signal_19163) ) ;
    buf_clk cell_14281 ( .C (clk), .D (signal_19168), .Q (signal_19169) ) ;
    buf_clk cell_14287 ( .C (clk), .D (signal_19174), .Q (signal_19175) ) ;
    buf_clk cell_14293 ( .C (clk), .D (signal_19180), .Q (signal_19181) ) ;
    buf_clk cell_14299 ( .C (clk), .D (signal_19186), .Q (signal_19187) ) ;
    buf_clk cell_14305 ( .C (clk), .D (signal_19192), .Q (signal_19193) ) ;
    buf_clk cell_14311 ( .C (clk), .D (signal_19198), .Q (signal_19199) ) ;
    buf_clk cell_14317 ( .C (clk), .D (signal_19204), .Q (signal_19205) ) ;
    buf_clk cell_14323 ( .C (clk), .D (signal_19210), .Q (signal_19211) ) ;
    buf_clk cell_14329 ( .C (clk), .D (signal_19216), .Q (signal_19217) ) ;
    buf_clk cell_14335 ( .C (clk), .D (signal_19222), .Q (signal_19223) ) ;
    buf_clk cell_14341 ( .C (clk), .D (signal_19228), .Q (signal_19229) ) ;
    buf_clk cell_14347 ( .C (clk), .D (signal_19234), .Q (signal_19235) ) ;
    buf_clk cell_14353 ( .C (clk), .D (signal_19240), .Q (signal_19241) ) ;
    buf_clk cell_14359 ( .C (clk), .D (signal_19246), .Q (signal_19247) ) ;
    buf_clk cell_14365 ( .C (clk), .D (signal_19252), .Q (signal_19253) ) ;
    buf_clk cell_14371 ( .C (clk), .D (signal_19258), .Q (signal_19259) ) ;
    buf_clk cell_14377 ( .C (clk), .D (signal_19264), .Q (signal_19265) ) ;
    buf_clk cell_14383 ( .C (clk), .D (signal_19270), .Q (signal_19271) ) ;
    buf_clk cell_14389 ( .C (clk), .D (signal_19276), .Q (signal_19277) ) ;
    buf_clk cell_14395 ( .C (clk), .D (signal_19282), .Q (signal_19283) ) ;
    buf_clk cell_14401 ( .C (clk), .D (signal_19288), .Q (signal_19289) ) ;
    buf_clk cell_14407 ( .C (clk), .D (signal_19294), .Q (signal_19295) ) ;
    buf_clk cell_14413 ( .C (clk), .D (signal_19300), .Q (signal_19301) ) ;
    buf_clk cell_14419 ( .C (clk), .D (signal_19306), .Q (signal_19307) ) ;
    buf_clk cell_14425 ( .C (clk), .D (signal_19312), .Q (signal_19313) ) ;
    buf_clk cell_14431 ( .C (clk), .D (signal_19318), .Q (signal_19319) ) ;
    buf_clk cell_14437 ( .C (clk), .D (signal_19324), .Q (signal_19325) ) ;
    buf_clk cell_14443 ( .C (clk), .D (signal_19330), .Q (signal_19331) ) ;
    buf_clk cell_14449 ( .C (clk), .D (signal_19336), .Q (signal_19337) ) ;
    buf_clk cell_14455 ( .C (clk), .D (signal_19342), .Q (signal_19343) ) ;
    buf_clk cell_14461 ( .C (clk), .D (signal_19348), .Q (signal_19349) ) ;
    buf_clk cell_14467 ( .C (clk), .D (signal_19354), .Q (signal_19355) ) ;
    buf_clk cell_14473 ( .C (clk), .D (signal_19360), .Q (signal_19361) ) ;
    buf_clk cell_14479 ( .C (clk), .D (signal_19366), .Q (signal_19367) ) ;
    buf_clk cell_14485 ( .C (clk), .D (signal_19372), .Q (signal_19373) ) ;
    buf_clk cell_14491 ( .C (clk), .D (signal_19378), .Q (signal_19379) ) ;
    buf_clk cell_14497 ( .C (clk), .D (signal_19384), .Q (signal_19385) ) ;
    buf_clk cell_14503 ( .C (clk), .D (signal_19390), .Q (signal_19391) ) ;
    buf_clk cell_14509 ( .C (clk), .D (signal_19396), .Q (signal_19397) ) ;
    buf_clk cell_14515 ( .C (clk), .D (signal_19402), .Q (signal_19403) ) ;
    buf_clk cell_14521 ( .C (clk), .D (signal_19408), .Q (signal_19409) ) ;
    buf_clk cell_14527 ( .C (clk), .D (signal_19414), .Q (signal_19415) ) ;
    buf_clk cell_14533 ( .C (clk), .D (signal_19420), .Q (signal_19421) ) ;
    buf_clk cell_14539 ( .C (clk), .D (signal_19426), .Q (signal_19427) ) ;
    buf_clk cell_14545 ( .C (clk), .D (signal_19432), .Q (signal_19433) ) ;
    buf_clk cell_14551 ( .C (clk), .D (signal_19438), .Q (signal_19439) ) ;
    buf_clk cell_14557 ( .C (clk), .D (signal_19444), .Q (signal_19445) ) ;
    buf_clk cell_14563 ( .C (clk), .D (signal_19450), .Q (signal_19451) ) ;
    buf_clk cell_14569 ( .C (clk), .D (signal_19456), .Q (signal_19457) ) ;
    buf_clk cell_14575 ( .C (clk), .D (signal_19462), .Q (signal_19463) ) ;
    buf_clk cell_14581 ( .C (clk), .D (signal_19468), .Q (signal_19469) ) ;
    buf_clk cell_14587 ( .C (clk), .D (signal_19474), .Q (signal_19475) ) ;
    buf_clk cell_14593 ( .C (clk), .D (signal_19480), .Q (signal_19481) ) ;
    buf_clk cell_14599 ( .C (clk), .D (signal_19486), .Q (signal_19487) ) ;
    buf_clk cell_14605 ( .C (clk), .D (signal_19492), .Q (signal_19493) ) ;
    buf_clk cell_14611 ( .C (clk), .D (signal_19498), .Q (signal_19499) ) ;
    buf_clk cell_14617 ( .C (clk), .D (signal_19504), .Q (signal_19505) ) ;
    buf_clk cell_14623 ( .C (clk), .D (signal_19510), .Q (signal_19511) ) ;
    buf_clk cell_14629 ( .C (clk), .D (signal_19516), .Q (signal_19517) ) ;
    buf_clk cell_14635 ( .C (clk), .D (signal_19522), .Q (signal_19523) ) ;
    buf_clk cell_14641 ( .C (clk), .D (signal_19528), .Q (signal_19529) ) ;
    buf_clk cell_14647 ( .C (clk), .D (signal_19534), .Q (signal_19535) ) ;
    buf_clk cell_14653 ( .C (clk), .D (signal_19540), .Q (signal_19541) ) ;
    buf_clk cell_14659 ( .C (clk), .D (signal_19546), .Q (signal_19547) ) ;
    buf_clk cell_14665 ( .C (clk), .D (signal_19552), .Q (signal_19553) ) ;
    buf_clk cell_14671 ( .C (clk), .D (signal_19558), .Q (signal_19559) ) ;
    buf_clk cell_14677 ( .C (clk), .D (signal_19564), .Q (signal_19565) ) ;
    buf_clk cell_14683 ( .C (clk), .D (signal_19570), .Q (signal_19571) ) ;
    buf_clk cell_14689 ( .C (clk), .D (signal_19576), .Q (signal_19577) ) ;
    buf_clk cell_14695 ( .C (clk), .D (signal_19582), .Q (signal_19583) ) ;
    buf_clk cell_14701 ( .C (clk), .D (signal_19588), .Q (signal_19589) ) ;
    buf_clk cell_14707 ( .C (clk), .D (signal_19594), .Q (signal_19595) ) ;
    buf_clk cell_14713 ( .C (clk), .D (signal_19600), .Q (signal_19601) ) ;
    buf_clk cell_14719 ( .C (clk), .D (signal_19606), .Q (signal_19607) ) ;
    buf_clk cell_14725 ( .C (clk), .D (signal_19612), .Q (signal_19613) ) ;
    buf_clk cell_14731 ( .C (clk), .D (signal_19618), .Q (signal_19619) ) ;
    buf_clk cell_14737 ( .C (clk), .D (signal_19624), .Q (signal_19625) ) ;
    buf_clk cell_14743 ( .C (clk), .D (signal_19630), .Q (signal_19631) ) ;
    buf_clk cell_14749 ( .C (clk), .D (signal_19636), .Q (signal_19637) ) ;
    buf_clk cell_14755 ( .C (clk), .D (signal_19642), .Q (signal_19643) ) ;
    buf_clk cell_14761 ( .C (clk), .D (signal_19648), .Q (signal_19649) ) ;
    buf_clk cell_14767 ( .C (clk), .D (signal_19654), .Q (signal_19655) ) ;
    buf_clk cell_14773 ( .C (clk), .D (signal_19660), .Q (signal_19661) ) ;
    buf_clk cell_14779 ( .C (clk), .D (signal_19666), .Q (signal_19667) ) ;
    buf_clk cell_14785 ( .C (clk), .D (signal_19672), .Q (signal_19673) ) ;
    buf_clk cell_14791 ( .C (clk), .D (signal_19678), .Q (signal_19679) ) ;
    buf_clk cell_14797 ( .C (clk), .D (signal_19684), .Q (signal_19685) ) ;
    buf_clk cell_14803 ( .C (clk), .D (signal_19690), .Q (signal_19691) ) ;
    buf_clk cell_14809 ( .C (clk), .D (signal_19696), .Q (signal_19697) ) ;
    buf_clk cell_14815 ( .C (clk), .D (signal_19702), .Q (signal_19703) ) ;
    buf_clk cell_14821 ( .C (clk), .D (signal_19708), .Q (signal_19709) ) ;
    buf_clk cell_14827 ( .C (clk), .D (signal_19714), .Q (signal_19715) ) ;
    buf_clk cell_14833 ( .C (clk), .D (signal_19720), .Q (signal_19721) ) ;
    buf_clk cell_14839 ( .C (clk), .D (signal_19726), .Q (signal_19727) ) ;
    buf_clk cell_14845 ( .C (clk), .D (signal_19732), .Q (signal_19733) ) ;
    buf_clk cell_14851 ( .C (clk), .D (signal_19738), .Q (signal_19739) ) ;
    buf_clk cell_14857 ( .C (clk), .D (signal_19744), .Q (signal_19745) ) ;
    buf_clk cell_14863 ( .C (clk), .D (signal_19750), .Q (signal_19751) ) ;
    buf_clk cell_14869 ( .C (clk), .D (signal_19756), .Q (signal_19757) ) ;
    buf_clk cell_14875 ( .C (clk), .D (signal_19762), .Q (signal_19763) ) ;
    buf_clk cell_14881 ( .C (clk), .D (signal_19768), .Q (signal_19769) ) ;
    buf_clk cell_14887 ( .C (clk), .D (signal_19774), .Q (signal_19775) ) ;
    buf_clk cell_14893 ( .C (clk), .D (signal_19780), .Q (signal_19781) ) ;
    buf_clk cell_14899 ( .C (clk), .D (signal_19786), .Q (signal_19787) ) ;
    buf_clk cell_14905 ( .C (clk), .D (signal_19792), .Q (signal_19793) ) ;
    buf_clk cell_14911 ( .C (clk), .D (signal_19798), .Q (signal_19799) ) ;
    buf_clk cell_14917 ( .C (clk), .D (signal_19804), .Q (signal_19805) ) ;
    buf_clk cell_14923 ( .C (clk), .D (signal_19810), .Q (signal_19811) ) ;
    buf_clk cell_14929 ( .C (clk), .D (signal_19816), .Q (signal_19817) ) ;
    buf_clk cell_14935 ( .C (clk), .D (signal_19822), .Q (signal_19823) ) ;
    buf_clk cell_14941 ( .C (clk), .D (signal_19828), .Q (signal_19829) ) ;
    buf_clk cell_14947 ( .C (clk), .D (signal_19834), .Q (signal_19835) ) ;
    buf_clk cell_14953 ( .C (clk), .D (signal_19840), .Q (signal_19841) ) ;
    buf_clk cell_14959 ( .C (clk), .D (signal_19846), .Q (signal_19847) ) ;
    buf_clk cell_14965 ( .C (clk), .D (signal_19852), .Q (signal_19853) ) ;
    buf_clk cell_14971 ( .C (clk), .D (signal_19858), .Q (signal_19859) ) ;
    buf_clk cell_14977 ( .C (clk), .D (signal_19864), .Q (signal_19865) ) ;
    buf_clk cell_14983 ( .C (clk), .D (signal_19870), .Q (signal_19871) ) ;
    buf_clk cell_14989 ( .C (clk), .D (signal_19876), .Q (signal_19877) ) ;
    buf_clk cell_14995 ( .C (clk), .D (signal_19882), .Q (signal_19883) ) ;
    buf_clk cell_15001 ( .C (clk), .D (signal_19888), .Q (signal_19889) ) ;
    buf_clk cell_15007 ( .C (clk), .D (signal_19894), .Q (signal_19895) ) ;
    buf_clk cell_15013 ( .C (clk), .D (signal_19900), .Q (signal_19901) ) ;
    buf_clk cell_15019 ( .C (clk), .D (signal_19906), .Q (signal_19907) ) ;
    buf_clk cell_15025 ( .C (clk), .D (signal_19912), .Q (signal_19913) ) ;
    buf_clk cell_15031 ( .C (clk), .D (signal_19918), .Q (signal_19919) ) ;
    buf_clk cell_15037 ( .C (clk), .D (signal_19924), .Q (signal_19925) ) ;
    buf_clk cell_15043 ( .C (clk), .D (signal_19930), .Q (signal_19931) ) ;
    buf_clk cell_15049 ( .C (clk), .D (signal_19936), .Q (signal_19937) ) ;
    buf_clk cell_15055 ( .C (clk), .D (signal_19942), .Q (signal_19943) ) ;
    buf_clk cell_15061 ( .C (clk), .D (signal_19948), .Q (signal_19949) ) ;
    buf_clk cell_15067 ( .C (clk), .D (signal_19954), .Q (signal_19955) ) ;
    buf_clk cell_15073 ( .C (clk), .D (signal_19960), .Q (signal_19961) ) ;
    buf_clk cell_15079 ( .C (clk), .D (signal_19966), .Q (signal_19967) ) ;
    buf_clk cell_15085 ( .C (clk), .D (signal_19972), .Q (signal_19973) ) ;
    buf_clk cell_15091 ( .C (clk), .D (signal_19978), .Q (signal_19979) ) ;
    buf_clk cell_15097 ( .C (clk), .D (signal_19984), .Q (signal_19985) ) ;
    buf_clk cell_15103 ( .C (clk), .D (signal_19990), .Q (signal_19991) ) ;
    buf_clk cell_15109 ( .C (clk), .D (signal_19996), .Q (signal_19997) ) ;
    buf_clk cell_15115 ( .C (clk), .D (signal_20002), .Q (signal_20003) ) ;
    buf_clk cell_15121 ( .C (clk), .D (signal_20008), .Q (signal_20009) ) ;
    buf_clk cell_15127 ( .C (clk), .D (signal_20014), .Q (signal_20015) ) ;
    buf_clk cell_15133 ( .C (clk), .D (signal_20020), .Q (signal_20021) ) ;
    buf_clk cell_15139 ( .C (clk), .D (signal_20026), .Q (signal_20027) ) ;
    buf_clk cell_15145 ( .C (clk), .D (signal_20032), .Q (signal_20033) ) ;
    buf_clk cell_15151 ( .C (clk), .D (signal_20038), .Q (signal_20039) ) ;
    buf_clk cell_15157 ( .C (clk), .D (signal_20044), .Q (signal_20045) ) ;
    buf_clk cell_15163 ( .C (clk), .D (signal_20050), .Q (signal_20051) ) ;
    buf_clk cell_15169 ( .C (clk), .D (signal_20056), .Q (signal_20057) ) ;
    buf_clk cell_15175 ( .C (clk), .D (signal_20062), .Q (signal_20063) ) ;
    buf_clk cell_15181 ( .C (clk), .D (signal_20068), .Q (signal_20069) ) ;
    buf_clk cell_15187 ( .C (clk), .D (signal_20074), .Q (signal_20075) ) ;
    buf_clk cell_15193 ( .C (clk), .D (signal_20080), .Q (signal_20081) ) ;
    buf_clk cell_15199 ( .C (clk), .D (signal_20086), .Q (signal_20087) ) ;
    buf_clk cell_15205 ( .C (clk), .D (signal_20092), .Q (signal_20093) ) ;
    buf_clk cell_15211 ( .C (clk), .D (signal_20098), .Q (signal_20099) ) ;
    buf_clk cell_15217 ( .C (clk), .D (signal_20104), .Q (signal_20105) ) ;
    buf_clk cell_15223 ( .C (clk), .D (signal_20110), .Q (signal_20111) ) ;
    buf_clk cell_15229 ( .C (clk), .D (signal_20116), .Q (signal_20117) ) ;
    buf_clk cell_15235 ( .C (clk), .D (signal_20122), .Q (signal_20123) ) ;
    buf_clk cell_15241 ( .C (clk), .D (signal_20128), .Q (signal_20129) ) ;
    buf_clk cell_15247 ( .C (clk), .D (signal_20134), .Q (signal_20135) ) ;
    buf_clk cell_15253 ( .C (clk), .D (signal_20140), .Q (signal_20141) ) ;
    buf_clk cell_15259 ( .C (clk), .D (signal_20146), .Q (signal_20147) ) ;
    buf_clk cell_15265 ( .C (clk), .D (signal_20152), .Q (signal_20153) ) ;
    buf_clk cell_15271 ( .C (clk), .D (signal_20158), .Q (signal_20159) ) ;
    buf_clk cell_15277 ( .C (clk), .D (signal_20164), .Q (signal_20165) ) ;
    buf_clk cell_15283 ( .C (clk), .D (signal_20170), .Q (signal_20171) ) ;
    buf_clk cell_15289 ( .C (clk), .D (signal_20176), .Q (signal_20177) ) ;
    buf_clk cell_15295 ( .C (clk), .D (signal_20182), .Q (signal_20183) ) ;
    buf_clk cell_15301 ( .C (clk), .D (signal_20188), .Q (signal_20189) ) ;
    buf_clk cell_15307 ( .C (clk), .D (signal_20194), .Q (signal_20195) ) ;
    buf_clk cell_15313 ( .C (clk), .D (signal_20200), .Q (signal_20201) ) ;
    buf_clk cell_15319 ( .C (clk), .D (signal_20206), .Q (signal_20207) ) ;
    buf_clk cell_15325 ( .C (clk), .D (signal_20212), .Q (signal_20213) ) ;
    buf_clk cell_15331 ( .C (clk), .D (signal_20218), .Q (signal_20219) ) ;
    buf_clk cell_15337 ( .C (clk), .D (signal_20224), .Q (signal_20225) ) ;
    buf_clk cell_15343 ( .C (clk), .D (signal_20230), .Q (signal_20231) ) ;
    buf_clk cell_15349 ( .C (clk), .D (signal_20236), .Q (signal_20237) ) ;
    buf_clk cell_15355 ( .C (clk), .D (signal_20242), .Q (signal_20243) ) ;
    buf_clk cell_15361 ( .C (clk), .D (signal_20248), .Q (signal_20249) ) ;
    buf_clk cell_15367 ( .C (clk), .D (signal_20254), .Q (signal_20255) ) ;
    buf_clk cell_15373 ( .C (clk), .D (signal_20260), .Q (signal_20261) ) ;
    buf_clk cell_15379 ( .C (clk), .D (signal_20266), .Q (signal_20267) ) ;
    buf_clk cell_15385 ( .C (clk), .D (signal_20272), .Q (signal_20273) ) ;
    buf_clk cell_15391 ( .C (clk), .D (signal_20278), .Q (signal_20279) ) ;
    buf_clk cell_15397 ( .C (clk), .D (signal_20284), .Q (signal_20285) ) ;
    buf_clk cell_15403 ( .C (clk), .D (signal_20290), .Q (signal_20291) ) ;
    buf_clk cell_15409 ( .C (clk), .D (signal_20296), .Q (signal_20297) ) ;
    buf_clk cell_15415 ( .C (clk), .D (signal_20302), .Q (signal_20303) ) ;
    buf_clk cell_15421 ( .C (clk), .D (signal_20308), .Q (signal_20309) ) ;
    buf_clk cell_15427 ( .C (clk), .D (signal_20314), .Q (signal_20315) ) ;
    buf_clk cell_15433 ( .C (clk), .D (signal_20320), .Q (signal_20321) ) ;
    buf_clk cell_15439 ( .C (clk), .D (signal_20326), .Q (signal_20327) ) ;
    buf_clk cell_15445 ( .C (clk), .D (signal_20332), .Q (signal_20333) ) ;
    buf_clk cell_15451 ( .C (clk), .D (signal_20338), .Q (signal_20339) ) ;
    buf_clk cell_15457 ( .C (clk), .D (signal_20344), .Q (signal_20345) ) ;
    buf_clk cell_15463 ( .C (clk), .D (signal_20350), .Q (signal_20351) ) ;
    buf_clk cell_15469 ( .C (clk), .D (signal_20356), .Q (signal_20357) ) ;
    buf_clk cell_15475 ( .C (clk), .D (signal_20362), .Q (signal_20363) ) ;
    buf_clk cell_15481 ( .C (clk), .D (signal_20368), .Q (signal_20369) ) ;
    buf_clk cell_15487 ( .C (clk), .D (signal_20374), .Q (signal_20375) ) ;
    buf_clk cell_15493 ( .C (clk), .D (signal_20380), .Q (signal_20381) ) ;
    buf_clk cell_15499 ( .C (clk), .D (signal_20386), .Q (signal_20387) ) ;
    buf_clk cell_15505 ( .C (clk), .D (signal_20392), .Q (signal_20393) ) ;
    buf_clk cell_15511 ( .C (clk), .D (signal_20398), .Q (signal_20399) ) ;
    buf_clk cell_15517 ( .C (clk), .D (signal_20404), .Q (signal_20405) ) ;
    buf_clk cell_15523 ( .C (clk), .D (signal_20410), .Q (signal_20411) ) ;
    buf_clk cell_15529 ( .C (clk), .D (signal_20416), .Q (signal_20417) ) ;
    buf_clk cell_15535 ( .C (clk), .D (signal_20422), .Q (signal_20423) ) ;
    buf_clk cell_15541 ( .C (clk), .D (signal_20428), .Q (signal_20429) ) ;
    buf_clk cell_15547 ( .C (clk), .D (signal_20434), .Q (signal_20435) ) ;
    buf_clk cell_15553 ( .C (clk), .D (signal_20440), .Q (signal_20441) ) ;
    buf_clk cell_15559 ( .C (clk), .D (signal_20446), .Q (signal_20447) ) ;
    buf_clk cell_15565 ( .C (clk), .D (signal_20452), .Q (signal_20453) ) ;
    buf_clk cell_15571 ( .C (clk), .D (signal_20458), .Q (signal_20459) ) ;
    buf_clk cell_15577 ( .C (clk), .D (signal_20464), .Q (signal_20465) ) ;
    buf_clk cell_15583 ( .C (clk), .D (signal_20470), .Q (signal_20471) ) ;
    buf_clk cell_15589 ( .C (clk), .D (signal_20476), .Q (signal_20477) ) ;
    buf_clk cell_15595 ( .C (clk), .D (signal_20482), .Q (signal_20483) ) ;
    buf_clk cell_15601 ( .C (clk), .D (signal_20488), .Q (signal_20489) ) ;
    buf_clk cell_15607 ( .C (clk), .D (signal_20494), .Q (signal_20495) ) ;
    buf_clk cell_15613 ( .C (clk), .D (signal_20500), .Q (signal_20501) ) ;
    buf_clk cell_15619 ( .C (clk), .D (signal_20506), .Q (signal_20507) ) ;
    buf_clk cell_15625 ( .C (clk), .D (signal_20512), .Q (signal_20513) ) ;
    buf_clk cell_15631 ( .C (clk), .D (signal_20518), .Q (signal_20519) ) ;
    buf_clk cell_15637 ( .C (clk), .D (signal_20524), .Q (signal_20525) ) ;
    buf_clk cell_15643 ( .C (clk), .D (signal_20530), .Q (signal_20531) ) ;
    buf_clk cell_15649 ( .C (clk), .D (signal_20536), .Q (signal_20537) ) ;
    buf_clk cell_15655 ( .C (clk), .D (signal_20542), .Q (signal_20543) ) ;
    buf_clk cell_15661 ( .C (clk), .D (signal_20548), .Q (signal_20549) ) ;
    buf_clk cell_15667 ( .C (clk), .D (signal_20554), .Q (signal_20555) ) ;
    buf_clk cell_15673 ( .C (clk), .D (signal_20560), .Q (signal_20561) ) ;
    buf_clk cell_15679 ( .C (clk), .D (signal_20566), .Q (signal_20567) ) ;
    buf_clk cell_15685 ( .C (clk), .D (signal_20572), .Q (signal_20573) ) ;
    buf_clk cell_15691 ( .C (clk), .D (signal_20578), .Q (signal_20579) ) ;
    buf_clk cell_15697 ( .C (clk), .D (signal_20584), .Q (signal_20585) ) ;
    buf_clk cell_15703 ( .C (clk), .D (signal_20590), .Q (signal_20591) ) ;
    buf_clk cell_15709 ( .C (clk), .D (signal_20596), .Q (signal_20597) ) ;
    buf_clk cell_15715 ( .C (clk), .D (signal_20602), .Q (signal_20603) ) ;
    buf_clk cell_15721 ( .C (clk), .D (signal_20608), .Q (signal_20609) ) ;
    buf_clk cell_15727 ( .C (clk), .D (signal_20614), .Q (signal_20615) ) ;
    buf_clk cell_15733 ( .C (clk), .D (signal_20620), .Q (signal_20621) ) ;
    buf_clk cell_15739 ( .C (clk), .D (signal_20626), .Q (signal_20627) ) ;
    buf_clk cell_15745 ( .C (clk), .D (signal_20632), .Q (signal_20633) ) ;
    buf_clk cell_15751 ( .C (clk), .D (signal_20638), .Q (signal_20639) ) ;
    buf_clk cell_15757 ( .C (clk), .D (signal_20644), .Q (signal_20645) ) ;
    buf_clk cell_15763 ( .C (clk), .D (signal_20650), .Q (signal_20651) ) ;
    buf_clk cell_15769 ( .C (clk), .D (signal_20656), .Q (signal_20657) ) ;
    buf_clk cell_15775 ( .C (clk), .D (signal_20662), .Q (signal_20663) ) ;
    buf_clk cell_15781 ( .C (clk), .D (signal_20668), .Q (signal_20669) ) ;
    buf_clk cell_15787 ( .C (clk), .D (signal_20674), .Q (signal_20675) ) ;
    buf_clk cell_15793 ( .C (clk), .D (signal_20680), .Q (signal_20681) ) ;
    buf_clk cell_15799 ( .C (clk), .D (signal_20686), .Q (signal_20687) ) ;
    buf_clk cell_15805 ( .C (clk), .D (signal_20692), .Q (signal_20693) ) ;
    buf_clk cell_15811 ( .C (clk), .D (signal_20698), .Q (signal_20699) ) ;
    buf_clk cell_15817 ( .C (clk), .D (signal_20704), .Q (signal_20705) ) ;
    buf_clk cell_15823 ( .C (clk), .D (signal_20710), .Q (signal_20711) ) ;
    buf_clk cell_15829 ( .C (clk), .D (signal_20716), .Q (signal_20717) ) ;
    buf_clk cell_15835 ( .C (clk), .D (signal_20722), .Q (signal_20723) ) ;
    buf_clk cell_15841 ( .C (clk), .D (signal_20728), .Q (signal_20729) ) ;
    buf_clk cell_15847 ( .C (clk), .D (signal_20734), .Q (signal_20735) ) ;
    buf_clk cell_15853 ( .C (clk), .D (signal_20740), .Q (signal_20741) ) ;
    buf_clk cell_15859 ( .C (clk), .D (signal_20746), .Q (signal_20747) ) ;
    buf_clk cell_15865 ( .C (clk), .D (signal_20752), .Q (signal_20753) ) ;
    buf_clk cell_15871 ( .C (clk), .D (signal_20758), .Q (signal_20759) ) ;
    buf_clk cell_15877 ( .C (clk), .D (signal_20764), .Q (signal_20765) ) ;
    buf_clk cell_15883 ( .C (clk), .D (signal_20770), .Q (signal_20771) ) ;
    buf_clk cell_15889 ( .C (clk), .D (signal_20776), .Q (signal_20777) ) ;
    buf_clk cell_15895 ( .C (clk), .D (signal_20782), .Q (signal_20783) ) ;
    buf_clk cell_15901 ( .C (clk), .D (signal_20788), .Q (signal_20789) ) ;
    buf_clk cell_15907 ( .C (clk), .D (signal_20794), .Q (signal_20795) ) ;
    buf_clk cell_15913 ( .C (clk), .D (signal_20800), .Q (signal_20801) ) ;
    buf_clk cell_15919 ( .C (clk), .D (signal_20806), .Q (signal_20807) ) ;
    buf_clk cell_15925 ( .C (clk), .D (signal_20812), .Q (signal_20813) ) ;
    buf_clk cell_15931 ( .C (clk), .D (signal_20818), .Q (signal_20819) ) ;
    buf_clk cell_15937 ( .C (clk), .D (signal_20824), .Q (signal_20825) ) ;
    buf_clk cell_15943 ( .C (clk), .D (signal_20830), .Q (signal_20831) ) ;
    buf_clk cell_15949 ( .C (clk), .D (signal_20836), .Q (signal_20837) ) ;
    buf_clk cell_15955 ( .C (clk), .D (signal_20842), .Q (signal_20843) ) ;
    buf_clk cell_15961 ( .C (clk), .D (signal_20848), .Q (signal_20849) ) ;
    buf_clk cell_15967 ( .C (clk), .D (signal_20854), .Q (signal_20855) ) ;
    buf_clk cell_15973 ( .C (clk), .D (signal_20860), .Q (signal_20861) ) ;
    buf_clk cell_15979 ( .C (clk), .D (signal_20866), .Q (signal_20867) ) ;
    buf_clk cell_15985 ( .C (clk), .D (signal_20872), .Q (signal_20873) ) ;
    buf_clk cell_15991 ( .C (clk), .D (signal_20878), .Q (signal_20879) ) ;
    buf_clk cell_15997 ( .C (clk), .D (signal_20884), .Q (signal_20885) ) ;
    buf_clk cell_16003 ( .C (clk), .D (signal_20890), .Q (signal_20891) ) ;
    buf_clk cell_16009 ( .C (clk), .D (signal_20896), .Q (signal_20897) ) ;
    buf_clk cell_16015 ( .C (clk), .D (signal_20902), .Q (signal_20903) ) ;
    buf_clk cell_16021 ( .C (clk), .D (signal_20908), .Q (signal_20909) ) ;
    buf_clk cell_16027 ( .C (clk), .D (signal_20914), .Q (signal_20915) ) ;
    buf_clk cell_16033 ( .C (clk), .D (signal_20920), .Q (signal_20921) ) ;
    buf_clk cell_16039 ( .C (clk), .D (signal_20926), .Q (signal_20927) ) ;
    buf_clk cell_16045 ( .C (clk), .D (signal_20932), .Q (signal_20933) ) ;
    buf_clk cell_16051 ( .C (clk), .D (signal_20938), .Q (signal_20939) ) ;
    buf_clk cell_16057 ( .C (clk), .D (signal_20944), .Q (signal_20945) ) ;
    buf_clk cell_16063 ( .C (clk), .D (signal_20950), .Q (signal_20951) ) ;
    buf_clk cell_16069 ( .C (clk), .D (signal_20956), .Q (signal_20957) ) ;
    buf_clk cell_16075 ( .C (clk), .D (signal_20962), .Q (signal_20963) ) ;
    buf_clk cell_16081 ( .C (clk), .D (signal_20968), .Q (signal_20969) ) ;
    buf_clk cell_16087 ( .C (clk), .D (signal_20974), .Q (signal_20975) ) ;
    buf_clk cell_16093 ( .C (clk), .D (signal_20980), .Q (signal_20981) ) ;
    buf_clk cell_16099 ( .C (clk), .D (signal_20986), .Q (signal_20987) ) ;
    buf_clk cell_16105 ( .C (clk), .D (signal_20992), .Q (signal_20993) ) ;
    buf_clk cell_16111 ( .C (clk), .D (signal_20998), .Q (signal_20999) ) ;
    buf_clk cell_16117 ( .C (clk), .D (signal_21004), .Q (signal_21005) ) ;
    buf_clk cell_16123 ( .C (clk), .D (signal_21010), .Q (signal_21011) ) ;
    buf_clk cell_16129 ( .C (clk), .D (signal_21016), .Q (signal_21017) ) ;
    buf_clk cell_16135 ( .C (clk), .D (signal_21022), .Q (signal_21023) ) ;
    buf_clk cell_16141 ( .C (clk), .D (signal_21028), .Q (signal_21029) ) ;
    buf_clk cell_16147 ( .C (clk), .D (signal_21034), .Q (signal_21035) ) ;
    buf_clk cell_16153 ( .C (clk), .D (signal_21040), .Q (signal_21041) ) ;
    buf_clk cell_16159 ( .C (clk), .D (signal_21046), .Q (signal_21047) ) ;
    buf_clk cell_16165 ( .C (clk), .D (signal_21052), .Q (signal_21053) ) ;
    buf_clk cell_16171 ( .C (clk), .D (signal_21058), .Q (signal_21059) ) ;
    buf_clk cell_16177 ( .C (clk), .D (signal_21064), .Q (signal_21065) ) ;
    buf_clk cell_16183 ( .C (clk), .D (signal_21070), .Q (signal_21071) ) ;
    buf_clk cell_16189 ( .C (clk), .D (signal_21076), .Q (signal_21077) ) ;
    buf_clk cell_16195 ( .C (clk), .D (signal_21082), .Q (signal_21083) ) ;
    buf_clk cell_16201 ( .C (clk), .D (signal_21088), .Q (signal_21089) ) ;
    buf_clk cell_16207 ( .C (clk), .D (signal_21094), .Q (signal_21095) ) ;
    buf_clk cell_16213 ( .C (clk), .D (signal_21100), .Q (signal_21101) ) ;
    buf_clk cell_16219 ( .C (clk), .D (signal_21106), .Q (signal_21107) ) ;
    buf_clk cell_16225 ( .C (clk), .D (signal_21112), .Q (signal_21113) ) ;
    buf_clk cell_16231 ( .C (clk), .D (signal_21118), .Q (signal_21119) ) ;
    buf_clk cell_16237 ( .C (clk), .D (signal_21124), .Q (signal_21125) ) ;
    buf_clk cell_16243 ( .C (clk), .D (signal_21130), .Q (signal_21131) ) ;
    buf_clk cell_16249 ( .C (clk), .D (signal_21136), .Q (signal_21137) ) ;
    buf_clk cell_16255 ( .C (clk), .D (signal_21142), .Q (signal_21143) ) ;
    buf_clk cell_16261 ( .C (clk), .D (signal_21148), .Q (signal_21149) ) ;
    buf_clk cell_16267 ( .C (clk), .D (signal_21154), .Q (signal_21155) ) ;
    buf_clk cell_16273 ( .C (clk), .D (signal_21160), .Q (signal_21161) ) ;
    buf_clk cell_16279 ( .C (clk), .D (signal_21166), .Q (signal_21167) ) ;
    buf_clk cell_16285 ( .C (clk), .D (signal_21172), .Q (signal_21173) ) ;
    buf_clk cell_16291 ( .C (clk), .D (signal_21178), .Q (signal_21179) ) ;
    buf_clk cell_16297 ( .C (clk), .D (signal_21184), .Q (signal_21185) ) ;
    buf_clk cell_16303 ( .C (clk), .D (signal_21190), .Q (signal_21191) ) ;
    buf_clk cell_16309 ( .C (clk), .D (signal_21196), .Q (signal_21197) ) ;
    buf_clk cell_16315 ( .C (clk), .D (signal_21202), .Q (signal_21203) ) ;
    buf_clk cell_16321 ( .C (clk), .D (signal_21208), .Q (signal_21209) ) ;
    buf_clk cell_16327 ( .C (clk), .D (signal_21214), .Q (signal_21215) ) ;
    buf_clk cell_16333 ( .C (clk), .D (signal_21220), .Q (signal_21221) ) ;
    buf_clk cell_16339 ( .C (clk), .D (signal_21226), .Q (signal_21227) ) ;
    buf_clk cell_16345 ( .C (clk), .D (signal_21232), .Q (signal_21233) ) ;
    buf_clk cell_16351 ( .C (clk), .D (signal_21238), .Q (signal_21239) ) ;
    buf_clk cell_16357 ( .C (clk), .D (signal_21244), .Q (signal_21245) ) ;
    buf_clk cell_16363 ( .C (clk), .D (signal_21250), .Q (signal_21251) ) ;
    buf_clk cell_16369 ( .C (clk), .D (signal_21256), .Q (signal_21257) ) ;
    buf_clk cell_16375 ( .C (clk), .D (signal_21262), .Q (signal_21263) ) ;
    buf_clk cell_16381 ( .C (clk), .D (signal_21268), .Q (signal_21269) ) ;
    buf_clk cell_16387 ( .C (clk), .D (signal_21274), .Q (signal_21275) ) ;
    buf_clk cell_16393 ( .C (clk), .D (signal_21280), .Q (signal_21281) ) ;
    buf_clk cell_16399 ( .C (clk), .D (signal_21286), .Q (signal_21287) ) ;
    buf_clk cell_16405 ( .C (clk), .D (signal_21292), .Q (signal_21293) ) ;
    buf_clk cell_16411 ( .C (clk), .D (signal_21298), .Q (signal_21299) ) ;
    buf_clk cell_16417 ( .C (clk), .D (signal_21304), .Q (signal_21305) ) ;
    buf_clk cell_16423 ( .C (clk), .D (signal_21310), .Q (signal_21311) ) ;
    buf_clk cell_16429 ( .C (clk), .D (signal_21316), .Q (signal_21317) ) ;
    buf_clk cell_16435 ( .C (clk), .D (signal_21322), .Q (signal_21323) ) ;
    buf_clk cell_16441 ( .C (clk), .D (signal_21328), .Q (signal_21329) ) ;
    buf_clk cell_16447 ( .C (clk), .D (signal_21334), .Q (signal_21335) ) ;
    buf_clk cell_16453 ( .C (clk), .D (signal_21340), .Q (signal_21341) ) ;
    buf_clk cell_16459 ( .C (clk), .D (signal_21346), .Q (signal_21347) ) ;
    buf_clk cell_16465 ( .C (clk), .D (signal_21352), .Q (signal_21353) ) ;
    buf_clk cell_16471 ( .C (clk), .D (signal_21358), .Q (signal_21359) ) ;
    buf_clk cell_16477 ( .C (clk), .D (signal_21364), .Q (signal_21365) ) ;
    buf_clk cell_16483 ( .C (clk), .D (signal_21370), .Q (signal_21371) ) ;
    buf_clk cell_16489 ( .C (clk), .D (signal_21376), .Q (signal_21377) ) ;
    buf_clk cell_16495 ( .C (clk), .D (signal_21382), .Q (signal_21383) ) ;
    buf_clk cell_16501 ( .C (clk), .D (signal_21388), .Q (signal_21389) ) ;
    buf_clk cell_16507 ( .C (clk), .D (signal_21394), .Q (signal_21395) ) ;
    buf_clk cell_16513 ( .C (clk), .D (signal_21400), .Q (signal_21401) ) ;
    buf_clk cell_16519 ( .C (clk), .D (signal_21406), .Q (signal_21407) ) ;
    buf_clk cell_16525 ( .C (clk), .D (signal_21412), .Q (signal_21413) ) ;
    buf_clk cell_16531 ( .C (clk), .D (signal_21418), .Q (signal_21419) ) ;
    buf_clk cell_16537 ( .C (clk), .D (signal_21424), .Q (signal_21425) ) ;
    buf_clk cell_16543 ( .C (clk), .D (signal_21430), .Q (signal_21431) ) ;
    buf_clk cell_16549 ( .C (clk), .D (signal_21436), .Q (signal_21437) ) ;
    buf_clk cell_16555 ( .C (clk), .D (signal_21442), .Q (signal_21443) ) ;
    buf_clk cell_16561 ( .C (clk), .D (signal_21448), .Q (signal_21449) ) ;
    buf_clk cell_16567 ( .C (clk), .D (signal_21454), .Q (signal_21455) ) ;
    buf_clk cell_16573 ( .C (clk), .D (signal_21460), .Q (signal_21461) ) ;
    buf_clk cell_16579 ( .C (clk), .D (signal_21466), .Q (signal_21467) ) ;
    buf_clk cell_16585 ( .C (clk), .D (signal_21472), .Q (signal_21473) ) ;
    buf_clk cell_16591 ( .C (clk), .D (signal_21478), .Q (signal_21479) ) ;
    buf_clk cell_16597 ( .C (clk), .D (signal_21484), .Q (signal_21485) ) ;
    buf_clk cell_16603 ( .C (clk), .D (signal_21490), .Q (signal_21491) ) ;
    buf_clk cell_16609 ( .C (clk), .D (signal_21496), .Q (signal_21497) ) ;
    buf_clk cell_16615 ( .C (clk), .D (signal_21502), .Q (signal_21503) ) ;
    buf_clk cell_16621 ( .C (clk), .D (signal_21508), .Q (signal_21509) ) ;
    buf_clk cell_16627 ( .C (clk), .D (signal_21514), .Q (signal_21515) ) ;
    buf_clk cell_16633 ( .C (clk), .D (signal_21520), .Q (signal_21521) ) ;
    buf_clk cell_16639 ( .C (clk), .D (signal_21526), .Q (signal_21527) ) ;
    buf_clk cell_16645 ( .C (clk), .D (signal_21532), .Q (signal_21533) ) ;
    buf_clk cell_16651 ( .C (clk), .D (signal_21538), .Q (signal_21539) ) ;
    buf_clk cell_16657 ( .C (clk), .D (signal_21544), .Q (signal_21545) ) ;
    buf_clk cell_16663 ( .C (clk), .D (signal_21550), .Q (signal_21551) ) ;
    buf_clk cell_16669 ( .C (clk), .D (signal_21556), .Q (signal_21557) ) ;
    buf_clk cell_16675 ( .C (clk), .D (signal_21562), .Q (signal_21563) ) ;
    buf_clk cell_16681 ( .C (clk), .D (signal_21568), .Q (signal_21569) ) ;
    buf_clk cell_16687 ( .C (clk), .D (signal_21574), .Q (signal_21575) ) ;
    buf_clk cell_16693 ( .C (clk), .D (signal_21580), .Q (signal_21581) ) ;
    buf_clk cell_16699 ( .C (clk), .D (signal_21586), .Q (signal_21587) ) ;
    buf_clk cell_16705 ( .C (clk), .D (signal_21592), .Q (signal_21593) ) ;
    buf_clk cell_16711 ( .C (clk), .D (signal_21598), .Q (signal_21599) ) ;
    buf_clk cell_16717 ( .C (clk), .D (signal_21604), .Q (signal_21605) ) ;
    buf_clk cell_16723 ( .C (clk), .D (signal_21610), .Q (signal_21611) ) ;
    buf_clk cell_16729 ( .C (clk), .D (signal_21616), .Q (signal_21617) ) ;
    buf_clk cell_16735 ( .C (clk), .D (signal_21622), .Q (signal_21623) ) ;
    buf_clk cell_16741 ( .C (clk), .D (signal_21628), .Q (signal_21629) ) ;
    buf_clk cell_16747 ( .C (clk), .D (signal_21634), .Q (signal_21635) ) ;
    buf_clk cell_16753 ( .C (clk), .D (signal_21640), .Q (signal_21641) ) ;
    buf_clk cell_16759 ( .C (clk), .D (signal_21646), .Q (signal_21647) ) ;
    buf_clk cell_16765 ( .C (clk), .D (signal_21652), .Q (signal_21653) ) ;
    buf_clk cell_16771 ( .C (clk), .D (signal_21658), .Q (signal_21659) ) ;
    buf_clk cell_16777 ( .C (clk), .D (signal_21664), .Q (signal_21665) ) ;
    buf_clk cell_16783 ( .C (clk), .D (signal_21670), .Q (signal_21671) ) ;
    buf_clk cell_16789 ( .C (clk), .D (signal_21676), .Q (signal_21677) ) ;
    buf_clk cell_16795 ( .C (clk), .D (signal_21682), .Q (signal_21683) ) ;
    buf_clk cell_16801 ( .C (clk), .D (signal_21688), .Q (signal_21689) ) ;
    buf_clk cell_16807 ( .C (clk), .D (signal_21694), .Q (signal_21695) ) ;
    buf_clk cell_16813 ( .C (clk), .D (signal_21700), .Q (signal_21701) ) ;
    buf_clk cell_16819 ( .C (clk), .D (signal_21706), .Q (signal_21707) ) ;
    buf_clk cell_16825 ( .C (clk), .D (signal_21712), .Q (signal_21713) ) ;
    buf_clk cell_16831 ( .C (clk), .D (signal_21718), .Q (signal_21719) ) ;
    buf_clk cell_16837 ( .C (clk), .D (signal_21724), .Q (signal_21725) ) ;
    buf_clk cell_16843 ( .C (clk), .D (signal_21730), .Q (signal_21731) ) ;
    buf_clk cell_16849 ( .C (clk), .D (signal_21736), .Q (signal_21737) ) ;
    buf_clk cell_16855 ( .C (clk), .D (signal_21742), .Q (signal_21743) ) ;
    buf_clk cell_16861 ( .C (clk), .D (signal_21748), .Q (signal_21749) ) ;
    buf_clk cell_16867 ( .C (clk), .D (signal_21754), .Q (signal_21755) ) ;
    buf_clk cell_16873 ( .C (clk), .D (signal_21760), .Q (signal_21761) ) ;
    buf_clk cell_16879 ( .C (clk), .D (signal_21766), .Q (signal_21767) ) ;
    buf_clk cell_16885 ( .C (clk), .D (signal_21772), .Q (signal_21773) ) ;
    buf_clk cell_16891 ( .C (clk), .D (signal_21778), .Q (signal_21779) ) ;
    buf_clk cell_16897 ( .C (clk), .D (signal_21784), .Q (signal_21785) ) ;
    buf_clk cell_16903 ( .C (clk), .D (signal_21790), .Q (signal_21791) ) ;
    buf_clk cell_16909 ( .C (clk), .D (signal_21796), .Q (signal_21797) ) ;
    buf_clk cell_16915 ( .C (clk), .D (signal_21802), .Q (signal_21803) ) ;
    buf_clk cell_16921 ( .C (clk), .D (signal_21808), .Q (signal_21809) ) ;
    buf_clk cell_16927 ( .C (clk), .D (signal_21814), .Q (signal_21815) ) ;
    buf_clk cell_16933 ( .C (clk), .D (signal_21820), .Q (signal_21821) ) ;
    buf_clk cell_16939 ( .C (clk), .D (signal_21826), .Q (signal_21827) ) ;
    buf_clk cell_16945 ( .C (clk), .D (signal_21832), .Q (signal_21833) ) ;
    buf_clk cell_16951 ( .C (clk), .D (signal_21838), .Q (signal_21839) ) ;
    buf_clk cell_16957 ( .C (clk), .D (signal_21844), .Q (signal_21845) ) ;
    buf_clk cell_16963 ( .C (clk), .D (signal_21850), .Q (signal_21851) ) ;
    buf_clk cell_16969 ( .C (clk), .D (signal_21856), .Q (signal_21857) ) ;
    buf_clk cell_16975 ( .C (clk), .D (signal_21862), .Q (signal_21863) ) ;
    buf_clk cell_16981 ( .C (clk), .D (signal_21868), .Q (signal_21869) ) ;
    buf_clk cell_16987 ( .C (clk), .D (signal_21874), .Q (signal_21875) ) ;
    buf_clk cell_16993 ( .C (clk), .D (signal_21880), .Q (signal_21881) ) ;
    buf_clk cell_16999 ( .C (clk), .D (signal_21886), .Q (signal_21887) ) ;
    buf_clk cell_17005 ( .C (clk), .D (signal_21892), .Q (signal_21893) ) ;
    buf_clk cell_17011 ( .C (clk), .D (signal_21898), .Q (signal_21899) ) ;
    buf_clk cell_17017 ( .C (clk), .D (signal_21904), .Q (signal_21905) ) ;
    buf_clk cell_17023 ( .C (clk), .D (signal_21910), .Q (signal_21911) ) ;
    buf_clk cell_17029 ( .C (clk), .D (signal_21916), .Q (signal_21917) ) ;
    buf_clk cell_17035 ( .C (clk), .D (signal_21922), .Q (signal_21923) ) ;
    buf_clk cell_17041 ( .C (clk), .D (signal_21928), .Q (signal_21929) ) ;
    buf_clk cell_17047 ( .C (clk), .D (signal_21934), .Q (signal_21935) ) ;
    buf_clk cell_17053 ( .C (clk), .D (signal_21940), .Q (signal_21941) ) ;
    buf_clk cell_17059 ( .C (clk), .D (signal_21946), .Q (signal_21947) ) ;
    buf_clk cell_17065 ( .C (clk), .D (signal_21952), .Q (signal_21953) ) ;
    buf_clk cell_17071 ( .C (clk), .D (signal_21958), .Q (signal_21959) ) ;
    buf_clk cell_17077 ( .C (clk), .D (signal_21964), .Q (signal_21965) ) ;
    buf_clk cell_17083 ( .C (clk), .D (signal_21970), .Q (signal_21971) ) ;
    buf_clk cell_17089 ( .C (clk), .D (signal_21976), .Q (signal_21977) ) ;
    buf_clk cell_17095 ( .C (clk), .D (signal_21982), .Q (signal_21983) ) ;
    buf_clk cell_17101 ( .C (clk), .D (signal_21988), .Q (signal_21989) ) ;
    buf_clk cell_17107 ( .C (clk), .D (signal_21994), .Q (signal_21995) ) ;
    buf_clk cell_17113 ( .C (clk), .D (signal_22000), .Q (signal_22001) ) ;
    buf_clk cell_17119 ( .C (clk), .D (signal_22006), .Q (signal_22007) ) ;
    buf_clk cell_17125 ( .C (clk), .D (signal_22012), .Q (signal_22013) ) ;
    buf_clk cell_17131 ( .C (clk), .D (signal_22018), .Q (signal_22019) ) ;
    buf_clk cell_17137 ( .C (clk), .D (signal_22024), .Q (signal_22025) ) ;
    buf_clk cell_17143 ( .C (clk), .D (signal_22030), .Q (signal_22031) ) ;
    buf_clk cell_17149 ( .C (clk), .D (signal_22036), .Q (signal_22037) ) ;
    buf_clk cell_17155 ( .C (clk), .D (signal_22042), .Q (signal_22043) ) ;
    buf_clk cell_17161 ( .C (clk), .D (signal_22048), .Q (signal_22049) ) ;
    buf_clk cell_17167 ( .C (clk), .D (signal_22054), .Q (signal_22055) ) ;
    buf_clk cell_17173 ( .C (clk), .D (signal_22060), .Q (signal_22061) ) ;
    buf_clk cell_17179 ( .C (clk), .D (signal_22066), .Q (signal_22067) ) ;
    buf_clk cell_17185 ( .C (clk), .D (signal_22072), .Q (signal_22073) ) ;
    buf_clk cell_17191 ( .C (clk), .D (signal_22078), .Q (signal_22079) ) ;
    buf_clk cell_17197 ( .C (clk), .D (signal_22084), .Q (signal_22085) ) ;
    buf_clk cell_17203 ( .C (clk), .D (signal_22090), .Q (signal_22091) ) ;
    buf_clk cell_17209 ( .C (clk), .D (signal_22096), .Q (signal_22097) ) ;
    buf_clk cell_17215 ( .C (clk), .D (signal_22102), .Q (signal_22103) ) ;
    buf_clk cell_17221 ( .C (clk), .D (signal_22108), .Q (signal_22109) ) ;
    buf_clk cell_17227 ( .C (clk), .D (signal_22114), .Q (signal_22115) ) ;
    buf_clk cell_17233 ( .C (clk), .D (signal_22120), .Q (signal_22121) ) ;
    buf_clk cell_17239 ( .C (clk), .D (signal_22126), .Q (signal_22127) ) ;
    buf_clk cell_17245 ( .C (clk), .D (signal_22132), .Q (signal_22133) ) ;
    buf_clk cell_17251 ( .C (clk), .D (signal_22138), .Q (signal_22139) ) ;
    buf_clk cell_17257 ( .C (clk), .D (signal_22144), .Q (signal_22145) ) ;
    buf_clk cell_17263 ( .C (clk), .D (signal_22150), .Q (signal_22151) ) ;
    buf_clk cell_17269 ( .C (clk), .D (signal_22156), .Q (signal_22157) ) ;
    buf_clk cell_17275 ( .C (clk), .D (signal_22162), .Q (signal_22163) ) ;
    buf_clk cell_17281 ( .C (clk), .D (signal_22168), .Q (signal_22169) ) ;
    buf_clk cell_17287 ( .C (clk), .D (signal_22174), .Q (signal_22175) ) ;
    buf_clk cell_17293 ( .C (clk), .D (signal_22180), .Q (signal_22181) ) ;
    buf_clk cell_17299 ( .C (clk), .D (signal_22186), .Q (signal_22187) ) ;
    buf_clk cell_17305 ( .C (clk), .D (signal_22192), .Q (signal_22193) ) ;
    buf_clk cell_17311 ( .C (clk), .D (signal_22198), .Q (signal_22199) ) ;
    buf_clk cell_17317 ( .C (clk), .D (signal_22204), .Q (signal_22205) ) ;
    buf_clk cell_17323 ( .C (clk), .D (signal_22210), .Q (signal_22211) ) ;
    buf_clk cell_17329 ( .C (clk), .D (signal_22216), .Q (signal_22217) ) ;
    buf_clk cell_17335 ( .C (clk), .D (signal_22222), .Q (signal_22223) ) ;
    buf_clk cell_17341 ( .C (clk), .D (signal_22228), .Q (signal_22229) ) ;
    buf_clk cell_17347 ( .C (clk), .D (signal_22234), .Q (signal_22235) ) ;
    buf_clk cell_17353 ( .C (clk), .D (signal_22240), .Q (signal_22241) ) ;
    buf_clk cell_17359 ( .C (clk), .D (signal_22246), .Q (signal_22247) ) ;
    buf_clk cell_17365 ( .C (clk), .D (signal_22252), .Q (signal_22253) ) ;
    buf_clk cell_17371 ( .C (clk), .D (signal_22258), .Q (signal_22259) ) ;
    buf_clk cell_17377 ( .C (clk), .D (signal_22264), .Q (signal_22265) ) ;
    buf_clk cell_17383 ( .C (clk), .D (signal_22270), .Q (signal_22271) ) ;
    buf_clk cell_17389 ( .C (clk), .D (signal_22276), .Q (signal_22277) ) ;
    buf_clk cell_17395 ( .C (clk), .D (signal_22282), .Q (signal_22283) ) ;
    buf_clk cell_17401 ( .C (clk), .D (signal_22288), .Q (signal_22289) ) ;
    buf_clk cell_17407 ( .C (clk), .D (signal_22294), .Q (signal_22295) ) ;
    buf_clk cell_17413 ( .C (clk), .D (signal_22300), .Q (signal_22301) ) ;
    buf_clk cell_17419 ( .C (clk), .D (signal_22306), .Q (signal_22307) ) ;
    buf_clk cell_17425 ( .C (clk), .D (signal_22312), .Q (signal_22313) ) ;
    buf_clk cell_17431 ( .C (clk), .D (signal_22318), .Q (signal_22319) ) ;
    buf_clk cell_17437 ( .C (clk), .D (signal_22324), .Q (signal_22325) ) ;
    buf_clk cell_17443 ( .C (clk), .D (signal_22330), .Q (signal_22331) ) ;
    buf_clk cell_17449 ( .C (clk), .D (signal_22336), .Q (signal_22337) ) ;
    buf_clk cell_17455 ( .C (clk), .D (signal_22342), .Q (signal_22343) ) ;
    buf_clk cell_17461 ( .C (clk), .D (signal_22348), .Q (signal_22349) ) ;
    buf_clk cell_17467 ( .C (clk), .D (signal_22354), .Q (signal_22355) ) ;
    buf_clk cell_17473 ( .C (clk), .D (signal_22360), .Q (signal_22361) ) ;
    buf_clk cell_17479 ( .C (clk), .D (signal_22366), .Q (signal_22367) ) ;
    buf_clk cell_17485 ( .C (clk), .D (signal_22372), .Q (signal_22373) ) ;
    buf_clk cell_17491 ( .C (clk), .D (signal_22378), .Q (signal_22379) ) ;
    buf_clk cell_17497 ( .C (clk), .D (signal_22384), .Q (signal_22385) ) ;
    buf_clk cell_17503 ( .C (clk), .D (signal_22390), .Q (signal_22391) ) ;
    buf_clk cell_17509 ( .C (clk), .D (signal_22396), .Q (signal_22397) ) ;
    buf_clk cell_17515 ( .C (clk), .D (signal_22402), .Q (signal_22403) ) ;
    buf_clk cell_17521 ( .C (clk), .D (signal_22408), .Q (signal_22409) ) ;
    buf_clk cell_17527 ( .C (clk), .D (signal_22414), .Q (signal_22415) ) ;
    buf_clk cell_17533 ( .C (clk), .D (signal_22420), .Q (signal_22421) ) ;
    buf_clk cell_17539 ( .C (clk), .D (signal_22426), .Q (signal_22427) ) ;
    buf_clk cell_17545 ( .C (clk), .D (signal_22432), .Q (signal_22433) ) ;
    buf_clk cell_17551 ( .C (clk), .D (signal_22438), .Q (signal_22439) ) ;
    buf_clk cell_17557 ( .C (clk), .D (signal_22444), .Q (signal_22445) ) ;
    buf_clk cell_17563 ( .C (clk), .D (signal_22450), .Q (signal_22451) ) ;
    buf_clk cell_17569 ( .C (clk), .D (signal_22456), .Q (signal_22457) ) ;
    buf_clk cell_17575 ( .C (clk), .D (signal_22462), .Q (signal_22463) ) ;
    buf_clk cell_17581 ( .C (clk), .D (signal_22468), .Q (signal_22469) ) ;
    buf_clk cell_17587 ( .C (clk), .D (signal_22474), .Q (signal_22475) ) ;
    buf_clk cell_17595 ( .C (clk), .D (signal_22482), .Q (signal_22483) ) ;
    buf_clk cell_17603 ( .C (clk), .D (signal_22490), .Q (signal_22491) ) ;
    buf_clk cell_17611 ( .C (clk), .D (signal_22498), .Q (signal_22499) ) ;
    buf_clk cell_17619 ( .C (clk), .D (signal_22506), .Q (signal_22507) ) ;
    buf_clk cell_17627 ( .C (clk), .D (signal_22514), .Q (signal_22515) ) ;
    buf_clk cell_17635 ( .C (clk), .D (signal_22522), .Q (signal_22523) ) ;
    buf_clk cell_17643 ( .C (clk), .D (signal_22530), .Q (signal_22531) ) ;
    buf_clk cell_17651 ( .C (clk), .D (signal_22538), .Q (signal_22539) ) ;
    buf_clk cell_17659 ( .C (clk), .D (signal_22546), .Q (signal_22547) ) ;
    buf_clk cell_17667 ( .C (clk), .D (signal_22554), .Q (signal_22555) ) ;
    buf_clk cell_17675 ( .C (clk), .D (signal_22562), .Q (signal_22563) ) ;
    buf_clk cell_17683 ( .C (clk), .D (signal_22570), .Q (signal_22571) ) ;
    buf_clk cell_17691 ( .C (clk), .D (signal_22578), .Q (signal_22579) ) ;
    buf_clk cell_17699 ( .C (clk), .D (signal_22586), .Q (signal_22587) ) ;
    buf_clk cell_17707 ( .C (clk), .D (signal_22594), .Q (signal_22595) ) ;
    buf_clk cell_17715 ( .C (clk), .D (signal_22602), .Q (signal_22603) ) ;
    buf_clk cell_17723 ( .C (clk), .D (signal_22610), .Q (signal_22611) ) ;
    buf_clk cell_17731 ( .C (clk), .D (signal_22618), .Q (signal_22619) ) ;
    buf_clk cell_17739 ( .C (clk), .D (signal_22626), .Q (signal_22627) ) ;
    buf_clk cell_17747 ( .C (clk), .D (signal_22634), .Q (signal_22635) ) ;
    buf_clk cell_17755 ( .C (clk), .D (signal_22642), .Q (signal_22643) ) ;
    buf_clk cell_17763 ( .C (clk), .D (signal_22650), .Q (signal_22651) ) ;
    buf_clk cell_17771 ( .C (clk), .D (signal_22658), .Q (signal_22659) ) ;
    buf_clk cell_17779 ( .C (clk), .D (signal_22666), .Q (signal_22667) ) ;
    buf_clk cell_17787 ( .C (clk), .D (signal_22674), .Q (signal_22675) ) ;
    buf_clk cell_17795 ( .C (clk), .D (signal_22682), .Q (signal_22683) ) ;
    buf_clk cell_17803 ( .C (clk), .D (signal_22690), .Q (signal_22691) ) ;
    buf_clk cell_17811 ( .C (clk), .D (signal_22698), .Q (signal_22699) ) ;
    buf_clk cell_17819 ( .C (clk), .D (signal_22706), .Q (signal_22707) ) ;
    buf_clk cell_17827 ( .C (clk), .D (signal_22714), .Q (signal_22715) ) ;
    buf_clk cell_17835 ( .C (clk), .D (signal_22722), .Q (signal_22723) ) ;
    buf_clk cell_17843 ( .C (clk), .D (signal_22730), .Q (signal_22731) ) ;
    buf_clk cell_17851 ( .C (clk), .D (signal_22738), .Q (signal_22739) ) ;
    buf_clk cell_17859 ( .C (clk), .D (signal_22746), .Q (signal_22747) ) ;
    buf_clk cell_17867 ( .C (clk), .D (signal_22754), .Q (signal_22755) ) ;
    buf_clk cell_17875 ( .C (clk), .D (signal_22762), .Q (signal_22763) ) ;
    buf_clk cell_17883 ( .C (clk), .D (signal_22770), .Q (signal_22771) ) ;
    buf_clk cell_17891 ( .C (clk), .D (signal_22778), .Q (signal_22779) ) ;
    buf_clk cell_17899 ( .C (clk), .D (signal_22786), .Q (signal_22787) ) ;
    buf_clk cell_17907 ( .C (clk), .D (signal_22794), .Q (signal_22795) ) ;
    buf_clk cell_17915 ( .C (clk), .D (signal_22802), .Q (signal_22803) ) ;
    buf_clk cell_17923 ( .C (clk), .D (signal_22810), .Q (signal_22811) ) ;
    buf_clk cell_17931 ( .C (clk), .D (signal_22818), .Q (signal_22819) ) ;
    buf_clk cell_17939 ( .C (clk), .D (signal_22826), .Q (signal_22827) ) ;
    buf_clk cell_17947 ( .C (clk), .D (signal_22834), .Q (signal_22835) ) ;
    buf_clk cell_17955 ( .C (clk), .D (signal_22842), .Q (signal_22843) ) ;
    buf_clk cell_17963 ( .C (clk), .D (signal_22850), .Q (signal_22851) ) ;
    buf_clk cell_17971 ( .C (clk), .D (signal_22858), .Q (signal_22859) ) ;
    buf_clk cell_17979 ( .C (clk), .D (signal_22866), .Q (signal_22867) ) ;
    buf_clk cell_17987 ( .C (clk), .D (signal_22874), .Q (signal_22875) ) ;
    buf_clk cell_17995 ( .C (clk), .D (signal_22882), .Q (signal_22883) ) ;
    buf_clk cell_18003 ( .C (clk), .D (signal_22890), .Q (signal_22891) ) ;
    buf_clk cell_18011 ( .C (clk), .D (signal_22898), .Q (signal_22899) ) ;
    buf_clk cell_18019 ( .C (clk), .D (signal_22906), .Q (signal_22907) ) ;
    buf_clk cell_18027 ( .C (clk), .D (signal_22914), .Q (signal_22915) ) ;
    buf_clk cell_18035 ( .C (clk), .D (signal_22922), .Q (signal_22923) ) ;
    buf_clk cell_18043 ( .C (clk), .D (signal_22930), .Q (signal_22931) ) ;
    buf_clk cell_18051 ( .C (clk), .D (signal_22938), .Q (signal_22939) ) ;
    buf_clk cell_18059 ( .C (clk), .D (signal_22946), .Q (signal_22947) ) ;
    buf_clk cell_18067 ( .C (clk), .D (signal_22954), .Q (signal_22955) ) ;
    buf_clk cell_18075 ( .C (clk), .D (signal_22962), .Q (signal_22963) ) ;
    buf_clk cell_18083 ( .C (clk), .D (signal_22970), .Q (signal_22971) ) ;
    buf_clk cell_18091 ( .C (clk), .D (signal_22978), .Q (signal_22979) ) ;
    buf_clk cell_18099 ( .C (clk), .D (signal_22986), .Q (signal_22987) ) ;
    buf_clk cell_18107 ( .C (clk), .D (signal_22994), .Q (signal_22995) ) ;
    buf_clk cell_18115 ( .C (clk), .D (signal_23002), .Q (signal_23003) ) ;
    buf_clk cell_18123 ( .C (clk), .D (signal_23010), .Q (signal_23011) ) ;
    buf_clk cell_18131 ( .C (clk), .D (signal_23018), .Q (signal_23019) ) ;
    buf_clk cell_18139 ( .C (clk), .D (signal_23026), .Q (signal_23027) ) ;
    buf_clk cell_18147 ( .C (clk), .D (signal_23034), .Q (signal_23035) ) ;
    buf_clk cell_18155 ( .C (clk), .D (signal_23042), .Q (signal_23043) ) ;
    buf_clk cell_18163 ( .C (clk), .D (signal_23050), .Q (signal_23051) ) ;
    buf_clk cell_18171 ( .C (clk), .D (signal_23058), .Q (signal_23059) ) ;
    buf_clk cell_18179 ( .C (clk), .D (signal_23066), .Q (signal_23067) ) ;
    buf_clk cell_18187 ( .C (clk), .D (signal_23074), .Q (signal_23075) ) ;
    buf_clk cell_18195 ( .C (clk), .D (signal_23082), .Q (signal_23083) ) ;
    buf_clk cell_18203 ( .C (clk), .D (signal_23090), .Q (signal_23091) ) ;
    buf_clk cell_18211 ( .C (clk), .D (signal_23098), .Q (signal_23099) ) ;
    buf_clk cell_18219 ( .C (clk), .D (signal_23106), .Q (signal_23107) ) ;
    buf_clk cell_18227 ( .C (clk), .D (signal_23114), .Q (signal_23115) ) ;
    buf_clk cell_18235 ( .C (clk), .D (signal_23122), .Q (signal_23123) ) ;
    buf_clk cell_18243 ( .C (clk), .D (signal_23130), .Q (signal_23131) ) ;
    buf_clk cell_18251 ( .C (clk), .D (signal_23138), .Q (signal_23139) ) ;
    buf_clk cell_18259 ( .C (clk), .D (signal_23146), .Q (signal_23147) ) ;
    buf_clk cell_18267 ( .C (clk), .D (signal_23154), .Q (signal_23155) ) ;
    buf_clk cell_18275 ( .C (clk), .D (signal_23162), .Q (signal_23163) ) ;
    buf_clk cell_18283 ( .C (clk), .D (signal_23170), .Q (signal_23171) ) ;
    buf_clk cell_18291 ( .C (clk), .D (signal_23178), .Q (signal_23179) ) ;
    buf_clk cell_18299 ( .C (clk), .D (signal_23186), .Q (signal_23187) ) ;
    buf_clk cell_18307 ( .C (clk), .D (signal_23194), .Q (signal_23195) ) ;
    buf_clk cell_18315 ( .C (clk), .D (signal_23202), .Q (signal_23203) ) ;
    buf_clk cell_18323 ( .C (clk), .D (signal_23210), .Q (signal_23211) ) ;
    buf_clk cell_18331 ( .C (clk), .D (signal_23218), .Q (signal_23219) ) ;
    buf_clk cell_18339 ( .C (clk), .D (signal_23226), .Q (signal_23227) ) ;
    buf_clk cell_18347 ( .C (clk), .D (signal_23234), .Q (signal_23235) ) ;
    buf_clk cell_18355 ( .C (clk), .D (signal_23242), .Q (signal_23243) ) ;
    buf_clk cell_18363 ( .C (clk), .D (signal_23250), .Q (signal_23251) ) ;
    buf_clk cell_18371 ( .C (clk), .D (signal_23258), .Q (signal_23259) ) ;
    buf_clk cell_18379 ( .C (clk), .D (signal_23266), .Q (signal_23267) ) ;
    buf_clk cell_18387 ( .C (clk), .D (signal_23274), .Q (signal_23275) ) ;
    buf_clk cell_18395 ( .C (clk), .D (signal_23282), .Q (signal_23283) ) ;
    buf_clk cell_18407 ( .C (clk), .D (signal_23294), .Q (signal_23295) ) ;
    buf_clk cell_18415 ( .C (clk), .D (signal_23302), .Q (signal_23303) ) ;
    buf_clk cell_18423 ( .C (clk), .D (signal_23310), .Q (signal_23311) ) ;
    buf_clk cell_18431 ( .C (clk), .D (signal_23318), .Q (signal_23319) ) ;
    buf_clk cell_18439 ( .C (clk), .D (signal_23326), .Q (signal_23327) ) ;
    buf_clk cell_18447 ( .C (clk), .D (signal_23334), .Q (signal_23335) ) ;
    buf_clk cell_18455 ( .C (clk), .D (signal_23342), .Q (signal_23343) ) ;
    buf_clk cell_18463 ( .C (clk), .D (signal_23350), .Q (signal_23351) ) ;
    buf_clk cell_18471 ( .C (clk), .D (signal_23358), .Q (signal_23359) ) ;
    buf_clk cell_18479 ( .C (clk), .D (signal_23366), .Q (signal_23367) ) ;
    buf_clk cell_18487 ( .C (clk), .D (signal_23374), .Q (signal_23375) ) ;
    buf_clk cell_18495 ( .C (clk), .D (signal_23382), .Q (signal_23383) ) ;
    buf_clk cell_18503 ( .C (clk), .D (signal_23390), .Q (signal_23391) ) ;
    buf_clk cell_18511 ( .C (clk), .D (signal_23398), .Q (signal_23399) ) ;
    buf_clk cell_18519 ( .C (clk), .D (signal_23406), .Q (signal_23407) ) ;
    buf_clk cell_18527 ( .C (clk), .D (signal_23414), .Q (signal_23415) ) ;
    buf_clk cell_18535 ( .C (clk), .D (signal_23422), .Q (signal_23423) ) ;
    buf_clk cell_18543 ( .C (clk), .D (signal_23430), .Q (signal_23431) ) ;
    buf_clk cell_18551 ( .C (clk), .D (signal_23438), .Q (signal_23439) ) ;
    buf_clk cell_18559 ( .C (clk), .D (signal_23446), .Q (signal_23447) ) ;
    buf_clk cell_18567 ( .C (clk), .D (signal_23454), .Q (signal_23455) ) ;
    buf_clk cell_18575 ( .C (clk), .D (signal_23462), .Q (signal_23463) ) ;
    buf_clk cell_18583 ( .C (clk), .D (signal_23470), .Q (signal_23471) ) ;
    buf_clk cell_18591 ( .C (clk), .D (signal_23478), .Q (signal_23479) ) ;
    buf_clk cell_18599 ( .C (clk), .D (signal_23486), .Q (signal_23487) ) ;
    buf_clk cell_18607 ( .C (clk), .D (signal_23494), .Q (signal_23495) ) ;
    buf_clk cell_18615 ( .C (clk), .D (signal_23502), .Q (signal_23503) ) ;
    buf_clk cell_18623 ( .C (clk), .D (signal_23510), .Q (signal_23511) ) ;
    buf_clk cell_18631 ( .C (clk), .D (signal_23518), .Q (signal_23519) ) ;
    buf_clk cell_18639 ( .C (clk), .D (signal_23526), .Q (signal_23527) ) ;
    buf_clk cell_18651 ( .C (clk), .D (signal_23538), .Q (signal_23539) ) ;
    buf_clk cell_18659 ( .C (clk), .D (signal_23546), .Q (signal_23547) ) ;
    buf_clk cell_18667 ( .C (clk), .D (signal_23554), .Q (signal_23555) ) ;
    buf_clk cell_18675 ( .C (clk), .D (signal_23562), .Q (signal_23563) ) ;
    buf_clk cell_18683 ( .C (clk), .D (signal_23570), .Q (signal_23571) ) ;
    buf_clk cell_18691 ( .C (clk), .D (signal_23578), .Q (signal_23579) ) ;
    buf_clk cell_18699 ( .C (clk), .D (signal_23586), .Q (signal_23587) ) ;
    buf_clk cell_18707 ( .C (clk), .D (signal_23594), .Q (signal_23595) ) ;
    buf_clk cell_18715 ( .C (clk), .D (signal_23602), .Q (signal_23603) ) ;
    buf_clk cell_18723 ( .C (clk), .D (signal_23610), .Q (signal_23611) ) ;
    buf_clk cell_18731 ( .C (clk), .D (signal_23618), .Q (signal_23619) ) ;
    buf_clk cell_18739 ( .C (clk), .D (signal_23626), .Q (signal_23627) ) ;
    buf_clk cell_18751 ( .C (clk), .D (signal_23638), .Q (signal_23639) ) ;
    buf_clk cell_18759 ( .C (clk), .D (signal_23646), .Q (signal_23647) ) ;
    buf_clk cell_18767 ( .C (clk), .D (signal_23654), .Q (signal_23655) ) ;
    buf_clk cell_18775 ( .C (clk), .D (signal_23662), .Q (signal_23663) ) ;
    buf_clk cell_18783 ( .C (clk), .D (signal_23670), .Q (signal_23671) ) ;
    buf_clk cell_18791 ( .C (clk), .D (signal_23678), .Q (signal_23679) ) ;
    buf_clk cell_18799 ( .C (clk), .D (signal_23686), .Q (signal_23687) ) ;
    buf_clk cell_18807 ( .C (clk), .D (signal_23694), .Q (signal_23695) ) ;
    buf_clk cell_18815 ( .C (clk), .D (signal_23702), .Q (signal_23703) ) ;
    buf_clk cell_18823 ( .C (clk), .D (signal_23710), .Q (signal_23711) ) ;
    buf_clk cell_18831 ( .C (clk), .D (signal_23718), .Q (signal_23719) ) ;
    buf_clk cell_18839 ( .C (clk), .D (signal_23726), .Q (signal_23727) ) ;
    buf_clk cell_18847 ( .C (clk), .D (signal_23734), .Q (signal_23735) ) ;
    buf_clk cell_18855 ( .C (clk), .D (signal_23742), .Q (signal_23743) ) ;
    buf_clk cell_18863 ( .C (clk), .D (signal_23750), .Q (signal_23751) ) ;
    buf_clk cell_18871 ( .C (clk), .D (signal_23758), .Q (signal_23759) ) ;
    buf_clk cell_18879 ( .C (clk), .D (signal_23766), .Q (signal_23767) ) ;
    buf_clk cell_18887 ( .C (clk), .D (signal_23774), .Q (signal_23775) ) ;
    buf_clk cell_18895 ( .C (clk), .D (signal_23782), .Q (signal_23783) ) ;
    buf_clk cell_18903 ( .C (clk), .D (signal_23790), .Q (signal_23791) ) ;
    buf_clk cell_18911 ( .C (clk), .D (signal_23798), .Q (signal_23799) ) ;
    buf_clk cell_18919 ( .C (clk), .D (signal_23806), .Q (signal_23807) ) ;
    buf_clk cell_18927 ( .C (clk), .D (signal_23814), .Q (signal_23815) ) ;
    buf_clk cell_18935 ( .C (clk), .D (signal_23822), .Q (signal_23823) ) ;
    buf_clk cell_18943 ( .C (clk), .D (signal_23830), .Q (signal_23831) ) ;
    buf_clk cell_18951 ( .C (clk), .D (signal_23838), .Q (signal_23839) ) ;
    buf_clk cell_18959 ( .C (clk), .D (signal_23846), .Q (signal_23847) ) ;
    buf_clk cell_18967 ( .C (clk), .D (signal_23854), .Q (signal_23855) ) ;
    buf_clk cell_18975 ( .C (clk), .D (signal_23862), .Q (signal_23863) ) ;
    buf_clk cell_18983 ( .C (clk), .D (signal_23870), .Q (signal_23871) ) ;
    buf_clk cell_18991 ( .C (clk), .D (signal_23878), .Q (signal_23879) ) ;
    buf_clk cell_18999 ( .C (clk), .D (signal_23886), .Q (signal_23887) ) ;
    buf_clk cell_19007 ( .C (clk), .D (signal_23894), .Q (signal_23895) ) ;
    buf_clk cell_19015 ( .C (clk), .D (signal_23902), .Q (signal_23903) ) ;
    buf_clk cell_19023 ( .C (clk), .D (signal_23910), .Q (signal_23911) ) ;
    buf_clk cell_19031 ( .C (clk), .D (signal_23918), .Q (signal_23919) ) ;
    buf_clk cell_19039 ( .C (clk), .D (signal_23926), .Q (signal_23927) ) ;
    buf_clk cell_19047 ( .C (clk), .D (signal_23934), .Q (signal_23935) ) ;
    buf_clk cell_19055 ( .C (clk), .D (signal_23942), .Q (signal_23943) ) ;
    buf_clk cell_19063 ( .C (clk), .D (signal_23950), .Q (signal_23951) ) ;
    buf_clk cell_19071 ( .C (clk), .D (signal_23958), .Q (signal_23959) ) ;
    buf_clk cell_19079 ( .C (clk), .D (signal_23966), .Q (signal_23967) ) ;
    buf_clk cell_19087 ( .C (clk), .D (signal_23974), .Q (signal_23975) ) ;
    buf_clk cell_19095 ( .C (clk), .D (signal_23982), .Q (signal_23983) ) ;
    buf_clk cell_19103 ( .C (clk), .D (signal_23990), .Q (signal_23991) ) ;
    buf_clk cell_19111 ( .C (clk), .D (signal_23998), .Q (signal_23999) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5241 ( .a ({signal_8758, signal_5420}), .b ({signal_8760, signal_5422}), .clk (clk), .r (Fresh[180]), .c ({signal_8837, signal_5477}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5242 ( .a ({signal_8759, signal_5421}), .b ({signal_8760, signal_5422}), .clk (clk), .r (Fresh[181]), .c ({signal_8838, signal_5478}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5243 ( .a ({signal_8762, signal_5439}), .b ({signal_8764, signal_5441}), .clk (clk), .r (Fresh[182]), .c ({signal_8839, signal_5479}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5244 ( .a ({signal_8763, signal_5440}), .b ({signal_8764, signal_5441}), .clk (clk), .r (Fresh[183]), .c ({signal_8840, signal_5480}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5245 ( .a ({signal_8766, signal_5458}), .b ({signal_8768, signal_5460}), .clk (clk), .r (Fresh[184]), .c ({signal_8841, signal_5481}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5246 ( .a ({signal_8767, signal_5459}), .b ({signal_8768, signal_5460}), .clk (clk), .r (Fresh[185]), .c ({signal_8842, signal_5482}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5247 ( .a ({signal_8742, signal_5462}), .b ({signal_8744, signal_5464}), .clk (clk), .r (Fresh[186]), .c ({signal_8769, signal_5483}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5248 ( .a ({signal_8743, signal_5463}), .b ({signal_8744, signal_5464}), .clk (clk), .r (Fresh[187]), .c ({signal_8770, signal_5484}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5249 ( .a ({signal_8746, signal_5466}), .b ({signal_8748, signal_5468}), .clk (clk), .r (Fresh[188]), .c ({signal_8771, signal_5485}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5250 ( .a ({signal_8747, signal_5467}), .b ({signal_8748, signal_5468}), .clk (clk), .r (Fresh[189]), .c ({signal_8772, signal_5486}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5251 ( .a ({signal_8750, signal_5470}), .b ({signal_8752, signal_5472}), .clk (clk), .r (Fresh[190]), .c ({signal_8773, signal_5487}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5252 ( .a ({signal_8751, signal_5471}), .b ({signal_8752, signal_5472}), .clk (clk), .r (Fresh[191]), .c ({signal_8774, signal_5488}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5253 ( .a ({signal_8754, signal_5474}), .b ({signal_8756, signal_5476}), .clk (clk), .r (Fresh[192]), .c ({signal_8775, signal_5489}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5254 ( .a ({signal_8755, signal_5475}), .b ({signal_8756, signal_5476}), .clk (clk), .r (Fresh[193]), .c ({signal_8776, signal_5490}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5321 ( .a ({signal_8778, signal_5492}), .b ({signal_8780, signal_5494}), .clk (clk), .r (Fresh[194]), .c ({signal_8849, signal_5557}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5322 ( .a ({signal_8779, signal_5493}), .b ({signal_8780, signal_5494}), .clk (clk), .r (Fresh[195]), .c ({signal_8850, signal_5558}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5323 ( .a ({signal_8782, signal_5496}), .b ({signal_8784, signal_5498}), .clk (clk), .r (Fresh[196]), .c ({signal_8851, signal_5559}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5324 ( .a ({signal_8783, signal_5497}), .b ({signal_8784, signal_5498}), .clk (clk), .r (Fresh[197]), .c ({signal_8852, signal_5560}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5325 ( .a ({signal_8786, signal_5500}), .b ({signal_8788, signal_5502}), .clk (clk), .r (Fresh[198]), .c ({signal_8853, signal_5561}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5326 ( .a ({signal_8787, signal_5501}), .b ({signal_8788, signal_5502}), .clk (clk), .r (Fresh[199]), .c ({signal_8854, signal_5562}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5327 ( .a ({signal_8790, signal_5504}), .b ({signal_8792, signal_5506}), .clk (clk), .r (Fresh[200]), .c ({signal_8855, signal_5563}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5328 ( .a ({signal_8791, signal_5505}), .b ({signal_8792, signal_5506}), .clk (clk), .r (Fresh[201]), .c ({signal_8856, signal_5564}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5329 ( .a ({signal_8794, signal_5508}), .b ({signal_8796, signal_5510}), .clk (clk), .r (Fresh[202]), .c ({signal_8857, signal_5565}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5330 ( .a ({signal_8795, signal_5509}), .b ({signal_8796, signal_5510}), .clk (clk), .r (Fresh[203]), .c ({signal_8858, signal_5566}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5331 ( .a ({signal_8798, signal_5512}), .b ({signal_8800, signal_5514}), .clk (clk), .r (Fresh[204]), .c ({signal_8859, signal_5567}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5332 ( .a ({signal_8799, signal_5513}), .b ({signal_8800, signal_5514}), .clk (clk), .r (Fresh[205]), .c ({signal_8860, signal_5568}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5333 ( .a ({signal_8802, signal_5516}), .b ({signal_8804, signal_5518}), .clk (clk), .r (Fresh[206]), .c ({signal_8861, signal_5569}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5334 ( .a ({signal_8803, signal_5517}), .b ({signal_8804, signal_5518}), .clk (clk), .r (Fresh[207]), .c ({signal_8862, signal_5570}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5335 ( .a ({signal_8758, signal_5420}), .b ({signal_8843, signal_5519}), .clk (clk), .r (Fresh[208]), .c ({signal_8921, signal_5571}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5336 ( .a ({signal_8806, signal_5522}), .b ({signal_8808, signal_5524}), .clk (clk), .r (Fresh[209]), .c ({signal_8863, signal_5572}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5337 ( .a ({signal_8807, signal_5523}), .b ({signal_8808, signal_5524}), .clk (clk), .r (Fresh[210]), .c ({signal_8864, signal_5573}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5338 ( .a ({signal_8810, signal_5526}), .b ({signal_8812, signal_5528}), .clk (clk), .r (Fresh[211]), .c ({signal_8865, signal_5574}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5339 ( .a ({signal_8811, signal_5527}), .b ({signal_8812, signal_5528}), .clk (clk), .r (Fresh[212]), .c ({signal_8866, signal_5575}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5340 ( .a ({signal_8814, signal_5530}), .b ({signal_8816, signal_5532}), .clk (clk), .r (Fresh[213]), .c ({signal_8867, signal_5576}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5341 ( .a ({signal_8815, signal_5531}), .b ({signal_8816, signal_5532}), .clk (clk), .r (Fresh[214]), .c ({signal_8868, signal_5577}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5342 ( .a ({signal_8762, signal_5439}), .b ({signal_8845, signal_5533}), .clk (clk), .r (Fresh[215]), .c ({signal_8922, signal_5578}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5343 ( .a ({signal_8818, signal_5536}), .b ({signal_8820, signal_5538}), .clk (clk), .r (Fresh[216]), .c ({signal_8869, signal_5579}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5344 ( .a ({signal_8819, signal_5537}), .b ({signal_8820, signal_5538}), .clk (clk), .r (Fresh[217]), .c ({signal_8870, signal_5580}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5345 ( .a ({signal_8822, signal_5540}), .b ({signal_8824, signal_5542}), .clk (clk), .r (Fresh[218]), .c ({signal_8871, signal_5581}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5346 ( .a ({signal_8823, signal_5541}), .b ({signal_8824, signal_5542}), .clk (clk), .r (Fresh[219]), .c ({signal_8872, signal_5582}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5347 ( .a ({signal_8826, signal_5544}), .b ({signal_8828, signal_5546}), .clk (clk), .r (Fresh[220]), .c ({signal_8873, signal_5583}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5348 ( .a ({signal_8827, signal_5545}), .b ({signal_8828, signal_5546}), .clk (clk), .r (Fresh[221]), .c ({signal_8874, signal_5584}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5349 ( .a ({signal_8766, signal_5458}), .b ({signal_8847, signal_5547}), .clk (clk), .r (Fresh[222]), .c ({signal_8923, signal_5585}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5350 ( .a ({signal_8742, signal_5462}), .b ({signal_8829, signal_5549}), .clk (clk), .r (Fresh[223]), .c ({signal_8875, signal_5586}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5351 ( .a ({signal_8746, signal_5466}), .b ({signal_8831, signal_5551}), .clk (clk), .r (Fresh[224]), .c ({signal_8876, signal_5587}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5352 ( .a ({signal_8750, signal_5470}), .b ({signal_8833, signal_5553}), .clk (clk), .r (Fresh[225]), .c ({signal_8877, signal_5588}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5353 ( .a ({signal_8754, signal_5474}), .b ({signal_8835, signal_5555}), .clk (clk), .r (Fresh[226]), .c ({signal_8878, signal_5589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5369 ( .a ({signal_12792, signal_12790}), .b ({signal_8837, signal_5477}), .c ({signal_8925, signal_5605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5370 ( .a ({signal_12796, signal_12794}), .b ({signal_8837, signal_5477}), .c ({signal_8926, signal_5606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5371 ( .a ({signal_8837, signal_5477}), .b ({signal_12800, signal_12798}), .c ({signal_8927, signal_5607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5379 ( .a ({signal_12804, signal_12802}), .b ({signal_8839, signal_5479}), .c ({signal_8929, signal_5615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5380 ( .a ({signal_12808, signal_12806}), .b ({signal_8839, signal_5479}), .c ({signal_8930, signal_5616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5381 ( .a ({signal_8839, signal_5479}), .b ({signal_12812, signal_12810}), .c ({signal_8931, signal_5617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5389 ( .a ({signal_12816, signal_12814}), .b ({signal_8841, signal_5481}), .c ({signal_8933, signal_5625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5390 ( .a ({signal_12820, signal_12818}), .b ({signal_8841, signal_5481}), .c ({signal_8934, signal_5626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5391 ( .a ({signal_8841, signal_5481}), .b ({signal_12824, signal_12822}), .c ({signal_8935, signal_5627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5393 ( .a ({signal_12828, signal_12826}), .b ({signal_8769, signal_5483}), .c ({signal_8906, signal_5629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5394 ( .a ({signal_12832, signal_12830}), .b ({signal_8769, signal_5483}), .c ({signal_8907, signal_5630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5395 ( .a ({signal_8769, signal_5483}), .b ({signal_12836, signal_12834}), .c ({signal_8908, signal_5631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5397 ( .a ({signal_12840, signal_12838}), .b ({signal_8771, signal_5485}), .c ({signal_8910, signal_5633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5398 ( .a ({signal_12844, signal_12842}), .b ({signal_8771, signal_5485}), .c ({signal_8911, signal_5634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5399 ( .a ({signal_8771, signal_5485}), .b ({signal_12848, signal_12846}), .c ({signal_8912, signal_5635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5401 ( .a ({signal_12852, signal_12850}), .b ({signal_8773, signal_5487}), .c ({signal_8914, signal_5637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5402 ( .a ({signal_12856, signal_12854}), .b ({signal_8773, signal_5487}), .c ({signal_8915, signal_5638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5403 ( .a ({signal_8773, signal_5487}), .b ({signal_12860, signal_12858}), .c ({signal_8916, signal_5639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5405 ( .a ({signal_12864, signal_12862}), .b ({signal_8775, signal_5489}), .c ({signal_8918, signal_5641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5406 ( .a ({signal_12868, signal_12866}), .b ({signal_8775, signal_5489}), .c ({signal_8919, signal_5642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5407 ( .a ({signal_8775, signal_5489}), .b ({signal_12872, signal_12870}), .c ({signal_8920, signal_5643}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5408 ( .a ({signal_8778, signal_5492}), .b ({signal_8879, signal_5590}), .clk (clk), .r (Fresh[227]), .c ({signal_8936, signal_5644}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5409 ( .a ({signal_8782, signal_5496}), .b ({signal_8881, signal_5592}), .clk (clk), .r (Fresh[228]), .c ({signal_8937, signal_5645}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5410 ( .a ({signal_8786, signal_5500}), .b ({signal_8883, signal_5594}), .clk (clk), .r (Fresh[229]), .c ({signal_8938, signal_5646}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5411 ( .a ({signal_8790, signal_5504}), .b ({signal_8885, signal_5596}), .clk (clk), .r (Fresh[230]), .c ({signal_8939, signal_5647}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5412 ( .a ({signal_8794, signal_5508}), .b ({signal_8887, signal_5598}), .clk (clk), .r (Fresh[231]), .c ({signal_8940, signal_5648}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5413 ( .a ({signal_8798, signal_5512}), .b ({signal_8889, signal_5600}), .clk (clk), .r (Fresh[232]), .c ({signal_8941, signal_5649}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5414 ( .a ({signal_8802, signal_5516}), .b ({signal_8891, signal_5602}), .clk (clk), .r (Fresh[233]), .c ({signal_8942, signal_5650}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5419 ( .a ({signal_8806, signal_5522}), .b ({signal_8893, signal_5608}), .clk (clk), .r (Fresh[234]), .c ({signal_8943, signal_5655}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5420 ( .a ({signal_8810, signal_5526}), .b ({signal_8895, signal_5610}), .clk (clk), .r (Fresh[235]), .c ({signal_8944, signal_5656}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5421 ( .a ({signal_8814, signal_5530}), .b ({signal_8897, signal_5612}), .clk (clk), .r (Fresh[236]), .c ({signal_8945, signal_5657}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5426 ( .a ({signal_8818, signal_5536}), .b ({signal_8899, signal_5618}), .clk (clk), .r (Fresh[237]), .c ({signal_8946, signal_5662}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5427 ( .a ({signal_8822, signal_5540}), .b ({signal_8901, signal_5620}), .clk (clk), .r (Fresh[238]), .c ({signal_8947, signal_5663}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5428 ( .a ({signal_8826, signal_5544}), .b ({signal_8903, signal_5622}), .clk (clk), .r (Fresh[239]), .c ({signal_8948, signal_5664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5450 ( .a ({signal_12876, signal_12874}), .b ({signal_8849, signal_5557}), .c ({signal_8966, signal_5686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5451 ( .a ({signal_12880, signal_12878}), .b ({signal_8849, signal_5557}), .c ({signal_8967, signal_5687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5452 ( .a ({signal_8849, signal_5557}), .b ({signal_12884, signal_12882}), .c ({signal_8968, signal_5688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5454 ( .a ({signal_12888, signal_12886}), .b ({signal_8851, signal_5559}), .c ({signal_8970, signal_5690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5455 ( .a ({signal_12892, signal_12890}), .b ({signal_8851, signal_5559}), .c ({signal_8971, signal_5691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5456 ( .a ({signal_8851, signal_5559}), .b ({signal_12896, signal_12894}), .c ({signal_8972, signal_5692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5458 ( .a ({signal_12900, signal_12898}), .b ({signal_8853, signal_5561}), .c ({signal_8974, signal_5694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5459 ( .a ({signal_12904, signal_12902}), .b ({signal_8853, signal_5561}), .c ({signal_8975, signal_5695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5460 ( .a ({signal_8853, signal_5561}), .b ({signal_12908, signal_12906}), .c ({signal_8976, signal_5696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5462 ( .a ({signal_12912, signal_12910}), .b ({signal_8855, signal_5563}), .c ({signal_8978, signal_5698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5463 ( .a ({signal_12916, signal_12914}), .b ({signal_8855, signal_5563}), .c ({signal_8979, signal_5699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5464 ( .a ({signal_8855, signal_5563}), .b ({signal_12920, signal_12918}), .c ({signal_8980, signal_5700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5466 ( .a ({signal_12924, signal_12922}), .b ({signal_8857, signal_5565}), .c ({signal_8982, signal_5702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5467 ( .a ({signal_12928, signal_12926}), .b ({signal_8857, signal_5565}), .c ({signal_8983, signal_5703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5468 ( .a ({signal_8857, signal_5565}), .b ({signal_12932, signal_12930}), .c ({signal_8984, signal_5704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5470 ( .a ({signal_12936, signal_12934}), .b ({signal_8859, signal_5567}), .c ({signal_8986, signal_5706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5471 ( .a ({signal_12940, signal_12938}), .b ({signal_8859, signal_5567}), .c ({signal_8987, signal_5707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5472 ( .a ({signal_8859, signal_5567}), .b ({signal_12944, signal_12942}), .c ({signal_8988, signal_5708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5474 ( .a ({signal_12948, signal_12946}), .b ({signal_8861, signal_5569}), .c ({signal_8990, signal_5710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5475 ( .a ({signal_12952, signal_12950}), .b ({signal_8861, signal_5569}), .c ({signal_8991, signal_5711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5476 ( .a ({signal_8861, signal_5569}), .b ({signal_12956, signal_12954}), .c ({signal_8992, signal_5712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5477 ( .a ({signal_8837, signal_5477}), .b ({signal_12960, signal_12958}), .c ({signal_9033, signal_5713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5479 ( .a ({signal_12964, signal_12962}), .b ({signal_8863, signal_5572}), .c ({signal_8994, signal_5715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5480 ( .a ({signal_12968, signal_12966}), .b ({signal_8863, signal_5572}), .c ({signal_8995, signal_5716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5481 ( .a ({signal_8863, signal_5572}), .b ({signal_12972, signal_12970}), .c ({signal_8996, signal_5717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5483 ( .a ({signal_12976, signal_12974}), .b ({signal_8865, signal_5574}), .c ({signal_8998, signal_5719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5484 ( .a ({signal_12980, signal_12978}), .b ({signal_8865, signal_5574}), .c ({signal_8999, signal_5720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5485 ( .a ({signal_8865, signal_5574}), .b ({signal_12984, signal_12982}), .c ({signal_9000, signal_5721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5487 ( .a ({signal_12988, signal_12986}), .b ({signal_8867, signal_5576}), .c ({signal_9002, signal_5723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5488 ( .a ({signal_12992, signal_12990}), .b ({signal_8867, signal_5576}), .c ({signal_9003, signal_5724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5489 ( .a ({signal_8867, signal_5576}), .b ({signal_12996, signal_12994}), .c ({signal_9004, signal_5725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5490 ( .a ({signal_8839, signal_5479}), .b ({signal_13000, signal_12998}), .c ({signal_9034, signal_5726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5492 ( .a ({signal_13004, signal_13002}), .b ({signal_8869, signal_5579}), .c ({signal_9006, signal_5728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5493 ( .a ({signal_13008, signal_13006}), .b ({signal_8869, signal_5579}), .c ({signal_9007, signal_5729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5494 ( .a ({signal_8869, signal_5579}), .b ({signal_13012, signal_13010}), .c ({signal_9008, signal_5730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5496 ( .a ({signal_13016, signal_13014}), .b ({signal_8871, signal_5581}), .c ({signal_9010, signal_5732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5497 ( .a ({signal_13020, signal_13018}), .b ({signal_8871, signal_5581}), .c ({signal_9011, signal_5733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5498 ( .a ({signal_8871, signal_5581}), .b ({signal_13024, signal_13022}), .c ({signal_9012, signal_5734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5500 ( .a ({signal_13028, signal_13026}), .b ({signal_8873, signal_5583}), .c ({signal_9014, signal_5736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5501 ( .a ({signal_13032, signal_13030}), .b ({signal_8873, signal_5583}), .c ({signal_9015, signal_5737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5502 ( .a ({signal_8873, signal_5583}), .b ({signal_13036, signal_13034}), .c ({signal_9016, signal_5738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5503 ( .a ({signal_8841, signal_5481}), .b ({signal_13040, signal_13038}), .c ({signal_9035, signal_5739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5504 ( .a ({signal_8769, signal_5483}), .b ({signal_13044, signal_13042}), .c ({signal_9017, signal_5740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5505 ( .a ({signal_8771, signal_5485}), .b ({signal_13048, signal_13046}), .c ({signal_9018, signal_5741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5506 ( .a ({signal_8773, signal_5487}), .b ({signal_13052, signal_13050}), .c ({signal_9019, signal_5742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5507 ( .a ({signal_8775, signal_5489}), .b ({signal_13056, signal_13054}), .c ({signal_9020, signal_5743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5560 ( .a ({signal_8849, signal_5557}), .b ({signal_13060, signal_13058}), .c ({signal_9088, signal_5796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5561 ( .a ({signal_8851, signal_5559}), .b ({signal_13064, signal_13062}), .c ({signal_9089, signal_5797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5562 ( .a ({signal_8853, signal_5561}), .b ({signal_13068, signal_13066}), .c ({signal_9090, signal_5798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5563 ( .a ({signal_8855, signal_5563}), .b ({signal_13072, signal_13070}), .c ({signal_9091, signal_5799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5564 ( .a ({signal_8857, signal_5565}), .b ({signal_13076, signal_13074}), .c ({signal_9092, signal_5800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5565 ( .a ({signal_8859, signal_5567}), .b ({signal_13080, signal_13078}), .c ({signal_9093, signal_5801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5566 ( .a ({signal_8861, signal_5569}), .b ({signal_13084, signal_13082}), .c ({signal_9094, signal_5802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5571 ( .a ({signal_8863, signal_5572}), .b ({signal_13088, signal_13086}), .c ({signal_9095, signal_5807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5572 ( .a ({signal_8865, signal_5574}), .b ({signal_13092, signal_13090}), .c ({signal_9096, signal_5808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5573 ( .a ({signal_8867, signal_5576}), .b ({signal_13096, signal_13094}), .c ({signal_9097, signal_5809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5578 ( .a ({signal_8869, signal_5579}), .b ({signal_13100, signal_13098}), .c ({signal_9098, signal_5814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5579 ( .a ({signal_8871, signal_5581}), .b ({signal_13104, signal_13102}), .c ({signal_9099, signal_5815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5580 ( .a ({signal_8873, signal_5583}), .b ({signal_13108, signal_13106}), .c ({signal_9100, signal_5816}) ) ;
    buf_clk cell_7902 ( .C (clk), .D (signal_12789), .Q (signal_12790) ) ;
    buf_clk cell_7904 ( .C (clk), .D (signal_12791), .Q (signal_12792) ) ;
    buf_clk cell_7906 ( .C (clk), .D (signal_12793), .Q (signal_12794) ) ;
    buf_clk cell_7908 ( .C (clk), .D (signal_12795), .Q (signal_12796) ) ;
    buf_clk cell_7910 ( .C (clk), .D (signal_12797), .Q (signal_12798) ) ;
    buf_clk cell_7912 ( .C (clk), .D (signal_12799), .Q (signal_12800) ) ;
    buf_clk cell_7914 ( .C (clk), .D (signal_12801), .Q (signal_12802) ) ;
    buf_clk cell_7916 ( .C (clk), .D (signal_12803), .Q (signal_12804) ) ;
    buf_clk cell_7918 ( .C (clk), .D (signal_12805), .Q (signal_12806) ) ;
    buf_clk cell_7920 ( .C (clk), .D (signal_12807), .Q (signal_12808) ) ;
    buf_clk cell_7922 ( .C (clk), .D (signal_12809), .Q (signal_12810) ) ;
    buf_clk cell_7924 ( .C (clk), .D (signal_12811), .Q (signal_12812) ) ;
    buf_clk cell_7926 ( .C (clk), .D (signal_12813), .Q (signal_12814) ) ;
    buf_clk cell_7928 ( .C (clk), .D (signal_12815), .Q (signal_12816) ) ;
    buf_clk cell_7930 ( .C (clk), .D (signal_12817), .Q (signal_12818) ) ;
    buf_clk cell_7932 ( .C (clk), .D (signal_12819), .Q (signal_12820) ) ;
    buf_clk cell_7934 ( .C (clk), .D (signal_12821), .Q (signal_12822) ) ;
    buf_clk cell_7936 ( .C (clk), .D (signal_12823), .Q (signal_12824) ) ;
    buf_clk cell_7938 ( .C (clk), .D (signal_12825), .Q (signal_12826) ) ;
    buf_clk cell_7940 ( .C (clk), .D (signal_12827), .Q (signal_12828) ) ;
    buf_clk cell_7942 ( .C (clk), .D (signal_12829), .Q (signal_12830) ) ;
    buf_clk cell_7944 ( .C (clk), .D (signal_12831), .Q (signal_12832) ) ;
    buf_clk cell_7946 ( .C (clk), .D (signal_12833), .Q (signal_12834) ) ;
    buf_clk cell_7948 ( .C (clk), .D (signal_12835), .Q (signal_12836) ) ;
    buf_clk cell_7950 ( .C (clk), .D (signal_12837), .Q (signal_12838) ) ;
    buf_clk cell_7952 ( .C (clk), .D (signal_12839), .Q (signal_12840) ) ;
    buf_clk cell_7954 ( .C (clk), .D (signal_12841), .Q (signal_12842) ) ;
    buf_clk cell_7956 ( .C (clk), .D (signal_12843), .Q (signal_12844) ) ;
    buf_clk cell_7958 ( .C (clk), .D (signal_12845), .Q (signal_12846) ) ;
    buf_clk cell_7960 ( .C (clk), .D (signal_12847), .Q (signal_12848) ) ;
    buf_clk cell_7962 ( .C (clk), .D (signal_12849), .Q (signal_12850) ) ;
    buf_clk cell_7964 ( .C (clk), .D (signal_12851), .Q (signal_12852) ) ;
    buf_clk cell_7966 ( .C (clk), .D (signal_12853), .Q (signal_12854) ) ;
    buf_clk cell_7968 ( .C (clk), .D (signal_12855), .Q (signal_12856) ) ;
    buf_clk cell_7970 ( .C (clk), .D (signal_12857), .Q (signal_12858) ) ;
    buf_clk cell_7972 ( .C (clk), .D (signal_12859), .Q (signal_12860) ) ;
    buf_clk cell_7974 ( .C (clk), .D (signal_12861), .Q (signal_12862) ) ;
    buf_clk cell_7976 ( .C (clk), .D (signal_12863), .Q (signal_12864) ) ;
    buf_clk cell_7978 ( .C (clk), .D (signal_12865), .Q (signal_12866) ) ;
    buf_clk cell_7980 ( .C (clk), .D (signal_12867), .Q (signal_12868) ) ;
    buf_clk cell_7982 ( .C (clk), .D (signal_12869), .Q (signal_12870) ) ;
    buf_clk cell_7984 ( .C (clk), .D (signal_12871), .Q (signal_12872) ) ;
    buf_clk cell_7986 ( .C (clk), .D (signal_12873), .Q (signal_12874) ) ;
    buf_clk cell_7988 ( .C (clk), .D (signal_12875), .Q (signal_12876) ) ;
    buf_clk cell_7990 ( .C (clk), .D (signal_12877), .Q (signal_12878) ) ;
    buf_clk cell_7992 ( .C (clk), .D (signal_12879), .Q (signal_12880) ) ;
    buf_clk cell_7994 ( .C (clk), .D (signal_12881), .Q (signal_12882) ) ;
    buf_clk cell_7996 ( .C (clk), .D (signal_12883), .Q (signal_12884) ) ;
    buf_clk cell_7998 ( .C (clk), .D (signal_12885), .Q (signal_12886) ) ;
    buf_clk cell_8000 ( .C (clk), .D (signal_12887), .Q (signal_12888) ) ;
    buf_clk cell_8002 ( .C (clk), .D (signal_12889), .Q (signal_12890) ) ;
    buf_clk cell_8004 ( .C (clk), .D (signal_12891), .Q (signal_12892) ) ;
    buf_clk cell_8006 ( .C (clk), .D (signal_12893), .Q (signal_12894) ) ;
    buf_clk cell_8008 ( .C (clk), .D (signal_12895), .Q (signal_12896) ) ;
    buf_clk cell_8010 ( .C (clk), .D (signal_12897), .Q (signal_12898) ) ;
    buf_clk cell_8012 ( .C (clk), .D (signal_12899), .Q (signal_12900) ) ;
    buf_clk cell_8014 ( .C (clk), .D (signal_12901), .Q (signal_12902) ) ;
    buf_clk cell_8016 ( .C (clk), .D (signal_12903), .Q (signal_12904) ) ;
    buf_clk cell_8018 ( .C (clk), .D (signal_12905), .Q (signal_12906) ) ;
    buf_clk cell_8020 ( .C (clk), .D (signal_12907), .Q (signal_12908) ) ;
    buf_clk cell_8022 ( .C (clk), .D (signal_12909), .Q (signal_12910) ) ;
    buf_clk cell_8024 ( .C (clk), .D (signal_12911), .Q (signal_12912) ) ;
    buf_clk cell_8026 ( .C (clk), .D (signal_12913), .Q (signal_12914) ) ;
    buf_clk cell_8028 ( .C (clk), .D (signal_12915), .Q (signal_12916) ) ;
    buf_clk cell_8030 ( .C (clk), .D (signal_12917), .Q (signal_12918) ) ;
    buf_clk cell_8032 ( .C (clk), .D (signal_12919), .Q (signal_12920) ) ;
    buf_clk cell_8034 ( .C (clk), .D (signal_12921), .Q (signal_12922) ) ;
    buf_clk cell_8036 ( .C (clk), .D (signal_12923), .Q (signal_12924) ) ;
    buf_clk cell_8038 ( .C (clk), .D (signal_12925), .Q (signal_12926) ) ;
    buf_clk cell_8040 ( .C (clk), .D (signal_12927), .Q (signal_12928) ) ;
    buf_clk cell_8042 ( .C (clk), .D (signal_12929), .Q (signal_12930) ) ;
    buf_clk cell_8044 ( .C (clk), .D (signal_12931), .Q (signal_12932) ) ;
    buf_clk cell_8046 ( .C (clk), .D (signal_12933), .Q (signal_12934) ) ;
    buf_clk cell_8048 ( .C (clk), .D (signal_12935), .Q (signal_12936) ) ;
    buf_clk cell_8050 ( .C (clk), .D (signal_12937), .Q (signal_12938) ) ;
    buf_clk cell_8052 ( .C (clk), .D (signal_12939), .Q (signal_12940) ) ;
    buf_clk cell_8054 ( .C (clk), .D (signal_12941), .Q (signal_12942) ) ;
    buf_clk cell_8056 ( .C (clk), .D (signal_12943), .Q (signal_12944) ) ;
    buf_clk cell_8058 ( .C (clk), .D (signal_12945), .Q (signal_12946) ) ;
    buf_clk cell_8060 ( .C (clk), .D (signal_12947), .Q (signal_12948) ) ;
    buf_clk cell_8062 ( .C (clk), .D (signal_12949), .Q (signal_12950) ) ;
    buf_clk cell_8064 ( .C (clk), .D (signal_12951), .Q (signal_12952) ) ;
    buf_clk cell_8066 ( .C (clk), .D (signal_12953), .Q (signal_12954) ) ;
    buf_clk cell_8068 ( .C (clk), .D (signal_12955), .Q (signal_12956) ) ;
    buf_clk cell_8070 ( .C (clk), .D (signal_12957), .Q (signal_12958) ) ;
    buf_clk cell_8072 ( .C (clk), .D (signal_12959), .Q (signal_12960) ) ;
    buf_clk cell_8074 ( .C (clk), .D (signal_12961), .Q (signal_12962) ) ;
    buf_clk cell_8076 ( .C (clk), .D (signal_12963), .Q (signal_12964) ) ;
    buf_clk cell_8078 ( .C (clk), .D (signal_12965), .Q (signal_12966) ) ;
    buf_clk cell_8080 ( .C (clk), .D (signal_12967), .Q (signal_12968) ) ;
    buf_clk cell_8082 ( .C (clk), .D (signal_12969), .Q (signal_12970) ) ;
    buf_clk cell_8084 ( .C (clk), .D (signal_12971), .Q (signal_12972) ) ;
    buf_clk cell_8086 ( .C (clk), .D (signal_12973), .Q (signal_12974) ) ;
    buf_clk cell_8088 ( .C (clk), .D (signal_12975), .Q (signal_12976) ) ;
    buf_clk cell_8090 ( .C (clk), .D (signal_12977), .Q (signal_12978) ) ;
    buf_clk cell_8092 ( .C (clk), .D (signal_12979), .Q (signal_12980) ) ;
    buf_clk cell_8094 ( .C (clk), .D (signal_12981), .Q (signal_12982) ) ;
    buf_clk cell_8096 ( .C (clk), .D (signal_12983), .Q (signal_12984) ) ;
    buf_clk cell_8098 ( .C (clk), .D (signal_12985), .Q (signal_12986) ) ;
    buf_clk cell_8100 ( .C (clk), .D (signal_12987), .Q (signal_12988) ) ;
    buf_clk cell_8102 ( .C (clk), .D (signal_12989), .Q (signal_12990) ) ;
    buf_clk cell_8104 ( .C (clk), .D (signal_12991), .Q (signal_12992) ) ;
    buf_clk cell_8106 ( .C (clk), .D (signal_12993), .Q (signal_12994) ) ;
    buf_clk cell_8108 ( .C (clk), .D (signal_12995), .Q (signal_12996) ) ;
    buf_clk cell_8110 ( .C (clk), .D (signal_12997), .Q (signal_12998) ) ;
    buf_clk cell_8112 ( .C (clk), .D (signal_12999), .Q (signal_13000) ) ;
    buf_clk cell_8114 ( .C (clk), .D (signal_13001), .Q (signal_13002) ) ;
    buf_clk cell_8116 ( .C (clk), .D (signal_13003), .Q (signal_13004) ) ;
    buf_clk cell_8118 ( .C (clk), .D (signal_13005), .Q (signal_13006) ) ;
    buf_clk cell_8120 ( .C (clk), .D (signal_13007), .Q (signal_13008) ) ;
    buf_clk cell_8122 ( .C (clk), .D (signal_13009), .Q (signal_13010) ) ;
    buf_clk cell_8124 ( .C (clk), .D (signal_13011), .Q (signal_13012) ) ;
    buf_clk cell_8126 ( .C (clk), .D (signal_13013), .Q (signal_13014) ) ;
    buf_clk cell_8128 ( .C (clk), .D (signal_13015), .Q (signal_13016) ) ;
    buf_clk cell_8130 ( .C (clk), .D (signal_13017), .Q (signal_13018) ) ;
    buf_clk cell_8132 ( .C (clk), .D (signal_13019), .Q (signal_13020) ) ;
    buf_clk cell_8134 ( .C (clk), .D (signal_13021), .Q (signal_13022) ) ;
    buf_clk cell_8136 ( .C (clk), .D (signal_13023), .Q (signal_13024) ) ;
    buf_clk cell_8138 ( .C (clk), .D (signal_13025), .Q (signal_13026) ) ;
    buf_clk cell_8140 ( .C (clk), .D (signal_13027), .Q (signal_13028) ) ;
    buf_clk cell_8142 ( .C (clk), .D (signal_13029), .Q (signal_13030) ) ;
    buf_clk cell_8144 ( .C (clk), .D (signal_13031), .Q (signal_13032) ) ;
    buf_clk cell_8146 ( .C (clk), .D (signal_13033), .Q (signal_13034) ) ;
    buf_clk cell_8148 ( .C (clk), .D (signal_13035), .Q (signal_13036) ) ;
    buf_clk cell_8150 ( .C (clk), .D (signal_13037), .Q (signal_13038) ) ;
    buf_clk cell_8152 ( .C (clk), .D (signal_13039), .Q (signal_13040) ) ;
    buf_clk cell_8154 ( .C (clk), .D (signal_13041), .Q (signal_13042) ) ;
    buf_clk cell_8156 ( .C (clk), .D (signal_13043), .Q (signal_13044) ) ;
    buf_clk cell_8158 ( .C (clk), .D (signal_13045), .Q (signal_13046) ) ;
    buf_clk cell_8160 ( .C (clk), .D (signal_13047), .Q (signal_13048) ) ;
    buf_clk cell_8162 ( .C (clk), .D (signal_13049), .Q (signal_13050) ) ;
    buf_clk cell_8164 ( .C (clk), .D (signal_13051), .Q (signal_13052) ) ;
    buf_clk cell_8166 ( .C (clk), .D (signal_13053), .Q (signal_13054) ) ;
    buf_clk cell_8168 ( .C (clk), .D (signal_13055), .Q (signal_13056) ) ;
    buf_clk cell_8170 ( .C (clk), .D (signal_13057), .Q (signal_13058) ) ;
    buf_clk cell_8172 ( .C (clk), .D (signal_13059), .Q (signal_13060) ) ;
    buf_clk cell_8174 ( .C (clk), .D (signal_13061), .Q (signal_13062) ) ;
    buf_clk cell_8176 ( .C (clk), .D (signal_13063), .Q (signal_13064) ) ;
    buf_clk cell_8178 ( .C (clk), .D (signal_13065), .Q (signal_13066) ) ;
    buf_clk cell_8180 ( .C (clk), .D (signal_13067), .Q (signal_13068) ) ;
    buf_clk cell_8182 ( .C (clk), .D (signal_13069), .Q (signal_13070) ) ;
    buf_clk cell_8184 ( .C (clk), .D (signal_13071), .Q (signal_13072) ) ;
    buf_clk cell_8186 ( .C (clk), .D (signal_13073), .Q (signal_13074) ) ;
    buf_clk cell_8188 ( .C (clk), .D (signal_13075), .Q (signal_13076) ) ;
    buf_clk cell_8190 ( .C (clk), .D (signal_13077), .Q (signal_13078) ) ;
    buf_clk cell_8192 ( .C (clk), .D (signal_13079), .Q (signal_13080) ) ;
    buf_clk cell_8194 ( .C (clk), .D (signal_13081), .Q (signal_13082) ) ;
    buf_clk cell_8196 ( .C (clk), .D (signal_13083), .Q (signal_13084) ) ;
    buf_clk cell_8198 ( .C (clk), .D (signal_13085), .Q (signal_13086) ) ;
    buf_clk cell_8200 ( .C (clk), .D (signal_13087), .Q (signal_13088) ) ;
    buf_clk cell_8202 ( .C (clk), .D (signal_13089), .Q (signal_13090) ) ;
    buf_clk cell_8204 ( .C (clk), .D (signal_13091), .Q (signal_13092) ) ;
    buf_clk cell_8206 ( .C (clk), .D (signal_13093), .Q (signal_13094) ) ;
    buf_clk cell_8208 ( .C (clk), .D (signal_13095), .Q (signal_13096) ) ;
    buf_clk cell_8210 ( .C (clk), .D (signal_13097), .Q (signal_13098) ) ;
    buf_clk cell_8212 ( .C (clk), .D (signal_13099), .Q (signal_13100) ) ;
    buf_clk cell_8214 ( .C (clk), .D (signal_13101), .Q (signal_13102) ) ;
    buf_clk cell_8216 ( .C (clk), .D (signal_13103), .Q (signal_13104) ) ;
    buf_clk cell_8218 ( .C (clk), .D (signal_13105), .Q (signal_13106) ) ;
    buf_clk cell_8220 ( .C (clk), .D (signal_13107), .Q (signal_13108) ) ;
    buf_clk cell_8544 ( .C (clk), .D (signal_13431), .Q (signal_13432) ) ;
    buf_clk cell_8552 ( .C (clk), .D (signal_13439), .Q (signal_13440) ) ;
    buf_clk cell_8560 ( .C (clk), .D (signal_13447), .Q (signal_13448) ) ;
    buf_clk cell_8568 ( .C (clk), .D (signal_13455), .Q (signal_13456) ) ;
    buf_clk cell_8576 ( .C (clk), .D (signal_13463), .Q (signal_13464) ) ;
    buf_clk cell_8584 ( .C (clk), .D (signal_13471), .Q (signal_13472) ) ;
    buf_clk cell_8592 ( .C (clk), .D (signal_13479), .Q (signal_13480) ) ;
    buf_clk cell_8600 ( .C (clk), .D (signal_13487), .Q (signal_13488) ) ;
    buf_clk cell_8608 ( .C (clk), .D (signal_13495), .Q (signal_13496) ) ;
    buf_clk cell_8616 ( .C (clk), .D (signal_13503), .Q (signal_13504) ) ;
    buf_clk cell_8624 ( .C (clk), .D (signal_13511), .Q (signal_13512) ) ;
    buf_clk cell_8632 ( .C (clk), .D (signal_13519), .Q (signal_13520) ) ;
    buf_clk cell_8640 ( .C (clk), .D (signal_13527), .Q (signal_13528) ) ;
    buf_clk cell_8648 ( .C (clk), .D (signal_13535), .Q (signal_13536) ) ;
    buf_clk cell_8656 ( .C (clk), .D (signal_13543), .Q (signal_13544) ) ;
    buf_clk cell_8664 ( .C (clk), .D (signal_13551), .Q (signal_13552) ) ;
    buf_clk cell_8672 ( .C (clk), .D (signal_13559), .Q (signal_13560) ) ;
    buf_clk cell_8680 ( .C (clk), .D (signal_13567), .Q (signal_13568) ) ;
    buf_clk cell_8688 ( .C (clk), .D (signal_13575), .Q (signal_13576) ) ;
    buf_clk cell_8696 ( .C (clk), .D (signal_13583), .Q (signal_13584) ) ;
    buf_clk cell_8704 ( .C (clk), .D (signal_13591), .Q (signal_13592) ) ;
    buf_clk cell_8712 ( .C (clk), .D (signal_13599), .Q (signal_13600) ) ;
    buf_clk cell_8720 ( .C (clk), .D (signal_13607), .Q (signal_13608) ) ;
    buf_clk cell_8728 ( .C (clk), .D (signal_13615), .Q (signal_13616) ) ;
    buf_clk cell_8736 ( .C (clk), .D (signal_13623), .Q (signal_13624) ) ;
    buf_clk cell_8744 ( .C (clk), .D (signal_13631), .Q (signal_13632) ) ;
    buf_clk cell_8752 ( .C (clk), .D (signal_13639), .Q (signal_13640) ) ;
    buf_clk cell_8760 ( .C (clk), .D (signal_13647), .Q (signal_13648) ) ;
    buf_clk cell_8768 ( .C (clk), .D (signal_13655), .Q (signal_13656) ) ;
    buf_clk cell_8776 ( .C (clk), .D (signal_13663), .Q (signal_13664) ) ;
    buf_clk cell_8784 ( .C (clk), .D (signal_13671), .Q (signal_13672) ) ;
    buf_clk cell_8792 ( .C (clk), .D (signal_13679), .Q (signal_13680) ) ;
    buf_clk cell_8800 ( .C (clk), .D (signal_13687), .Q (signal_13688) ) ;
    buf_clk cell_8808 ( .C (clk), .D (signal_13695), .Q (signal_13696) ) ;
    buf_clk cell_8816 ( .C (clk), .D (signal_13703), .Q (signal_13704) ) ;
    buf_clk cell_8824 ( .C (clk), .D (signal_13711), .Q (signal_13712) ) ;
    buf_clk cell_8832 ( .C (clk), .D (signal_13719), .Q (signal_13720) ) ;
    buf_clk cell_8840 ( .C (clk), .D (signal_13727), .Q (signal_13728) ) ;
    buf_clk cell_8848 ( .C (clk), .D (signal_13735), .Q (signal_13736) ) ;
    buf_clk cell_8856 ( .C (clk), .D (signal_13743), .Q (signal_13744) ) ;
    buf_clk cell_8864 ( .C (clk), .D (signal_13751), .Q (signal_13752) ) ;
    buf_clk cell_8872 ( .C (clk), .D (signal_13759), .Q (signal_13760) ) ;
    buf_clk cell_8880 ( .C (clk), .D (signal_13767), .Q (signal_13768) ) ;
    buf_clk cell_8888 ( .C (clk), .D (signal_13775), .Q (signal_13776) ) ;
    buf_clk cell_8896 ( .C (clk), .D (signal_13783), .Q (signal_13784) ) ;
    buf_clk cell_8904 ( .C (clk), .D (signal_13791), .Q (signal_13792) ) ;
    buf_clk cell_8912 ( .C (clk), .D (signal_13799), .Q (signal_13800) ) ;
    buf_clk cell_8920 ( .C (clk), .D (signal_13807), .Q (signal_13808) ) ;
    buf_clk cell_8928 ( .C (clk), .D (signal_13815), .Q (signal_13816) ) ;
    buf_clk cell_8936 ( .C (clk), .D (signal_13823), .Q (signal_13824) ) ;
    buf_clk cell_8944 ( .C (clk), .D (signal_13831), .Q (signal_13832) ) ;
    buf_clk cell_8952 ( .C (clk), .D (signal_13839), .Q (signal_13840) ) ;
    buf_clk cell_8960 ( .C (clk), .D (signal_13847), .Q (signal_13848) ) ;
    buf_clk cell_8968 ( .C (clk), .D (signal_13855), .Q (signal_13856) ) ;
    buf_clk cell_8976 ( .C (clk), .D (signal_13863), .Q (signal_13864) ) ;
    buf_clk cell_8984 ( .C (clk), .D (signal_13871), .Q (signal_13872) ) ;
    buf_clk cell_8992 ( .C (clk), .D (signal_13879), .Q (signal_13880) ) ;
    buf_clk cell_9000 ( .C (clk), .D (signal_13887), .Q (signal_13888) ) ;
    buf_clk cell_9008 ( .C (clk), .D (signal_13895), .Q (signal_13896) ) ;
    buf_clk cell_9016 ( .C (clk), .D (signal_13903), .Q (signal_13904) ) ;
    buf_clk cell_9024 ( .C (clk), .D (signal_13911), .Q (signal_13912) ) ;
    buf_clk cell_9032 ( .C (clk), .D (signal_13919), .Q (signal_13920) ) ;
    buf_clk cell_9040 ( .C (clk), .D (signal_13927), .Q (signal_13928) ) ;
    buf_clk cell_9048 ( .C (clk), .D (signal_13935), .Q (signal_13936) ) ;
    buf_clk cell_9056 ( .C (clk), .D (signal_13943), .Q (signal_13944) ) ;
    buf_clk cell_9064 ( .C (clk), .D (signal_13951), .Q (signal_13952) ) ;
    buf_clk cell_9072 ( .C (clk), .D (signal_13959), .Q (signal_13960) ) ;
    buf_clk cell_9080 ( .C (clk), .D (signal_13967), .Q (signal_13968) ) ;
    buf_clk cell_9088 ( .C (clk), .D (signal_13975), .Q (signal_13976) ) ;
    buf_clk cell_9096 ( .C (clk), .D (signal_13983), .Q (signal_13984) ) ;
    buf_clk cell_9104 ( .C (clk), .D (signal_13991), .Q (signal_13992) ) ;
    buf_clk cell_9112 ( .C (clk), .D (signal_13999), .Q (signal_14000) ) ;
    buf_clk cell_9120 ( .C (clk), .D (signal_14007), .Q (signal_14008) ) ;
    buf_clk cell_9128 ( .C (clk), .D (signal_14015), .Q (signal_14016) ) ;
    buf_clk cell_9136 ( .C (clk), .D (signal_14023), .Q (signal_14024) ) ;
    buf_clk cell_9144 ( .C (clk), .D (signal_14031), .Q (signal_14032) ) ;
    buf_clk cell_9152 ( .C (clk), .D (signal_14039), .Q (signal_14040) ) ;
    buf_clk cell_9160 ( .C (clk), .D (signal_14047), .Q (signal_14048) ) ;
    buf_clk cell_9168 ( .C (clk), .D (signal_14055), .Q (signal_14056) ) ;
    buf_clk cell_9176 ( .C (clk), .D (signal_14063), .Q (signal_14064) ) ;
    buf_clk cell_9184 ( .C (clk), .D (signal_14071), .Q (signal_14072) ) ;
    buf_clk cell_9192 ( .C (clk), .D (signal_14079), .Q (signal_14080) ) ;
    buf_clk cell_9200 ( .C (clk), .D (signal_14087), .Q (signal_14088) ) ;
    buf_clk cell_9208 ( .C (clk), .D (signal_14095), .Q (signal_14096) ) ;
    buf_clk cell_9216 ( .C (clk), .D (signal_14103), .Q (signal_14104) ) ;
    buf_clk cell_9224 ( .C (clk), .D (signal_14111), .Q (signal_14112) ) ;
    buf_clk cell_9232 ( .C (clk), .D (signal_14119), .Q (signal_14120) ) ;
    buf_clk cell_9240 ( .C (clk), .D (signal_14127), .Q (signal_14128) ) ;
    buf_clk cell_9248 ( .C (clk), .D (signal_14135), .Q (signal_14136) ) ;
    buf_clk cell_9256 ( .C (clk), .D (signal_14143), .Q (signal_14144) ) ;
    buf_clk cell_9264 ( .C (clk), .D (signal_14151), .Q (signal_14152) ) ;
    buf_clk cell_9272 ( .C (clk), .D (signal_14159), .Q (signal_14160) ) ;
    buf_clk cell_9280 ( .C (clk), .D (signal_14167), .Q (signal_14168) ) ;
    buf_clk cell_9288 ( .C (clk), .D (signal_14175), .Q (signal_14176) ) ;
    buf_clk cell_9296 ( .C (clk), .D (signal_14183), .Q (signal_14184) ) ;
    buf_clk cell_9304 ( .C (clk), .D (signal_14191), .Q (signal_14192) ) ;
    buf_clk cell_9312 ( .C (clk), .D (signal_14199), .Q (signal_14200) ) ;
    buf_clk cell_9320 ( .C (clk), .D (signal_14207), .Q (signal_14208) ) ;
    buf_clk cell_9328 ( .C (clk), .D (signal_14215), .Q (signal_14216) ) ;
    buf_clk cell_9336 ( .C (clk), .D (signal_14223), .Q (signal_14224) ) ;
    buf_clk cell_9344 ( .C (clk), .D (signal_14231), .Q (signal_14232) ) ;
    buf_clk cell_9352 ( .C (clk), .D (signal_14239), .Q (signal_14240) ) ;
    buf_clk cell_9360 ( .C (clk), .D (signal_14247), .Q (signal_14248) ) ;
    buf_clk cell_9368 ( .C (clk), .D (signal_14255), .Q (signal_14256) ) ;
    buf_clk cell_9376 ( .C (clk), .D (signal_14263), .Q (signal_14264) ) ;
    buf_clk cell_9384 ( .C (clk), .D (signal_14271), .Q (signal_14272) ) ;
    buf_clk cell_9392 ( .C (clk), .D (signal_14279), .Q (signal_14280) ) ;
    buf_clk cell_9400 ( .C (clk), .D (signal_14287), .Q (signal_14288) ) ;
    buf_clk cell_9408 ( .C (clk), .D (signal_14295), .Q (signal_14296) ) ;
    buf_clk cell_9416 ( .C (clk), .D (signal_14303), .Q (signal_14304) ) ;
    buf_clk cell_9424 ( .C (clk), .D (signal_14311), .Q (signal_14312) ) ;
    buf_clk cell_9432 ( .C (clk), .D (signal_14319), .Q (signal_14320) ) ;
    buf_clk cell_9440 ( .C (clk), .D (signal_14327), .Q (signal_14328) ) ;
    buf_clk cell_9448 ( .C (clk), .D (signal_14335), .Q (signal_14336) ) ;
    buf_clk cell_9456 ( .C (clk), .D (signal_14343), .Q (signal_14344) ) ;
    buf_clk cell_9464 ( .C (clk), .D (signal_14351), .Q (signal_14352) ) ;
    buf_clk cell_9472 ( .C (clk), .D (signal_14359), .Q (signal_14360) ) ;
    buf_clk cell_9480 ( .C (clk), .D (signal_14367), .Q (signal_14368) ) ;
    buf_clk cell_9488 ( .C (clk), .D (signal_14375), .Q (signal_14376) ) ;
    buf_clk cell_9496 ( .C (clk), .D (signal_14383), .Q (signal_14384) ) ;
    buf_clk cell_9504 ( .C (clk), .D (signal_14391), .Q (signal_14392) ) ;
    buf_clk cell_9512 ( .C (clk), .D (signal_14399), .Q (signal_14400) ) ;
    buf_clk cell_9520 ( .C (clk), .D (signal_14407), .Q (signal_14408) ) ;
    buf_clk cell_9528 ( .C (clk), .D (signal_14415), .Q (signal_14416) ) ;
    buf_clk cell_9536 ( .C (clk), .D (signal_14423), .Q (signal_14424) ) ;
    buf_clk cell_9544 ( .C (clk), .D (signal_14431), .Q (signal_14432) ) ;
    buf_clk cell_9552 ( .C (clk), .D (signal_14439), .Q (signal_14440) ) ;
    buf_clk cell_9560 ( .C (clk), .D (signal_14447), .Q (signal_14448) ) ;
    buf_clk cell_9568 ( .C (clk), .D (signal_14455), .Q (signal_14456) ) ;
    buf_clk cell_9576 ( .C (clk), .D (signal_14463), .Q (signal_14464) ) ;
    buf_clk cell_9584 ( .C (clk), .D (signal_14471), .Q (signal_14472) ) ;
    buf_clk cell_9592 ( .C (clk), .D (signal_14479), .Q (signal_14480) ) ;
    buf_clk cell_9600 ( .C (clk), .D (signal_14487), .Q (signal_14488) ) ;
    buf_clk cell_9608 ( .C (clk), .D (signal_14495), .Q (signal_14496) ) ;
    buf_clk cell_9616 ( .C (clk), .D (signal_14503), .Q (signal_14504) ) ;
    buf_clk cell_9624 ( .C (clk), .D (signal_14511), .Q (signal_14512) ) ;
    buf_clk cell_9632 ( .C (clk), .D (signal_14519), .Q (signal_14520) ) ;
    buf_clk cell_9640 ( .C (clk), .D (signal_14527), .Q (signal_14528) ) ;
    buf_clk cell_9648 ( .C (clk), .D (signal_14535), .Q (signal_14536) ) ;
    buf_clk cell_9656 ( .C (clk), .D (signal_14543), .Q (signal_14544) ) ;
    buf_clk cell_9664 ( .C (clk), .D (signal_14551), .Q (signal_14552) ) ;
    buf_clk cell_9672 ( .C (clk), .D (signal_14559), .Q (signal_14560) ) ;
    buf_clk cell_9680 ( .C (clk), .D (signal_14567), .Q (signal_14568) ) ;
    buf_clk cell_9688 ( .C (clk), .D (signal_14575), .Q (signal_14576) ) ;
    buf_clk cell_9696 ( .C (clk), .D (signal_14583), .Q (signal_14584) ) ;
    buf_clk cell_9704 ( .C (clk), .D (signal_14591), .Q (signal_14592) ) ;
    buf_clk cell_9712 ( .C (clk), .D (signal_14599), .Q (signal_14600) ) ;
    buf_clk cell_9720 ( .C (clk), .D (signal_14607), .Q (signal_14608) ) ;
    buf_clk cell_9728 ( .C (clk), .D (signal_14615), .Q (signal_14616) ) ;
    buf_clk cell_9736 ( .C (clk), .D (signal_14623), .Q (signal_14624) ) ;
    buf_clk cell_9744 ( .C (clk), .D (signal_14631), .Q (signal_14632) ) ;
    buf_clk cell_9752 ( .C (clk), .D (signal_14639), .Q (signal_14640) ) ;
    buf_clk cell_9760 ( .C (clk), .D (signal_14647), .Q (signal_14648) ) ;
    buf_clk cell_9768 ( .C (clk), .D (signal_14655), .Q (signal_14656) ) ;
    buf_clk cell_9776 ( .C (clk), .D (signal_14663), .Q (signal_14664) ) ;
    buf_clk cell_9784 ( .C (clk), .D (signal_14671), .Q (signal_14672) ) ;
    buf_clk cell_9792 ( .C (clk), .D (signal_14679), .Q (signal_14680) ) ;
    buf_clk cell_9800 ( .C (clk), .D (signal_14687), .Q (signal_14688) ) ;
    buf_clk cell_9808 ( .C (clk), .D (signal_14695), .Q (signal_14696) ) ;
    buf_clk cell_9816 ( .C (clk), .D (signal_14703), .Q (signal_14704) ) ;
    buf_clk cell_9824 ( .C (clk), .D (signal_14711), .Q (signal_14712) ) ;
    buf_clk cell_9832 ( .C (clk), .D (signal_14719), .Q (signal_14720) ) ;
    buf_clk cell_9840 ( .C (clk), .D (signal_14727), .Q (signal_14728) ) ;
    buf_clk cell_9848 ( .C (clk), .D (signal_14735), .Q (signal_14736) ) ;
    buf_clk cell_9856 ( .C (clk), .D (signal_14743), .Q (signal_14744) ) ;
    buf_clk cell_9864 ( .C (clk), .D (signal_14751), .Q (signal_14752) ) ;
    buf_clk cell_9872 ( .C (clk), .D (signal_14759), .Q (signal_14760) ) ;
    buf_clk cell_9880 ( .C (clk), .D (signal_14767), .Q (signal_14768) ) ;
    buf_clk cell_9888 ( .C (clk), .D (signal_14775), .Q (signal_14776) ) ;
    buf_clk cell_9896 ( .C (clk), .D (signal_14783), .Q (signal_14784) ) ;
    buf_clk cell_9904 ( .C (clk), .D (signal_14791), .Q (signal_14792) ) ;
    buf_clk cell_9912 ( .C (clk), .D (signal_14799), .Q (signal_14800) ) ;
    buf_clk cell_9920 ( .C (clk), .D (signal_14807), .Q (signal_14808) ) ;
    buf_clk cell_9928 ( .C (clk), .D (signal_14815), .Q (signal_14816) ) ;
    buf_clk cell_9936 ( .C (clk), .D (signal_14823), .Q (signal_14824) ) ;
    buf_clk cell_9944 ( .C (clk), .D (signal_14831), .Q (signal_14832) ) ;
    buf_clk cell_9952 ( .C (clk), .D (signal_14839), .Q (signal_14840) ) ;
    buf_clk cell_9960 ( .C (clk), .D (signal_14847), .Q (signal_14848) ) ;
    buf_clk cell_9968 ( .C (clk), .D (signal_14855), .Q (signal_14856) ) ;
    buf_clk cell_9976 ( .C (clk), .D (signal_14863), .Q (signal_14864) ) ;
    buf_clk cell_9984 ( .C (clk), .D (signal_14871), .Q (signal_14872) ) ;
    buf_clk cell_9992 ( .C (clk), .D (signal_14879), .Q (signal_14880) ) ;
    buf_clk cell_10000 ( .C (clk), .D (signal_14887), .Q (signal_14888) ) ;
    buf_clk cell_10008 ( .C (clk), .D (signal_14895), .Q (signal_14896) ) ;
    buf_clk cell_10016 ( .C (clk), .D (signal_14903), .Q (signal_14904) ) ;
    buf_clk cell_10024 ( .C (clk), .D (signal_14911), .Q (signal_14912) ) ;
    buf_clk cell_10032 ( .C (clk), .D (signal_14919), .Q (signal_14920) ) ;
    buf_clk cell_10040 ( .C (clk), .D (signal_14927), .Q (signal_14928) ) ;
    buf_clk cell_10048 ( .C (clk), .D (signal_14935), .Q (signal_14936) ) ;
    buf_clk cell_10056 ( .C (clk), .D (signal_14943), .Q (signal_14944) ) ;
    buf_clk cell_10064 ( .C (clk), .D (signal_14951), .Q (signal_14952) ) ;
    buf_clk cell_10072 ( .C (clk), .D (signal_14959), .Q (signal_14960) ) ;
    buf_clk cell_10080 ( .C (clk), .D (signal_14967), .Q (signal_14968) ) ;
    buf_clk cell_10088 ( .C (clk), .D (signal_14975), .Q (signal_14976) ) ;
    buf_clk cell_10096 ( .C (clk), .D (signal_14983), .Q (signal_14984) ) ;
    buf_clk cell_10104 ( .C (clk), .D (signal_14991), .Q (signal_14992) ) ;
    buf_clk cell_10112 ( .C (clk), .D (signal_14999), .Q (signal_15000) ) ;
    buf_clk cell_10120 ( .C (clk), .D (signal_15007), .Q (signal_15008) ) ;
    buf_clk cell_10128 ( .C (clk), .D (signal_15015), .Q (signal_15016) ) ;
    buf_clk cell_10136 ( .C (clk), .D (signal_15023), .Q (signal_15024) ) ;
    buf_clk cell_10144 ( .C (clk), .D (signal_15031), .Q (signal_15032) ) ;
    buf_clk cell_10152 ( .C (clk), .D (signal_15039), .Q (signal_15040) ) ;
    buf_clk cell_10160 ( .C (clk), .D (signal_15047), .Q (signal_15048) ) ;
    buf_clk cell_10168 ( .C (clk), .D (signal_15055), .Q (signal_15056) ) ;
    buf_clk cell_10176 ( .C (clk), .D (signal_15063), .Q (signal_15064) ) ;
    buf_clk cell_10184 ( .C (clk), .D (signal_15071), .Q (signal_15072) ) ;
    buf_clk cell_10192 ( .C (clk), .D (signal_15079), .Q (signal_15080) ) ;
    buf_clk cell_10200 ( .C (clk), .D (signal_15087), .Q (signal_15088) ) ;
    buf_clk cell_10208 ( .C (clk), .D (signal_15095), .Q (signal_15096) ) ;
    buf_clk cell_10216 ( .C (clk), .D (signal_15103), .Q (signal_15104) ) ;
    buf_clk cell_10224 ( .C (clk), .D (signal_15111), .Q (signal_15112) ) ;
    buf_clk cell_10232 ( .C (clk), .D (signal_15119), .Q (signal_15120) ) ;
    buf_clk cell_10240 ( .C (clk), .D (signal_15127), .Q (signal_15128) ) ;
    buf_clk cell_10248 ( .C (clk), .D (signal_15135), .Q (signal_15136) ) ;
    buf_clk cell_10256 ( .C (clk), .D (signal_15143), .Q (signal_15144) ) ;
    buf_clk cell_10264 ( .C (clk), .D (signal_15151), .Q (signal_15152) ) ;
    buf_clk cell_10272 ( .C (clk), .D (signal_15159), .Q (signal_15160) ) ;
    buf_clk cell_10280 ( .C (clk), .D (signal_15167), .Q (signal_15168) ) ;
    buf_clk cell_10288 ( .C (clk), .D (signal_15175), .Q (signal_15176) ) ;
    buf_clk cell_10296 ( .C (clk), .D (signal_15183), .Q (signal_15184) ) ;
    buf_clk cell_10304 ( .C (clk), .D (signal_15191), .Q (signal_15192) ) ;
    buf_clk cell_10312 ( .C (clk), .D (signal_15199), .Q (signal_15200) ) ;
    buf_clk cell_10320 ( .C (clk), .D (signal_15207), .Q (signal_15208) ) ;
    buf_clk cell_10328 ( .C (clk), .D (signal_15215), .Q (signal_15216) ) ;
    buf_clk cell_10336 ( .C (clk), .D (signal_15223), .Q (signal_15224) ) ;
    buf_clk cell_10344 ( .C (clk), .D (signal_15231), .Q (signal_15232) ) ;
    buf_clk cell_10352 ( .C (clk), .D (signal_15239), .Q (signal_15240) ) ;
    buf_clk cell_10360 ( .C (clk), .D (signal_15247), .Q (signal_15248) ) ;
    buf_clk cell_10368 ( .C (clk), .D (signal_15255), .Q (signal_15256) ) ;
    buf_clk cell_10376 ( .C (clk), .D (signal_15263), .Q (signal_15264) ) ;
    buf_clk cell_10384 ( .C (clk), .D (signal_15271), .Q (signal_15272) ) ;
    buf_clk cell_10392 ( .C (clk), .D (signal_15279), .Q (signal_15280) ) ;
    buf_clk cell_10400 ( .C (clk), .D (signal_15287), .Q (signal_15288) ) ;
    buf_clk cell_10408 ( .C (clk), .D (signal_15295), .Q (signal_15296) ) ;
    buf_clk cell_10416 ( .C (clk), .D (signal_15303), .Q (signal_15304) ) ;
    buf_clk cell_10424 ( .C (clk), .D (signal_15311), .Q (signal_15312) ) ;
    buf_clk cell_10432 ( .C (clk), .D (signal_15319), .Q (signal_15320) ) ;
    buf_clk cell_10440 ( .C (clk), .D (signal_15327), .Q (signal_15328) ) ;
    buf_clk cell_10448 ( .C (clk), .D (signal_15335), .Q (signal_15336) ) ;
    buf_clk cell_10456 ( .C (clk), .D (signal_15343), .Q (signal_15344) ) ;
    buf_clk cell_10464 ( .C (clk), .D (signal_15351), .Q (signal_15352) ) ;
    buf_clk cell_10472 ( .C (clk), .D (signal_15359), .Q (signal_15360) ) ;
    buf_clk cell_10480 ( .C (clk), .D (signal_15367), .Q (signal_15368) ) ;
    buf_clk cell_10488 ( .C (clk), .D (signal_15375), .Q (signal_15376) ) ;
    buf_clk cell_10496 ( .C (clk), .D (signal_15383), .Q (signal_15384) ) ;
    buf_clk cell_10504 ( .C (clk), .D (signal_15391), .Q (signal_15392) ) ;
    buf_clk cell_10512 ( .C (clk), .D (signal_15399), .Q (signal_15400) ) ;
    buf_clk cell_10520 ( .C (clk), .D (signal_15407), .Q (signal_15408) ) ;
    buf_clk cell_10528 ( .C (clk), .D (signal_15415), .Q (signal_15416) ) ;
    buf_clk cell_10536 ( .C (clk), .D (signal_15423), .Q (signal_15424) ) ;
    buf_clk cell_10544 ( .C (clk), .D (signal_15431), .Q (signal_15432) ) ;
    buf_clk cell_10552 ( .C (clk), .D (signal_15439), .Q (signal_15440) ) ;
    buf_clk cell_10560 ( .C (clk), .D (signal_15447), .Q (signal_15448) ) ;
    buf_clk cell_10568 ( .C (clk), .D (signal_15455), .Q (signal_15456) ) ;
    buf_clk cell_10576 ( .C (clk), .D (signal_15463), .Q (signal_15464) ) ;
    buf_clk cell_10584 ( .C (clk), .D (signal_15471), .Q (signal_15472) ) ;
    buf_clk cell_10592 ( .C (clk), .D (signal_15479), .Q (signal_15480) ) ;
    buf_clk cell_10600 ( .C (clk), .D (signal_15487), .Q (signal_15488) ) ;
    buf_clk cell_10608 ( .C (clk), .D (signal_15495), .Q (signal_15496) ) ;
    buf_clk cell_10616 ( .C (clk), .D (signal_15503), .Q (signal_15504) ) ;
    buf_clk cell_10624 ( .C (clk), .D (signal_15511), .Q (signal_15512) ) ;
    buf_clk cell_10632 ( .C (clk), .D (signal_15519), .Q (signal_15520) ) ;
    buf_clk cell_10640 ( .C (clk), .D (signal_15527), .Q (signal_15528) ) ;
    buf_clk cell_10648 ( .C (clk), .D (signal_15535), .Q (signal_15536) ) ;
    buf_clk cell_10656 ( .C (clk), .D (signal_15543), .Q (signal_15544) ) ;
    buf_clk cell_10664 ( .C (clk), .D (signal_15551), .Q (signal_15552) ) ;
    buf_clk cell_10672 ( .C (clk), .D (signal_15559), .Q (signal_15560) ) ;
    buf_clk cell_10680 ( .C (clk), .D (signal_15567), .Q (signal_15568) ) ;
    buf_clk cell_10688 ( .C (clk), .D (signal_15575), .Q (signal_15576) ) ;
    buf_clk cell_10696 ( .C (clk), .D (signal_15583), .Q (signal_15584) ) ;
    buf_clk cell_10704 ( .C (clk), .D (signal_15591), .Q (signal_15592) ) ;
    buf_clk cell_10712 ( .C (clk), .D (signal_15599), .Q (signal_15600) ) ;
    buf_clk cell_10720 ( .C (clk), .D (signal_15607), .Q (signal_15608) ) ;
    buf_clk cell_10728 ( .C (clk), .D (signal_15615), .Q (signal_15616) ) ;
    buf_clk cell_10736 ( .C (clk), .D (signal_15623), .Q (signal_15624) ) ;
    buf_clk cell_10744 ( .C (clk), .D (signal_15631), .Q (signal_15632) ) ;
    buf_clk cell_10752 ( .C (clk), .D (signal_15639), .Q (signal_15640) ) ;
    buf_clk cell_10760 ( .C (clk), .D (signal_15647), .Q (signal_15648) ) ;
    buf_clk cell_10768 ( .C (clk), .D (signal_15655), .Q (signal_15656) ) ;
    buf_clk cell_10776 ( .C (clk), .D (signal_15663), .Q (signal_15664) ) ;
    buf_clk cell_10784 ( .C (clk), .D (signal_15671), .Q (signal_15672) ) ;
    buf_clk cell_10792 ( .C (clk), .D (signal_15679), .Q (signal_15680) ) ;
    buf_clk cell_10800 ( .C (clk), .D (signal_15687), .Q (signal_15688) ) ;
    buf_clk cell_10808 ( .C (clk), .D (signal_15695), .Q (signal_15696) ) ;
    buf_clk cell_10816 ( .C (clk), .D (signal_15703), .Q (signal_15704) ) ;
    buf_clk cell_10824 ( .C (clk), .D (signal_15711), .Q (signal_15712) ) ;
    buf_clk cell_10832 ( .C (clk), .D (signal_15719), .Q (signal_15720) ) ;
    buf_clk cell_10840 ( .C (clk), .D (signal_15727), .Q (signal_15728) ) ;
    buf_clk cell_10848 ( .C (clk), .D (signal_15735), .Q (signal_15736) ) ;
    buf_clk cell_10856 ( .C (clk), .D (signal_15743), .Q (signal_15744) ) ;
    buf_clk cell_10864 ( .C (clk), .D (signal_15751), .Q (signal_15752) ) ;
    buf_clk cell_10872 ( .C (clk), .D (signal_15759), .Q (signal_15760) ) ;
    buf_clk cell_10880 ( .C (clk), .D (signal_15767), .Q (signal_15768) ) ;
    buf_clk cell_10888 ( .C (clk), .D (signal_15775), .Q (signal_15776) ) ;
    buf_clk cell_10896 ( .C (clk), .D (signal_15783), .Q (signal_15784) ) ;
    buf_clk cell_10904 ( .C (clk), .D (signal_15791), .Q (signal_15792) ) ;
    buf_clk cell_10912 ( .C (clk), .D (signal_15799), .Q (signal_15800) ) ;
    buf_clk cell_10920 ( .C (clk), .D (signal_15807), .Q (signal_15808) ) ;
    buf_clk cell_10928 ( .C (clk), .D (signal_15815), .Q (signal_15816) ) ;
    buf_clk cell_10936 ( .C (clk), .D (signal_15823), .Q (signal_15824) ) ;
    buf_clk cell_10944 ( .C (clk), .D (signal_15831), .Q (signal_15832) ) ;
    buf_clk cell_10952 ( .C (clk), .D (signal_15839), .Q (signal_15840) ) ;
    buf_clk cell_10960 ( .C (clk), .D (signal_15847), .Q (signal_15848) ) ;
    buf_clk cell_10968 ( .C (clk), .D (signal_15855), .Q (signal_15856) ) ;
    buf_clk cell_10976 ( .C (clk), .D (signal_15863), .Q (signal_15864) ) ;
    buf_clk cell_10984 ( .C (clk), .D (signal_15871), .Q (signal_15872) ) ;
    buf_clk cell_10992 ( .C (clk), .D (signal_15879), .Q (signal_15880) ) ;
    buf_clk cell_11000 ( .C (clk), .D (signal_15887), .Q (signal_15888) ) ;
    buf_clk cell_11008 ( .C (clk), .D (signal_15895), .Q (signal_15896) ) ;
    buf_clk cell_11016 ( .C (clk), .D (signal_15903), .Q (signal_15904) ) ;
    buf_clk cell_11024 ( .C (clk), .D (signal_15911), .Q (signal_15912) ) ;
    buf_clk cell_11032 ( .C (clk), .D (signal_15919), .Q (signal_15920) ) ;
    buf_clk cell_11040 ( .C (clk), .D (signal_15927), .Q (signal_15928) ) ;
    buf_clk cell_11048 ( .C (clk), .D (signal_15935), .Q (signal_15936) ) ;
    buf_clk cell_11056 ( .C (clk), .D (signal_15943), .Q (signal_15944) ) ;
    buf_clk cell_11064 ( .C (clk), .D (signal_15951), .Q (signal_15952) ) ;
    buf_clk cell_11072 ( .C (clk), .D (signal_15959), .Q (signal_15960) ) ;
    buf_clk cell_11080 ( .C (clk), .D (signal_15967), .Q (signal_15968) ) ;
    buf_clk cell_11088 ( .C (clk), .D (signal_15975), .Q (signal_15976) ) ;
    buf_clk cell_11096 ( .C (clk), .D (signal_15983), .Q (signal_15984) ) ;
    buf_clk cell_11104 ( .C (clk), .D (signal_15991), .Q (signal_15992) ) ;
    buf_clk cell_11112 ( .C (clk), .D (signal_15999), .Q (signal_16000) ) ;
    buf_clk cell_11120 ( .C (clk), .D (signal_16007), .Q (signal_16008) ) ;
    buf_clk cell_11128 ( .C (clk), .D (signal_16015), .Q (signal_16016) ) ;
    buf_clk cell_11136 ( .C (clk), .D (signal_16023), .Q (signal_16024) ) ;
    buf_clk cell_11144 ( .C (clk), .D (signal_16031), .Q (signal_16032) ) ;
    buf_clk cell_11152 ( .C (clk), .D (signal_16039), .Q (signal_16040) ) ;
    buf_clk cell_11160 ( .C (clk), .D (signal_16047), .Q (signal_16048) ) ;
    buf_clk cell_11168 ( .C (clk), .D (signal_16055), .Q (signal_16056) ) ;
    buf_clk cell_11176 ( .C (clk), .D (signal_16063), .Q (signal_16064) ) ;
    buf_clk cell_11184 ( .C (clk), .D (signal_16071), .Q (signal_16072) ) ;
    buf_clk cell_11192 ( .C (clk), .D (signal_16079), .Q (signal_16080) ) ;
    buf_clk cell_11200 ( .C (clk), .D (signal_16087), .Q (signal_16088) ) ;
    buf_clk cell_11208 ( .C (clk), .D (signal_16095), .Q (signal_16096) ) ;
    buf_clk cell_11216 ( .C (clk), .D (signal_16103), .Q (signal_16104) ) ;
    buf_clk cell_11224 ( .C (clk), .D (signal_16111), .Q (signal_16112) ) ;
    buf_clk cell_11232 ( .C (clk), .D (signal_16119), .Q (signal_16120) ) ;
    buf_clk cell_11240 ( .C (clk), .D (signal_16127), .Q (signal_16128) ) ;
    buf_clk cell_11248 ( .C (clk), .D (signal_16135), .Q (signal_16136) ) ;
    buf_clk cell_11256 ( .C (clk), .D (signal_16143), .Q (signal_16144) ) ;
    buf_clk cell_11264 ( .C (clk), .D (signal_16151), .Q (signal_16152) ) ;
    buf_clk cell_11272 ( .C (clk), .D (signal_16159), .Q (signal_16160) ) ;
    buf_clk cell_11280 ( .C (clk), .D (signal_16167), .Q (signal_16168) ) ;
    buf_clk cell_11288 ( .C (clk), .D (signal_16175), .Q (signal_16176) ) ;
    buf_clk cell_11296 ( .C (clk), .D (signal_16183), .Q (signal_16184) ) ;
    buf_clk cell_11304 ( .C (clk), .D (signal_16191), .Q (signal_16192) ) ;
    buf_clk cell_11312 ( .C (clk), .D (signal_16199), .Q (signal_16200) ) ;
    buf_clk cell_11320 ( .C (clk), .D (signal_16207), .Q (signal_16208) ) ;
    buf_clk cell_11328 ( .C (clk), .D (signal_16215), .Q (signal_16216) ) ;
    buf_clk cell_11336 ( .C (clk), .D (signal_16223), .Q (signal_16224) ) ;
    buf_clk cell_11344 ( .C (clk), .D (signal_16231), .Q (signal_16232) ) ;
    buf_clk cell_11352 ( .C (clk), .D (signal_16239), .Q (signal_16240) ) ;
    buf_clk cell_11360 ( .C (clk), .D (signal_16247), .Q (signal_16248) ) ;
    buf_clk cell_11368 ( .C (clk), .D (signal_16255), .Q (signal_16256) ) ;
    buf_clk cell_11376 ( .C (clk), .D (signal_16263), .Q (signal_16264) ) ;
    buf_clk cell_11384 ( .C (clk), .D (signal_16271), .Q (signal_16272) ) ;
    buf_clk cell_11392 ( .C (clk), .D (signal_16279), .Q (signal_16280) ) ;
    buf_clk cell_11400 ( .C (clk), .D (signal_16287), .Q (signal_16288) ) ;
    buf_clk cell_11408 ( .C (clk), .D (signal_16295), .Q (signal_16296) ) ;
    buf_clk cell_11416 ( .C (clk), .D (signal_16303), .Q (signal_16304) ) ;
    buf_clk cell_11424 ( .C (clk), .D (signal_16311), .Q (signal_16312) ) ;
    buf_clk cell_11432 ( .C (clk), .D (signal_16319), .Q (signal_16320) ) ;
    buf_clk cell_11440 ( .C (clk), .D (signal_16327), .Q (signal_16328) ) ;
    buf_clk cell_11448 ( .C (clk), .D (signal_16335), .Q (signal_16336) ) ;
    buf_clk cell_11456 ( .C (clk), .D (signal_16343), .Q (signal_16344) ) ;
    buf_clk cell_11464 ( .C (clk), .D (signal_16351), .Q (signal_16352) ) ;
    buf_clk cell_11472 ( .C (clk), .D (signal_16359), .Q (signal_16360) ) ;
    buf_clk cell_11480 ( .C (clk), .D (signal_16367), .Q (signal_16368) ) ;
    buf_clk cell_11488 ( .C (clk), .D (signal_16375), .Q (signal_16376) ) ;
    buf_clk cell_11496 ( .C (clk), .D (signal_16383), .Q (signal_16384) ) ;
    buf_clk cell_11504 ( .C (clk), .D (signal_16391), .Q (signal_16392) ) ;
    buf_clk cell_11512 ( .C (clk), .D (signal_16399), .Q (signal_16400) ) ;
    buf_clk cell_11520 ( .C (clk), .D (signal_16407), .Q (signal_16408) ) ;
    buf_clk cell_11528 ( .C (clk), .D (signal_16415), .Q (signal_16416) ) ;
    buf_clk cell_11536 ( .C (clk), .D (signal_16423), .Q (signal_16424) ) ;
    buf_clk cell_11544 ( .C (clk), .D (signal_16431), .Q (signal_16432) ) ;
    buf_clk cell_11552 ( .C (clk), .D (signal_16439), .Q (signal_16440) ) ;
    buf_clk cell_11560 ( .C (clk), .D (signal_16447), .Q (signal_16448) ) ;
    buf_clk cell_11568 ( .C (clk), .D (signal_16455), .Q (signal_16456) ) ;
    buf_clk cell_11576 ( .C (clk), .D (signal_16463), .Q (signal_16464) ) ;
    buf_clk cell_11584 ( .C (clk), .D (signal_16471), .Q (signal_16472) ) ;
    buf_clk cell_11592 ( .C (clk), .D (signal_16479), .Q (signal_16480) ) ;
    buf_clk cell_11600 ( .C (clk), .D (signal_16487), .Q (signal_16488) ) ;
    buf_clk cell_11608 ( .C (clk), .D (signal_16495), .Q (signal_16496) ) ;
    buf_clk cell_11616 ( .C (clk), .D (signal_16503), .Q (signal_16504) ) ;
    buf_clk cell_11624 ( .C (clk), .D (signal_16511), .Q (signal_16512) ) ;
    buf_clk cell_11632 ( .C (clk), .D (signal_16519), .Q (signal_16520) ) ;
    buf_clk cell_11640 ( .C (clk), .D (signal_16527), .Q (signal_16528) ) ;
    buf_clk cell_11648 ( .C (clk), .D (signal_16535), .Q (signal_16536) ) ;
    buf_clk cell_11656 ( .C (clk), .D (signal_16543), .Q (signal_16544) ) ;
    buf_clk cell_11664 ( .C (clk), .D (signal_16551), .Q (signal_16552) ) ;
    buf_clk cell_11672 ( .C (clk), .D (signal_16559), .Q (signal_16560) ) ;
    buf_clk cell_11680 ( .C (clk), .D (signal_16567), .Q (signal_16568) ) ;
    buf_clk cell_11688 ( .C (clk), .D (signal_16575), .Q (signal_16576) ) ;
    buf_clk cell_11696 ( .C (clk), .D (signal_16583), .Q (signal_16584) ) ;
    buf_clk cell_11704 ( .C (clk), .D (signal_16591), .Q (signal_16592) ) ;
    buf_clk cell_11712 ( .C (clk), .D (signal_16599), .Q (signal_16600) ) ;
    buf_clk cell_11720 ( .C (clk), .D (signal_16607), .Q (signal_16608) ) ;
    buf_clk cell_11728 ( .C (clk), .D (signal_16615), .Q (signal_16616) ) ;
    buf_clk cell_11736 ( .C (clk), .D (signal_16623), .Q (signal_16624) ) ;
    buf_clk cell_11744 ( .C (clk), .D (signal_16631), .Q (signal_16632) ) ;
    buf_clk cell_11752 ( .C (clk), .D (signal_16639), .Q (signal_16640) ) ;
    buf_clk cell_11760 ( .C (clk), .D (signal_16647), .Q (signal_16648) ) ;
    buf_clk cell_11768 ( .C (clk), .D (signal_16655), .Q (signal_16656) ) ;
    buf_clk cell_11776 ( .C (clk), .D (signal_16663), .Q (signal_16664) ) ;
    buf_clk cell_11784 ( .C (clk), .D (signal_16671), .Q (signal_16672) ) ;
    buf_clk cell_11792 ( .C (clk), .D (signal_16679), .Q (signal_16680) ) ;
    buf_clk cell_11800 ( .C (clk), .D (signal_16687), .Q (signal_16688) ) ;
    buf_clk cell_11808 ( .C (clk), .D (signal_16695), .Q (signal_16696) ) ;
    buf_clk cell_11816 ( .C (clk), .D (signal_16703), .Q (signal_16704) ) ;
    buf_clk cell_11824 ( .C (clk), .D (signal_16711), .Q (signal_16712) ) ;
    buf_clk cell_11832 ( .C (clk), .D (signal_16719), .Q (signal_16720) ) ;
    buf_clk cell_11840 ( .C (clk), .D (signal_16727), .Q (signal_16728) ) ;
    buf_clk cell_11848 ( .C (clk), .D (signal_16735), .Q (signal_16736) ) ;
    buf_clk cell_11856 ( .C (clk), .D (signal_16743), .Q (signal_16744) ) ;
    buf_clk cell_11864 ( .C (clk), .D (signal_16751), .Q (signal_16752) ) ;
    buf_clk cell_11872 ( .C (clk), .D (signal_16759), .Q (signal_16760) ) ;
    buf_clk cell_11880 ( .C (clk), .D (signal_16767), .Q (signal_16768) ) ;
    buf_clk cell_11888 ( .C (clk), .D (signal_16775), .Q (signal_16776) ) ;
    buf_clk cell_11896 ( .C (clk), .D (signal_16783), .Q (signal_16784) ) ;
    buf_clk cell_11904 ( .C (clk), .D (signal_16791), .Q (signal_16792) ) ;
    buf_clk cell_11912 ( .C (clk), .D (signal_16799), .Q (signal_16800) ) ;
    buf_clk cell_11920 ( .C (clk), .D (signal_16807), .Q (signal_16808) ) ;
    buf_clk cell_11928 ( .C (clk), .D (signal_16815), .Q (signal_16816) ) ;
    buf_clk cell_11936 ( .C (clk), .D (signal_16823), .Q (signal_16824) ) ;
    buf_clk cell_11944 ( .C (clk), .D (signal_16831), .Q (signal_16832) ) ;
    buf_clk cell_11952 ( .C (clk), .D (signal_16839), .Q (signal_16840) ) ;
    buf_clk cell_11960 ( .C (clk), .D (signal_16847), .Q (signal_16848) ) ;
    buf_clk cell_11968 ( .C (clk), .D (signal_16855), .Q (signal_16856) ) ;
    buf_clk cell_11976 ( .C (clk), .D (signal_16863), .Q (signal_16864) ) ;
    buf_clk cell_11984 ( .C (clk), .D (signal_16871), .Q (signal_16872) ) ;
    buf_clk cell_11992 ( .C (clk), .D (signal_16879), .Q (signal_16880) ) ;
    buf_clk cell_12000 ( .C (clk), .D (signal_16887), .Q (signal_16888) ) ;
    buf_clk cell_12008 ( .C (clk), .D (signal_16895), .Q (signal_16896) ) ;
    buf_clk cell_12016 ( .C (clk), .D (signal_16903), .Q (signal_16904) ) ;
    buf_clk cell_12024 ( .C (clk), .D (signal_16911), .Q (signal_16912) ) ;
    buf_clk cell_12032 ( .C (clk), .D (signal_16919), .Q (signal_16920) ) ;
    buf_clk cell_12040 ( .C (clk), .D (signal_16927), .Q (signal_16928) ) ;
    buf_clk cell_12048 ( .C (clk), .D (signal_16935), .Q (signal_16936) ) ;
    buf_clk cell_12056 ( .C (clk), .D (signal_16943), .Q (signal_16944) ) ;
    buf_clk cell_12064 ( .C (clk), .D (signal_16951), .Q (signal_16952) ) ;
    buf_clk cell_12072 ( .C (clk), .D (signal_16959), .Q (signal_16960) ) ;
    buf_clk cell_12080 ( .C (clk), .D (signal_16967), .Q (signal_16968) ) ;
    buf_clk cell_12088 ( .C (clk), .D (signal_16975), .Q (signal_16976) ) ;
    buf_clk cell_12096 ( .C (clk), .D (signal_16983), .Q (signal_16984) ) ;
    buf_clk cell_12104 ( .C (clk), .D (signal_16991), .Q (signal_16992) ) ;
    buf_clk cell_12112 ( .C (clk), .D (signal_16999), .Q (signal_17000) ) ;
    buf_clk cell_12120 ( .C (clk), .D (signal_17007), .Q (signal_17008) ) ;
    buf_clk cell_12128 ( .C (clk), .D (signal_17015), .Q (signal_17016) ) ;
    buf_clk cell_12136 ( .C (clk), .D (signal_17023), .Q (signal_17024) ) ;
    buf_clk cell_12144 ( .C (clk), .D (signal_17031), .Q (signal_17032) ) ;
    buf_clk cell_12152 ( .C (clk), .D (signal_17039), .Q (signal_17040) ) ;
    buf_clk cell_12160 ( .C (clk), .D (signal_17047), .Q (signal_17048) ) ;
    buf_clk cell_12168 ( .C (clk), .D (signal_17055), .Q (signal_17056) ) ;
    buf_clk cell_12176 ( .C (clk), .D (signal_17063), .Q (signal_17064) ) ;
    buf_clk cell_12184 ( .C (clk), .D (signal_17071), .Q (signal_17072) ) ;
    buf_clk cell_12192 ( .C (clk), .D (signal_17079), .Q (signal_17080) ) ;
    buf_clk cell_12200 ( .C (clk), .D (signal_17087), .Q (signal_17088) ) ;
    buf_clk cell_12208 ( .C (clk), .D (signal_17095), .Q (signal_17096) ) ;
    buf_clk cell_12216 ( .C (clk), .D (signal_17103), .Q (signal_17104) ) ;
    buf_clk cell_12224 ( .C (clk), .D (signal_17111), .Q (signal_17112) ) ;
    buf_clk cell_12232 ( .C (clk), .D (signal_17119), .Q (signal_17120) ) ;
    buf_clk cell_12240 ( .C (clk), .D (signal_17127), .Q (signal_17128) ) ;
    buf_clk cell_12248 ( .C (clk), .D (signal_17135), .Q (signal_17136) ) ;
    buf_clk cell_12256 ( .C (clk), .D (signal_17143), .Q (signal_17144) ) ;
    buf_clk cell_12264 ( .C (clk), .D (signal_17151), .Q (signal_17152) ) ;
    buf_clk cell_12272 ( .C (clk), .D (signal_17159), .Q (signal_17160) ) ;
    buf_clk cell_12280 ( .C (clk), .D (signal_17167), .Q (signal_17168) ) ;
    buf_clk cell_12288 ( .C (clk), .D (signal_17175), .Q (signal_17176) ) ;
    buf_clk cell_12296 ( .C (clk), .D (signal_17183), .Q (signal_17184) ) ;
    buf_clk cell_12304 ( .C (clk), .D (signal_17191), .Q (signal_17192) ) ;
    buf_clk cell_12312 ( .C (clk), .D (signal_17199), .Q (signal_17200) ) ;
    buf_clk cell_12320 ( .C (clk), .D (signal_17207), .Q (signal_17208) ) ;
    buf_clk cell_12328 ( .C (clk), .D (signal_17215), .Q (signal_17216) ) ;
    buf_clk cell_12336 ( .C (clk), .D (signal_17223), .Q (signal_17224) ) ;
    buf_clk cell_12344 ( .C (clk), .D (signal_17231), .Q (signal_17232) ) ;
    buf_clk cell_12352 ( .C (clk), .D (signal_17239), .Q (signal_17240) ) ;
    buf_clk cell_12360 ( .C (clk), .D (signal_17247), .Q (signal_17248) ) ;
    buf_clk cell_12368 ( .C (clk), .D (signal_17255), .Q (signal_17256) ) ;
    buf_clk cell_12376 ( .C (clk), .D (signal_17263), .Q (signal_17264) ) ;
    buf_clk cell_12384 ( .C (clk), .D (signal_17271), .Q (signal_17272) ) ;
    buf_clk cell_12392 ( .C (clk), .D (signal_17279), .Q (signal_17280) ) ;
    buf_clk cell_12400 ( .C (clk), .D (signal_17287), .Q (signal_17288) ) ;
    buf_clk cell_12408 ( .C (clk), .D (signal_17295), .Q (signal_17296) ) ;
    buf_clk cell_12416 ( .C (clk), .D (signal_17303), .Q (signal_17304) ) ;
    buf_clk cell_12424 ( .C (clk), .D (signal_17311), .Q (signal_17312) ) ;
    buf_clk cell_12432 ( .C (clk), .D (signal_17319), .Q (signal_17320) ) ;
    buf_clk cell_12440 ( .C (clk), .D (signal_17327), .Q (signal_17328) ) ;
    buf_clk cell_12448 ( .C (clk), .D (signal_17335), .Q (signal_17336) ) ;
    buf_clk cell_12456 ( .C (clk), .D (signal_17343), .Q (signal_17344) ) ;
    buf_clk cell_12464 ( .C (clk), .D (signal_17351), .Q (signal_17352) ) ;
    buf_clk cell_12472 ( .C (clk), .D (signal_17359), .Q (signal_17360) ) ;
    buf_clk cell_12480 ( .C (clk), .D (signal_17367), .Q (signal_17368) ) ;
    buf_clk cell_12488 ( .C (clk), .D (signal_17375), .Q (signal_17376) ) ;
    buf_clk cell_12496 ( .C (clk), .D (signal_17383), .Q (signal_17384) ) ;
    buf_clk cell_12504 ( .C (clk), .D (signal_17391), .Q (signal_17392) ) ;
    buf_clk cell_12512 ( .C (clk), .D (signal_17399), .Q (signal_17400) ) ;
    buf_clk cell_12520 ( .C (clk), .D (signal_17407), .Q (signal_17408) ) ;
    buf_clk cell_12528 ( .C (clk), .D (signal_17415), .Q (signal_17416) ) ;
    buf_clk cell_12536 ( .C (clk), .D (signal_17423), .Q (signal_17424) ) ;
    buf_clk cell_12544 ( .C (clk), .D (signal_17431), .Q (signal_17432) ) ;
    buf_clk cell_12552 ( .C (clk), .D (signal_17439), .Q (signal_17440) ) ;
    buf_clk cell_12560 ( .C (clk), .D (signal_17447), .Q (signal_17448) ) ;
    buf_clk cell_12568 ( .C (clk), .D (signal_17455), .Q (signal_17456) ) ;
    buf_clk cell_12576 ( .C (clk), .D (signal_17463), .Q (signal_17464) ) ;
    buf_clk cell_12584 ( .C (clk), .D (signal_17471), .Q (signal_17472) ) ;
    buf_clk cell_12592 ( .C (clk), .D (signal_17479), .Q (signal_17480) ) ;
    buf_clk cell_12600 ( .C (clk), .D (signal_17487), .Q (signal_17488) ) ;
    buf_clk cell_12608 ( .C (clk), .D (signal_17495), .Q (signal_17496) ) ;
    buf_clk cell_12616 ( .C (clk), .D (signal_17503), .Q (signal_17504) ) ;
    buf_clk cell_12624 ( .C (clk), .D (signal_17511), .Q (signal_17512) ) ;
    buf_clk cell_12632 ( .C (clk), .D (signal_17519), .Q (signal_17520) ) ;
    buf_clk cell_12640 ( .C (clk), .D (signal_17527), .Q (signal_17528) ) ;
    buf_clk cell_12648 ( .C (clk), .D (signal_17535), .Q (signal_17536) ) ;
    buf_clk cell_12656 ( .C (clk), .D (signal_17543), .Q (signal_17544) ) ;
    buf_clk cell_12664 ( .C (clk), .D (signal_17551), .Q (signal_17552) ) ;
    buf_clk cell_12672 ( .C (clk), .D (signal_17559), .Q (signal_17560) ) ;
    buf_clk cell_12680 ( .C (clk), .D (signal_17567), .Q (signal_17568) ) ;
    buf_clk cell_12688 ( .C (clk), .D (signal_17575), .Q (signal_17576) ) ;
    buf_clk cell_12696 ( .C (clk), .D (signal_17583), .Q (signal_17584) ) ;
    buf_clk cell_12704 ( .C (clk), .D (signal_17591), .Q (signal_17592) ) ;
    buf_clk cell_12712 ( .C (clk), .D (signal_17599), .Q (signal_17600) ) ;
    buf_clk cell_12720 ( .C (clk), .D (signal_17607), .Q (signal_17608) ) ;
    buf_clk cell_12728 ( .C (clk), .D (signal_17615), .Q (signal_17616) ) ;
    buf_clk cell_12736 ( .C (clk), .D (signal_17623), .Q (signal_17624) ) ;
    buf_clk cell_12744 ( .C (clk), .D (signal_17631), .Q (signal_17632) ) ;
    buf_clk cell_12752 ( .C (clk), .D (signal_17639), .Q (signal_17640) ) ;
    buf_clk cell_12760 ( .C (clk), .D (signal_17647), .Q (signal_17648) ) ;
    buf_clk cell_12768 ( .C (clk), .D (signal_17655), .Q (signal_17656) ) ;
    buf_clk cell_12776 ( .C (clk), .D (signal_17663), .Q (signal_17664) ) ;
    buf_clk cell_12784 ( .C (clk), .D (signal_17671), .Q (signal_17672) ) ;
    buf_clk cell_12792 ( .C (clk), .D (signal_17679), .Q (signal_17680) ) ;
    buf_clk cell_12800 ( .C (clk), .D (signal_17687), .Q (signal_17688) ) ;
    buf_clk cell_12808 ( .C (clk), .D (signal_17695), .Q (signal_17696) ) ;
    buf_clk cell_12816 ( .C (clk), .D (signal_17703), .Q (signal_17704) ) ;
    buf_clk cell_12824 ( .C (clk), .D (signal_17711), .Q (signal_17712) ) ;
    buf_clk cell_12832 ( .C (clk), .D (signal_17719), .Q (signal_17720) ) ;
    buf_clk cell_12840 ( .C (clk), .D (signal_17727), .Q (signal_17728) ) ;
    buf_clk cell_12848 ( .C (clk), .D (signal_17735), .Q (signal_17736) ) ;
    buf_clk cell_12856 ( .C (clk), .D (signal_17743), .Q (signal_17744) ) ;
    buf_clk cell_12864 ( .C (clk), .D (signal_17751), .Q (signal_17752) ) ;
    buf_clk cell_12872 ( .C (clk), .D (signal_17759), .Q (signal_17760) ) ;
    buf_clk cell_12880 ( .C (clk), .D (signal_17767), .Q (signal_17768) ) ;
    buf_clk cell_12888 ( .C (clk), .D (signal_17775), .Q (signal_17776) ) ;
    buf_clk cell_12896 ( .C (clk), .D (signal_17783), .Q (signal_17784) ) ;
    buf_clk cell_12904 ( .C (clk), .D (signal_17791), .Q (signal_17792) ) ;
    buf_clk cell_12912 ( .C (clk), .D (signal_17799), .Q (signal_17800) ) ;
    buf_clk cell_12920 ( .C (clk), .D (signal_17807), .Q (signal_17808) ) ;
    buf_clk cell_12928 ( .C (clk), .D (signal_17815), .Q (signal_17816) ) ;
    buf_clk cell_12936 ( .C (clk), .D (signal_17823), .Q (signal_17824) ) ;
    buf_clk cell_12944 ( .C (clk), .D (signal_17831), .Q (signal_17832) ) ;
    buf_clk cell_12952 ( .C (clk), .D (signal_17839), .Q (signal_17840) ) ;
    buf_clk cell_12960 ( .C (clk), .D (signal_17847), .Q (signal_17848) ) ;
    buf_clk cell_12968 ( .C (clk), .D (signal_17855), .Q (signal_17856) ) ;
    buf_clk cell_12976 ( .C (clk), .D (signal_17863), .Q (signal_17864) ) ;
    buf_clk cell_12984 ( .C (clk), .D (signal_17871), .Q (signal_17872) ) ;
    buf_clk cell_12992 ( .C (clk), .D (signal_17879), .Q (signal_17880) ) ;
    buf_clk cell_13000 ( .C (clk), .D (signal_17887), .Q (signal_17888) ) ;
    buf_clk cell_13008 ( .C (clk), .D (signal_17895), .Q (signal_17896) ) ;
    buf_clk cell_13016 ( .C (clk), .D (signal_17903), .Q (signal_17904) ) ;
    buf_clk cell_13024 ( .C (clk), .D (signal_17911), .Q (signal_17912) ) ;
    buf_clk cell_13032 ( .C (clk), .D (signal_17919), .Q (signal_17920) ) ;
    buf_clk cell_13040 ( .C (clk), .D (signal_17927), .Q (signal_17928) ) ;
    buf_clk cell_13048 ( .C (clk), .D (signal_17935), .Q (signal_17936) ) ;
    buf_clk cell_13056 ( .C (clk), .D (signal_17943), .Q (signal_17944) ) ;
    buf_clk cell_13064 ( .C (clk), .D (signal_17951), .Q (signal_17952) ) ;
    buf_clk cell_13072 ( .C (clk), .D (signal_17959), .Q (signal_17960) ) ;
    buf_clk cell_13080 ( .C (clk), .D (signal_17967), .Q (signal_17968) ) ;
    buf_clk cell_13088 ( .C (clk), .D (signal_17975), .Q (signal_17976) ) ;
    buf_clk cell_13096 ( .C (clk), .D (signal_17983), .Q (signal_17984) ) ;
    buf_clk cell_13104 ( .C (clk), .D (signal_17991), .Q (signal_17992) ) ;
    buf_clk cell_13112 ( .C (clk), .D (signal_17999), .Q (signal_18000) ) ;
    buf_clk cell_13120 ( .C (clk), .D (signal_18007), .Q (signal_18008) ) ;
    buf_clk cell_13128 ( .C (clk), .D (signal_18015), .Q (signal_18016) ) ;
    buf_clk cell_13136 ( .C (clk), .D (signal_18023), .Q (signal_18024) ) ;
    buf_clk cell_13144 ( .C (clk), .D (signal_18031), .Q (signal_18032) ) ;
    buf_clk cell_13152 ( .C (clk), .D (signal_18039), .Q (signal_18040) ) ;
    buf_clk cell_13160 ( .C (clk), .D (signal_18047), .Q (signal_18048) ) ;
    buf_clk cell_13168 ( .C (clk), .D (signal_18055), .Q (signal_18056) ) ;
    buf_clk cell_13176 ( .C (clk), .D (signal_18063), .Q (signal_18064) ) ;
    buf_clk cell_13184 ( .C (clk), .D (signal_18071), .Q (signal_18072) ) ;
    buf_clk cell_13192 ( .C (clk), .D (signal_18079), .Q (signal_18080) ) ;
    buf_clk cell_13200 ( .C (clk), .D (signal_18087), .Q (signal_18088) ) ;
    buf_clk cell_13208 ( .C (clk), .D (signal_18095), .Q (signal_18096) ) ;
    buf_clk cell_13216 ( .C (clk), .D (signal_18103), .Q (signal_18104) ) ;
    buf_clk cell_13224 ( .C (clk), .D (signal_18111), .Q (signal_18112) ) ;
    buf_clk cell_13232 ( .C (clk), .D (signal_18119), .Q (signal_18120) ) ;
    buf_clk cell_13240 ( .C (clk), .D (signal_18127), .Q (signal_18128) ) ;
    buf_clk cell_13248 ( .C (clk), .D (signal_18135), .Q (signal_18136) ) ;
    buf_clk cell_13256 ( .C (clk), .D (signal_18143), .Q (signal_18144) ) ;
    buf_clk cell_13264 ( .C (clk), .D (signal_18151), .Q (signal_18152) ) ;
    buf_clk cell_13272 ( .C (clk), .D (signal_18159), .Q (signal_18160) ) ;
    buf_clk cell_13280 ( .C (clk), .D (signal_18167), .Q (signal_18168) ) ;
    buf_clk cell_13286 ( .C (clk), .D (signal_18173), .Q (signal_18174) ) ;
    buf_clk cell_13292 ( .C (clk), .D (signal_18179), .Q (signal_18180) ) ;
    buf_clk cell_13298 ( .C (clk), .D (signal_18185), .Q (signal_18186) ) ;
    buf_clk cell_13304 ( .C (clk), .D (signal_18191), .Q (signal_18192) ) ;
    buf_clk cell_13310 ( .C (clk), .D (signal_18197), .Q (signal_18198) ) ;
    buf_clk cell_13316 ( .C (clk), .D (signal_18203), .Q (signal_18204) ) ;
    buf_clk cell_13322 ( .C (clk), .D (signal_18209), .Q (signal_18210) ) ;
    buf_clk cell_13328 ( .C (clk), .D (signal_18215), .Q (signal_18216) ) ;
    buf_clk cell_13334 ( .C (clk), .D (signal_18221), .Q (signal_18222) ) ;
    buf_clk cell_13340 ( .C (clk), .D (signal_18227), .Q (signal_18228) ) ;
    buf_clk cell_13346 ( .C (clk), .D (signal_18233), .Q (signal_18234) ) ;
    buf_clk cell_13352 ( .C (clk), .D (signal_18239), .Q (signal_18240) ) ;
    buf_clk cell_13358 ( .C (clk), .D (signal_18245), .Q (signal_18246) ) ;
    buf_clk cell_13364 ( .C (clk), .D (signal_18251), .Q (signal_18252) ) ;
    buf_clk cell_13370 ( .C (clk), .D (signal_18257), .Q (signal_18258) ) ;
    buf_clk cell_13376 ( .C (clk), .D (signal_18263), .Q (signal_18264) ) ;
    buf_clk cell_13382 ( .C (clk), .D (signal_18269), .Q (signal_18270) ) ;
    buf_clk cell_13388 ( .C (clk), .D (signal_18275), .Q (signal_18276) ) ;
    buf_clk cell_13394 ( .C (clk), .D (signal_18281), .Q (signal_18282) ) ;
    buf_clk cell_13400 ( .C (clk), .D (signal_18287), .Q (signal_18288) ) ;
    buf_clk cell_13406 ( .C (clk), .D (signal_18293), .Q (signal_18294) ) ;
    buf_clk cell_13412 ( .C (clk), .D (signal_18299), .Q (signal_18300) ) ;
    buf_clk cell_13418 ( .C (clk), .D (signal_18305), .Q (signal_18306) ) ;
    buf_clk cell_13424 ( .C (clk), .D (signal_18311), .Q (signal_18312) ) ;
    buf_clk cell_13430 ( .C (clk), .D (signal_18317), .Q (signal_18318) ) ;
    buf_clk cell_13436 ( .C (clk), .D (signal_18323), .Q (signal_18324) ) ;
    buf_clk cell_13442 ( .C (clk), .D (signal_18329), .Q (signal_18330) ) ;
    buf_clk cell_13448 ( .C (clk), .D (signal_18335), .Q (signal_18336) ) ;
    buf_clk cell_13454 ( .C (clk), .D (signal_18341), .Q (signal_18342) ) ;
    buf_clk cell_13460 ( .C (clk), .D (signal_18347), .Q (signal_18348) ) ;
    buf_clk cell_13466 ( .C (clk), .D (signal_18353), .Q (signal_18354) ) ;
    buf_clk cell_13472 ( .C (clk), .D (signal_18359), .Q (signal_18360) ) ;
    buf_clk cell_13478 ( .C (clk), .D (signal_18365), .Q (signal_18366) ) ;
    buf_clk cell_13484 ( .C (clk), .D (signal_18371), .Q (signal_18372) ) ;
    buf_clk cell_13490 ( .C (clk), .D (signal_18377), .Q (signal_18378) ) ;
    buf_clk cell_13496 ( .C (clk), .D (signal_18383), .Q (signal_18384) ) ;
    buf_clk cell_13502 ( .C (clk), .D (signal_18389), .Q (signal_18390) ) ;
    buf_clk cell_13508 ( .C (clk), .D (signal_18395), .Q (signal_18396) ) ;
    buf_clk cell_13514 ( .C (clk), .D (signal_18401), .Q (signal_18402) ) ;
    buf_clk cell_13520 ( .C (clk), .D (signal_18407), .Q (signal_18408) ) ;
    buf_clk cell_13526 ( .C (clk), .D (signal_18413), .Q (signal_18414) ) ;
    buf_clk cell_13532 ( .C (clk), .D (signal_18419), .Q (signal_18420) ) ;
    buf_clk cell_13538 ( .C (clk), .D (signal_18425), .Q (signal_18426) ) ;
    buf_clk cell_13544 ( .C (clk), .D (signal_18431), .Q (signal_18432) ) ;
    buf_clk cell_13550 ( .C (clk), .D (signal_18437), .Q (signal_18438) ) ;
    buf_clk cell_13556 ( .C (clk), .D (signal_18443), .Q (signal_18444) ) ;
    buf_clk cell_13562 ( .C (clk), .D (signal_18449), .Q (signal_18450) ) ;
    buf_clk cell_13568 ( .C (clk), .D (signal_18455), .Q (signal_18456) ) ;
    buf_clk cell_13574 ( .C (clk), .D (signal_18461), .Q (signal_18462) ) ;
    buf_clk cell_13580 ( .C (clk), .D (signal_18467), .Q (signal_18468) ) ;
    buf_clk cell_13586 ( .C (clk), .D (signal_18473), .Q (signal_18474) ) ;
    buf_clk cell_13592 ( .C (clk), .D (signal_18479), .Q (signal_18480) ) ;
    buf_clk cell_13598 ( .C (clk), .D (signal_18485), .Q (signal_18486) ) ;
    buf_clk cell_13604 ( .C (clk), .D (signal_18491), .Q (signal_18492) ) ;
    buf_clk cell_13610 ( .C (clk), .D (signal_18497), .Q (signal_18498) ) ;
    buf_clk cell_13616 ( .C (clk), .D (signal_18503), .Q (signal_18504) ) ;
    buf_clk cell_13622 ( .C (clk), .D (signal_18509), .Q (signal_18510) ) ;
    buf_clk cell_13628 ( .C (clk), .D (signal_18515), .Q (signal_18516) ) ;
    buf_clk cell_13634 ( .C (clk), .D (signal_18521), .Q (signal_18522) ) ;
    buf_clk cell_13640 ( .C (clk), .D (signal_18527), .Q (signal_18528) ) ;
    buf_clk cell_13646 ( .C (clk), .D (signal_18533), .Q (signal_18534) ) ;
    buf_clk cell_13652 ( .C (clk), .D (signal_18539), .Q (signal_18540) ) ;
    buf_clk cell_13658 ( .C (clk), .D (signal_18545), .Q (signal_18546) ) ;
    buf_clk cell_13664 ( .C (clk), .D (signal_18551), .Q (signal_18552) ) ;
    buf_clk cell_13670 ( .C (clk), .D (signal_18557), .Q (signal_18558) ) ;
    buf_clk cell_13676 ( .C (clk), .D (signal_18563), .Q (signal_18564) ) ;
    buf_clk cell_13682 ( .C (clk), .D (signal_18569), .Q (signal_18570) ) ;
    buf_clk cell_13688 ( .C (clk), .D (signal_18575), .Q (signal_18576) ) ;
    buf_clk cell_13694 ( .C (clk), .D (signal_18581), .Q (signal_18582) ) ;
    buf_clk cell_13700 ( .C (clk), .D (signal_18587), .Q (signal_18588) ) ;
    buf_clk cell_13706 ( .C (clk), .D (signal_18593), .Q (signal_18594) ) ;
    buf_clk cell_13712 ( .C (clk), .D (signal_18599), .Q (signal_18600) ) ;
    buf_clk cell_13718 ( .C (clk), .D (signal_18605), .Q (signal_18606) ) ;
    buf_clk cell_13724 ( .C (clk), .D (signal_18611), .Q (signal_18612) ) ;
    buf_clk cell_13730 ( .C (clk), .D (signal_18617), .Q (signal_18618) ) ;
    buf_clk cell_13736 ( .C (clk), .D (signal_18623), .Q (signal_18624) ) ;
    buf_clk cell_13742 ( .C (clk), .D (signal_18629), .Q (signal_18630) ) ;
    buf_clk cell_13748 ( .C (clk), .D (signal_18635), .Q (signal_18636) ) ;
    buf_clk cell_13754 ( .C (clk), .D (signal_18641), .Q (signal_18642) ) ;
    buf_clk cell_13760 ( .C (clk), .D (signal_18647), .Q (signal_18648) ) ;
    buf_clk cell_13766 ( .C (clk), .D (signal_18653), .Q (signal_18654) ) ;
    buf_clk cell_13772 ( .C (clk), .D (signal_18659), .Q (signal_18660) ) ;
    buf_clk cell_13778 ( .C (clk), .D (signal_18665), .Q (signal_18666) ) ;
    buf_clk cell_13784 ( .C (clk), .D (signal_18671), .Q (signal_18672) ) ;
    buf_clk cell_13790 ( .C (clk), .D (signal_18677), .Q (signal_18678) ) ;
    buf_clk cell_13796 ( .C (clk), .D (signal_18683), .Q (signal_18684) ) ;
    buf_clk cell_13802 ( .C (clk), .D (signal_18689), .Q (signal_18690) ) ;
    buf_clk cell_13808 ( .C (clk), .D (signal_18695), .Q (signal_18696) ) ;
    buf_clk cell_13814 ( .C (clk), .D (signal_18701), .Q (signal_18702) ) ;
    buf_clk cell_13820 ( .C (clk), .D (signal_18707), .Q (signal_18708) ) ;
    buf_clk cell_13826 ( .C (clk), .D (signal_18713), .Q (signal_18714) ) ;
    buf_clk cell_13832 ( .C (clk), .D (signal_18719), .Q (signal_18720) ) ;
    buf_clk cell_13838 ( .C (clk), .D (signal_18725), .Q (signal_18726) ) ;
    buf_clk cell_13844 ( .C (clk), .D (signal_18731), .Q (signal_18732) ) ;
    buf_clk cell_13850 ( .C (clk), .D (signal_18737), .Q (signal_18738) ) ;
    buf_clk cell_13856 ( .C (clk), .D (signal_18743), .Q (signal_18744) ) ;
    buf_clk cell_13862 ( .C (clk), .D (signal_18749), .Q (signal_18750) ) ;
    buf_clk cell_13868 ( .C (clk), .D (signal_18755), .Q (signal_18756) ) ;
    buf_clk cell_13874 ( .C (clk), .D (signal_18761), .Q (signal_18762) ) ;
    buf_clk cell_13880 ( .C (clk), .D (signal_18767), .Q (signal_18768) ) ;
    buf_clk cell_13886 ( .C (clk), .D (signal_18773), .Q (signal_18774) ) ;
    buf_clk cell_13892 ( .C (clk), .D (signal_18779), .Q (signal_18780) ) ;
    buf_clk cell_13898 ( .C (clk), .D (signal_18785), .Q (signal_18786) ) ;
    buf_clk cell_13904 ( .C (clk), .D (signal_18791), .Q (signal_18792) ) ;
    buf_clk cell_13910 ( .C (clk), .D (signal_18797), .Q (signal_18798) ) ;
    buf_clk cell_13916 ( .C (clk), .D (signal_18803), .Q (signal_18804) ) ;
    buf_clk cell_13922 ( .C (clk), .D (signal_18809), .Q (signal_18810) ) ;
    buf_clk cell_13928 ( .C (clk), .D (signal_18815), .Q (signal_18816) ) ;
    buf_clk cell_13934 ( .C (clk), .D (signal_18821), .Q (signal_18822) ) ;
    buf_clk cell_13940 ( .C (clk), .D (signal_18827), .Q (signal_18828) ) ;
    buf_clk cell_13946 ( .C (clk), .D (signal_18833), .Q (signal_18834) ) ;
    buf_clk cell_13952 ( .C (clk), .D (signal_18839), .Q (signal_18840) ) ;
    buf_clk cell_13958 ( .C (clk), .D (signal_18845), .Q (signal_18846) ) ;
    buf_clk cell_13964 ( .C (clk), .D (signal_18851), .Q (signal_18852) ) ;
    buf_clk cell_13970 ( .C (clk), .D (signal_18857), .Q (signal_18858) ) ;
    buf_clk cell_13976 ( .C (clk), .D (signal_18863), .Q (signal_18864) ) ;
    buf_clk cell_13982 ( .C (clk), .D (signal_18869), .Q (signal_18870) ) ;
    buf_clk cell_13988 ( .C (clk), .D (signal_18875), .Q (signal_18876) ) ;
    buf_clk cell_13994 ( .C (clk), .D (signal_18881), .Q (signal_18882) ) ;
    buf_clk cell_14000 ( .C (clk), .D (signal_18887), .Q (signal_18888) ) ;
    buf_clk cell_14006 ( .C (clk), .D (signal_18893), .Q (signal_18894) ) ;
    buf_clk cell_14012 ( .C (clk), .D (signal_18899), .Q (signal_18900) ) ;
    buf_clk cell_14018 ( .C (clk), .D (signal_18905), .Q (signal_18906) ) ;
    buf_clk cell_14024 ( .C (clk), .D (signal_18911), .Q (signal_18912) ) ;
    buf_clk cell_14030 ( .C (clk), .D (signal_18917), .Q (signal_18918) ) ;
    buf_clk cell_14036 ( .C (clk), .D (signal_18923), .Q (signal_18924) ) ;
    buf_clk cell_14042 ( .C (clk), .D (signal_18929), .Q (signal_18930) ) ;
    buf_clk cell_14048 ( .C (clk), .D (signal_18935), .Q (signal_18936) ) ;
    buf_clk cell_14054 ( .C (clk), .D (signal_18941), .Q (signal_18942) ) ;
    buf_clk cell_14060 ( .C (clk), .D (signal_18947), .Q (signal_18948) ) ;
    buf_clk cell_14066 ( .C (clk), .D (signal_18953), .Q (signal_18954) ) ;
    buf_clk cell_14072 ( .C (clk), .D (signal_18959), .Q (signal_18960) ) ;
    buf_clk cell_14078 ( .C (clk), .D (signal_18965), .Q (signal_18966) ) ;
    buf_clk cell_14084 ( .C (clk), .D (signal_18971), .Q (signal_18972) ) ;
    buf_clk cell_14090 ( .C (clk), .D (signal_18977), .Q (signal_18978) ) ;
    buf_clk cell_14096 ( .C (clk), .D (signal_18983), .Q (signal_18984) ) ;
    buf_clk cell_14102 ( .C (clk), .D (signal_18989), .Q (signal_18990) ) ;
    buf_clk cell_14108 ( .C (clk), .D (signal_18995), .Q (signal_18996) ) ;
    buf_clk cell_14114 ( .C (clk), .D (signal_19001), .Q (signal_19002) ) ;
    buf_clk cell_14120 ( .C (clk), .D (signal_19007), .Q (signal_19008) ) ;
    buf_clk cell_14126 ( .C (clk), .D (signal_19013), .Q (signal_19014) ) ;
    buf_clk cell_14132 ( .C (clk), .D (signal_19019), .Q (signal_19020) ) ;
    buf_clk cell_14138 ( .C (clk), .D (signal_19025), .Q (signal_19026) ) ;
    buf_clk cell_14144 ( .C (clk), .D (signal_19031), .Q (signal_19032) ) ;
    buf_clk cell_14150 ( .C (clk), .D (signal_19037), .Q (signal_19038) ) ;
    buf_clk cell_14156 ( .C (clk), .D (signal_19043), .Q (signal_19044) ) ;
    buf_clk cell_14162 ( .C (clk), .D (signal_19049), .Q (signal_19050) ) ;
    buf_clk cell_14168 ( .C (clk), .D (signal_19055), .Q (signal_19056) ) ;
    buf_clk cell_14174 ( .C (clk), .D (signal_19061), .Q (signal_19062) ) ;
    buf_clk cell_14180 ( .C (clk), .D (signal_19067), .Q (signal_19068) ) ;
    buf_clk cell_14186 ( .C (clk), .D (signal_19073), .Q (signal_19074) ) ;
    buf_clk cell_14192 ( .C (clk), .D (signal_19079), .Q (signal_19080) ) ;
    buf_clk cell_14198 ( .C (clk), .D (signal_19085), .Q (signal_19086) ) ;
    buf_clk cell_14204 ( .C (clk), .D (signal_19091), .Q (signal_19092) ) ;
    buf_clk cell_14210 ( .C (clk), .D (signal_19097), .Q (signal_19098) ) ;
    buf_clk cell_14216 ( .C (clk), .D (signal_19103), .Q (signal_19104) ) ;
    buf_clk cell_14222 ( .C (clk), .D (signal_19109), .Q (signal_19110) ) ;
    buf_clk cell_14228 ( .C (clk), .D (signal_19115), .Q (signal_19116) ) ;
    buf_clk cell_14234 ( .C (clk), .D (signal_19121), .Q (signal_19122) ) ;
    buf_clk cell_14240 ( .C (clk), .D (signal_19127), .Q (signal_19128) ) ;
    buf_clk cell_14246 ( .C (clk), .D (signal_19133), .Q (signal_19134) ) ;
    buf_clk cell_14252 ( .C (clk), .D (signal_19139), .Q (signal_19140) ) ;
    buf_clk cell_14258 ( .C (clk), .D (signal_19145), .Q (signal_19146) ) ;
    buf_clk cell_14264 ( .C (clk), .D (signal_19151), .Q (signal_19152) ) ;
    buf_clk cell_14270 ( .C (clk), .D (signal_19157), .Q (signal_19158) ) ;
    buf_clk cell_14276 ( .C (clk), .D (signal_19163), .Q (signal_19164) ) ;
    buf_clk cell_14282 ( .C (clk), .D (signal_19169), .Q (signal_19170) ) ;
    buf_clk cell_14288 ( .C (clk), .D (signal_19175), .Q (signal_19176) ) ;
    buf_clk cell_14294 ( .C (clk), .D (signal_19181), .Q (signal_19182) ) ;
    buf_clk cell_14300 ( .C (clk), .D (signal_19187), .Q (signal_19188) ) ;
    buf_clk cell_14306 ( .C (clk), .D (signal_19193), .Q (signal_19194) ) ;
    buf_clk cell_14312 ( .C (clk), .D (signal_19199), .Q (signal_19200) ) ;
    buf_clk cell_14318 ( .C (clk), .D (signal_19205), .Q (signal_19206) ) ;
    buf_clk cell_14324 ( .C (clk), .D (signal_19211), .Q (signal_19212) ) ;
    buf_clk cell_14330 ( .C (clk), .D (signal_19217), .Q (signal_19218) ) ;
    buf_clk cell_14336 ( .C (clk), .D (signal_19223), .Q (signal_19224) ) ;
    buf_clk cell_14342 ( .C (clk), .D (signal_19229), .Q (signal_19230) ) ;
    buf_clk cell_14348 ( .C (clk), .D (signal_19235), .Q (signal_19236) ) ;
    buf_clk cell_14354 ( .C (clk), .D (signal_19241), .Q (signal_19242) ) ;
    buf_clk cell_14360 ( .C (clk), .D (signal_19247), .Q (signal_19248) ) ;
    buf_clk cell_14366 ( .C (clk), .D (signal_19253), .Q (signal_19254) ) ;
    buf_clk cell_14372 ( .C (clk), .D (signal_19259), .Q (signal_19260) ) ;
    buf_clk cell_14378 ( .C (clk), .D (signal_19265), .Q (signal_19266) ) ;
    buf_clk cell_14384 ( .C (clk), .D (signal_19271), .Q (signal_19272) ) ;
    buf_clk cell_14390 ( .C (clk), .D (signal_19277), .Q (signal_19278) ) ;
    buf_clk cell_14396 ( .C (clk), .D (signal_19283), .Q (signal_19284) ) ;
    buf_clk cell_14402 ( .C (clk), .D (signal_19289), .Q (signal_19290) ) ;
    buf_clk cell_14408 ( .C (clk), .D (signal_19295), .Q (signal_19296) ) ;
    buf_clk cell_14414 ( .C (clk), .D (signal_19301), .Q (signal_19302) ) ;
    buf_clk cell_14420 ( .C (clk), .D (signal_19307), .Q (signal_19308) ) ;
    buf_clk cell_14426 ( .C (clk), .D (signal_19313), .Q (signal_19314) ) ;
    buf_clk cell_14432 ( .C (clk), .D (signal_19319), .Q (signal_19320) ) ;
    buf_clk cell_14438 ( .C (clk), .D (signal_19325), .Q (signal_19326) ) ;
    buf_clk cell_14444 ( .C (clk), .D (signal_19331), .Q (signal_19332) ) ;
    buf_clk cell_14450 ( .C (clk), .D (signal_19337), .Q (signal_19338) ) ;
    buf_clk cell_14456 ( .C (clk), .D (signal_19343), .Q (signal_19344) ) ;
    buf_clk cell_14462 ( .C (clk), .D (signal_19349), .Q (signal_19350) ) ;
    buf_clk cell_14468 ( .C (clk), .D (signal_19355), .Q (signal_19356) ) ;
    buf_clk cell_14474 ( .C (clk), .D (signal_19361), .Q (signal_19362) ) ;
    buf_clk cell_14480 ( .C (clk), .D (signal_19367), .Q (signal_19368) ) ;
    buf_clk cell_14486 ( .C (clk), .D (signal_19373), .Q (signal_19374) ) ;
    buf_clk cell_14492 ( .C (clk), .D (signal_19379), .Q (signal_19380) ) ;
    buf_clk cell_14498 ( .C (clk), .D (signal_19385), .Q (signal_19386) ) ;
    buf_clk cell_14504 ( .C (clk), .D (signal_19391), .Q (signal_19392) ) ;
    buf_clk cell_14510 ( .C (clk), .D (signal_19397), .Q (signal_19398) ) ;
    buf_clk cell_14516 ( .C (clk), .D (signal_19403), .Q (signal_19404) ) ;
    buf_clk cell_14522 ( .C (clk), .D (signal_19409), .Q (signal_19410) ) ;
    buf_clk cell_14528 ( .C (clk), .D (signal_19415), .Q (signal_19416) ) ;
    buf_clk cell_14534 ( .C (clk), .D (signal_19421), .Q (signal_19422) ) ;
    buf_clk cell_14540 ( .C (clk), .D (signal_19427), .Q (signal_19428) ) ;
    buf_clk cell_14546 ( .C (clk), .D (signal_19433), .Q (signal_19434) ) ;
    buf_clk cell_14552 ( .C (clk), .D (signal_19439), .Q (signal_19440) ) ;
    buf_clk cell_14558 ( .C (clk), .D (signal_19445), .Q (signal_19446) ) ;
    buf_clk cell_14564 ( .C (clk), .D (signal_19451), .Q (signal_19452) ) ;
    buf_clk cell_14570 ( .C (clk), .D (signal_19457), .Q (signal_19458) ) ;
    buf_clk cell_14576 ( .C (clk), .D (signal_19463), .Q (signal_19464) ) ;
    buf_clk cell_14582 ( .C (clk), .D (signal_19469), .Q (signal_19470) ) ;
    buf_clk cell_14588 ( .C (clk), .D (signal_19475), .Q (signal_19476) ) ;
    buf_clk cell_14594 ( .C (clk), .D (signal_19481), .Q (signal_19482) ) ;
    buf_clk cell_14600 ( .C (clk), .D (signal_19487), .Q (signal_19488) ) ;
    buf_clk cell_14606 ( .C (clk), .D (signal_19493), .Q (signal_19494) ) ;
    buf_clk cell_14612 ( .C (clk), .D (signal_19499), .Q (signal_19500) ) ;
    buf_clk cell_14618 ( .C (clk), .D (signal_19505), .Q (signal_19506) ) ;
    buf_clk cell_14624 ( .C (clk), .D (signal_19511), .Q (signal_19512) ) ;
    buf_clk cell_14630 ( .C (clk), .D (signal_19517), .Q (signal_19518) ) ;
    buf_clk cell_14636 ( .C (clk), .D (signal_19523), .Q (signal_19524) ) ;
    buf_clk cell_14642 ( .C (clk), .D (signal_19529), .Q (signal_19530) ) ;
    buf_clk cell_14648 ( .C (clk), .D (signal_19535), .Q (signal_19536) ) ;
    buf_clk cell_14654 ( .C (clk), .D (signal_19541), .Q (signal_19542) ) ;
    buf_clk cell_14660 ( .C (clk), .D (signal_19547), .Q (signal_19548) ) ;
    buf_clk cell_14666 ( .C (clk), .D (signal_19553), .Q (signal_19554) ) ;
    buf_clk cell_14672 ( .C (clk), .D (signal_19559), .Q (signal_19560) ) ;
    buf_clk cell_14678 ( .C (clk), .D (signal_19565), .Q (signal_19566) ) ;
    buf_clk cell_14684 ( .C (clk), .D (signal_19571), .Q (signal_19572) ) ;
    buf_clk cell_14690 ( .C (clk), .D (signal_19577), .Q (signal_19578) ) ;
    buf_clk cell_14696 ( .C (clk), .D (signal_19583), .Q (signal_19584) ) ;
    buf_clk cell_14702 ( .C (clk), .D (signal_19589), .Q (signal_19590) ) ;
    buf_clk cell_14708 ( .C (clk), .D (signal_19595), .Q (signal_19596) ) ;
    buf_clk cell_14714 ( .C (clk), .D (signal_19601), .Q (signal_19602) ) ;
    buf_clk cell_14720 ( .C (clk), .D (signal_19607), .Q (signal_19608) ) ;
    buf_clk cell_14726 ( .C (clk), .D (signal_19613), .Q (signal_19614) ) ;
    buf_clk cell_14732 ( .C (clk), .D (signal_19619), .Q (signal_19620) ) ;
    buf_clk cell_14738 ( .C (clk), .D (signal_19625), .Q (signal_19626) ) ;
    buf_clk cell_14744 ( .C (clk), .D (signal_19631), .Q (signal_19632) ) ;
    buf_clk cell_14750 ( .C (clk), .D (signal_19637), .Q (signal_19638) ) ;
    buf_clk cell_14756 ( .C (clk), .D (signal_19643), .Q (signal_19644) ) ;
    buf_clk cell_14762 ( .C (clk), .D (signal_19649), .Q (signal_19650) ) ;
    buf_clk cell_14768 ( .C (clk), .D (signal_19655), .Q (signal_19656) ) ;
    buf_clk cell_14774 ( .C (clk), .D (signal_19661), .Q (signal_19662) ) ;
    buf_clk cell_14780 ( .C (clk), .D (signal_19667), .Q (signal_19668) ) ;
    buf_clk cell_14786 ( .C (clk), .D (signal_19673), .Q (signal_19674) ) ;
    buf_clk cell_14792 ( .C (clk), .D (signal_19679), .Q (signal_19680) ) ;
    buf_clk cell_14798 ( .C (clk), .D (signal_19685), .Q (signal_19686) ) ;
    buf_clk cell_14804 ( .C (clk), .D (signal_19691), .Q (signal_19692) ) ;
    buf_clk cell_14810 ( .C (clk), .D (signal_19697), .Q (signal_19698) ) ;
    buf_clk cell_14816 ( .C (clk), .D (signal_19703), .Q (signal_19704) ) ;
    buf_clk cell_14822 ( .C (clk), .D (signal_19709), .Q (signal_19710) ) ;
    buf_clk cell_14828 ( .C (clk), .D (signal_19715), .Q (signal_19716) ) ;
    buf_clk cell_14834 ( .C (clk), .D (signal_19721), .Q (signal_19722) ) ;
    buf_clk cell_14840 ( .C (clk), .D (signal_19727), .Q (signal_19728) ) ;
    buf_clk cell_14846 ( .C (clk), .D (signal_19733), .Q (signal_19734) ) ;
    buf_clk cell_14852 ( .C (clk), .D (signal_19739), .Q (signal_19740) ) ;
    buf_clk cell_14858 ( .C (clk), .D (signal_19745), .Q (signal_19746) ) ;
    buf_clk cell_14864 ( .C (clk), .D (signal_19751), .Q (signal_19752) ) ;
    buf_clk cell_14870 ( .C (clk), .D (signal_19757), .Q (signal_19758) ) ;
    buf_clk cell_14876 ( .C (clk), .D (signal_19763), .Q (signal_19764) ) ;
    buf_clk cell_14882 ( .C (clk), .D (signal_19769), .Q (signal_19770) ) ;
    buf_clk cell_14888 ( .C (clk), .D (signal_19775), .Q (signal_19776) ) ;
    buf_clk cell_14894 ( .C (clk), .D (signal_19781), .Q (signal_19782) ) ;
    buf_clk cell_14900 ( .C (clk), .D (signal_19787), .Q (signal_19788) ) ;
    buf_clk cell_14906 ( .C (clk), .D (signal_19793), .Q (signal_19794) ) ;
    buf_clk cell_14912 ( .C (clk), .D (signal_19799), .Q (signal_19800) ) ;
    buf_clk cell_14918 ( .C (clk), .D (signal_19805), .Q (signal_19806) ) ;
    buf_clk cell_14924 ( .C (clk), .D (signal_19811), .Q (signal_19812) ) ;
    buf_clk cell_14930 ( .C (clk), .D (signal_19817), .Q (signal_19818) ) ;
    buf_clk cell_14936 ( .C (clk), .D (signal_19823), .Q (signal_19824) ) ;
    buf_clk cell_14942 ( .C (clk), .D (signal_19829), .Q (signal_19830) ) ;
    buf_clk cell_14948 ( .C (clk), .D (signal_19835), .Q (signal_19836) ) ;
    buf_clk cell_14954 ( .C (clk), .D (signal_19841), .Q (signal_19842) ) ;
    buf_clk cell_14960 ( .C (clk), .D (signal_19847), .Q (signal_19848) ) ;
    buf_clk cell_14966 ( .C (clk), .D (signal_19853), .Q (signal_19854) ) ;
    buf_clk cell_14972 ( .C (clk), .D (signal_19859), .Q (signal_19860) ) ;
    buf_clk cell_14978 ( .C (clk), .D (signal_19865), .Q (signal_19866) ) ;
    buf_clk cell_14984 ( .C (clk), .D (signal_19871), .Q (signal_19872) ) ;
    buf_clk cell_14990 ( .C (clk), .D (signal_19877), .Q (signal_19878) ) ;
    buf_clk cell_14996 ( .C (clk), .D (signal_19883), .Q (signal_19884) ) ;
    buf_clk cell_15002 ( .C (clk), .D (signal_19889), .Q (signal_19890) ) ;
    buf_clk cell_15008 ( .C (clk), .D (signal_19895), .Q (signal_19896) ) ;
    buf_clk cell_15014 ( .C (clk), .D (signal_19901), .Q (signal_19902) ) ;
    buf_clk cell_15020 ( .C (clk), .D (signal_19907), .Q (signal_19908) ) ;
    buf_clk cell_15026 ( .C (clk), .D (signal_19913), .Q (signal_19914) ) ;
    buf_clk cell_15032 ( .C (clk), .D (signal_19919), .Q (signal_19920) ) ;
    buf_clk cell_15038 ( .C (clk), .D (signal_19925), .Q (signal_19926) ) ;
    buf_clk cell_15044 ( .C (clk), .D (signal_19931), .Q (signal_19932) ) ;
    buf_clk cell_15050 ( .C (clk), .D (signal_19937), .Q (signal_19938) ) ;
    buf_clk cell_15056 ( .C (clk), .D (signal_19943), .Q (signal_19944) ) ;
    buf_clk cell_15062 ( .C (clk), .D (signal_19949), .Q (signal_19950) ) ;
    buf_clk cell_15068 ( .C (clk), .D (signal_19955), .Q (signal_19956) ) ;
    buf_clk cell_15074 ( .C (clk), .D (signal_19961), .Q (signal_19962) ) ;
    buf_clk cell_15080 ( .C (clk), .D (signal_19967), .Q (signal_19968) ) ;
    buf_clk cell_15086 ( .C (clk), .D (signal_19973), .Q (signal_19974) ) ;
    buf_clk cell_15092 ( .C (clk), .D (signal_19979), .Q (signal_19980) ) ;
    buf_clk cell_15098 ( .C (clk), .D (signal_19985), .Q (signal_19986) ) ;
    buf_clk cell_15104 ( .C (clk), .D (signal_19991), .Q (signal_19992) ) ;
    buf_clk cell_15110 ( .C (clk), .D (signal_19997), .Q (signal_19998) ) ;
    buf_clk cell_15116 ( .C (clk), .D (signal_20003), .Q (signal_20004) ) ;
    buf_clk cell_15122 ( .C (clk), .D (signal_20009), .Q (signal_20010) ) ;
    buf_clk cell_15128 ( .C (clk), .D (signal_20015), .Q (signal_20016) ) ;
    buf_clk cell_15134 ( .C (clk), .D (signal_20021), .Q (signal_20022) ) ;
    buf_clk cell_15140 ( .C (clk), .D (signal_20027), .Q (signal_20028) ) ;
    buf_clk cell_15146 ( .C (clk), .D (signal_20033), .Q (signal_20034) ) ;
    buf_clk cell_15152 ( .C (clk), .D (signal_20039), .Q (signal_20040) ) ;
    buf_clk cell_15158 ( .C (clk), .D (signal_20045), .Q (signal_20046) ) ;
    buf_clk cell_15164 ( .C (clk), .D (signal_20051), .Q (signal_20052) ) ;
    buf_clk cell_15170 ( .C (clk), .D (signal_20057), .Q (signal_20058) ) ;
    buf_clk cell_15176 ( .C (clk), .D (signal_20063), .Q (signal_20064) ) ;
    buf_clk cell_15182 ( .C (clk), .D (signal_20069), .Q (signal_20070) ) ;
    buf_clk cell_15188 ( .C (clk), .D (signal_20075), .Q (signal_20076) ) ;
    buf_clk cell_15194 ( .C (clk), .D (signal_20081), .Q (signal_20082) ) ;
    buf_clk cell_15200 ( .C (clk), .D (signal_20087), .Q (signal_20088) ) ;
    buf_clk cell_15206 ( .C (clk), .D (signal_20093), .Q (signal_20094) ) ;
    buf_clk cell_15212 ( .C (clk), .D (signal_20099), .Q (signal_20100) ) ;
    buf_clk cell_15218 ( .C (clk), .D (signal_20105), .Q (signal_20106) ) ;
    buf_clk cell_15224 ( .C (clk), .D (signal_20111), .Q (signal_20112) ) ;
    buf_clk cell_15230 ( .C (clk), .D (signal_20117), .Q (signal_20118) ) ;
    buf_clk cell_15236 ( .C (clk), .D (signal_20123), .Q (signal_20124) ) ;
    buf_clk cell_15242 ( .C (clk), .D (signal_20129), .Q (signal_20130) ) ;
    buf_clk cell_15248 ( .C (clk), .D (signal_20135), .Q (signal_20136) ) ;
    buf_clk cell_15254 ( .C (clk), .D (signal_20141), .Q (signal_20142) ) ;
    buf_clk cell_15260 ( .C (clk), .D (signal_20147), .Q (signal_20148) ) ;
    buf_clk cell_15266 ( .C (clk), .D (signal_20153), .Q (signal_20154) ) ;
    buf_clk cell_15272 ( .C (clk), .D (signal_20159), .Q (signal_20160) ) ;
    buf_clk cell_15278 ( .C (clk), .D (signal_20165), .Q (signal_20166) ) ;
    buf_clk cell_15284 ( .C (clk), .D (signal_20171), .Q (signal_20172) ) ;
    buf_clk cell_15290 ( .C (clk), .D (signal_20177), .Q (signal_20178) ) ;
    buf_clk cell_15296 ( .C (clk), .D (signal_20183), .Q (signal_20184) ) ;
    buf_clk cell_15302 ( .C (clk), .D (signal_20189), .Q (signal_20190) ) ;
    buf_clk cell_15308 ( .C (clk), .D (signal_20195), .Q (signal_20196) ) ;
    buf_clk cell_15314 ( .C (clk), .D (signal_20201), .Q (signal_20202) ) ;
    buf_clk cell_15320 ( .C (clk), .D (signal_20207), .Q (signal_20208) ) ;
    buf_clk cell_15326 ( .C (clk), .D (signal_20213), .Q (signal_20214) ) ;
    buf_clk cell_15332 ( .C (clk), .D (signal_20219), .Q (signal_20220) ) ;
    buf_clk cell_15338 ( .C (clk), .D (signal_20225), .Q (signal_20226) ) ;
    buf_clk cell_15344 ( .C (clk), .D (signal_20231), .Q (signal_20232) ) ;
    buf_clk cell_15350 ( .C (clk), .D (signal_20237), .Q (signal_20238) ) ;
    buf_clk cell_15356 ( .C (clk), .D (signal_20243), .Q (signal_20244) ) ;
    buf_clk cell_15362 ( .C (clk), .D (signal_20249), .Q (signal_20250) ) ;
    buf_clk cell_15368 ( .C (clk), .D (signal_20255), .Q (signal_20256) ) ;
    buf_clk cell_15374 ( .C (clk), .D (signal_20261), .Q (signal_20262) ) ;
    buf_clk cell_15380 ( .C (clk), .D (signal_20267), .Q (signal_20268) ) ;
    buf_clk cell_15386 ( .C (clk), .D (signal_20273), .Q (signal_20274) ) ;
    buf_clk cell_15392 ( .C (clk), .D (signal_20279), .Q (signal_20280) ) ;
    buf_clk cell_15398 ( .C (clk), .D (signal_20285), .Q (signal_20286) ) ;
    buf_clk cell_15404 ( .C (clk), .D (signal_20291), .Q (signal_20292) ) ;
    buf_clk cell_15410 ( .C (clk), .D (signal_20297), .Q (signal_20298) ) ;
    buf_clk cell_15416 ( .C (clk), .D (signal_20303), .Q (signal_20304) ) ;
    buf_clk cell_15422 ( .C (clk), .D (signal_20309), .Q (signal_20310) ) ;
    buf_clk cell_15428 ( .C (clk), .D (signal_20315), .Q (signal_20316) ) ;
    buf_clk cell_15434 ( .C (clk), .D (signal_20321), .Q (signal_20322) ) ;
    buf_clk cell_15440 ( .C (clk), .D (signal_20327), .Q (signal_20328) ) ;
    buf_clk cell_15446 ( .C (clk), .D (signal_20333), .Q (signal_20334) ) ;
    buf_clk cell_15452 ( .C (clk), .D (signal_20339), .Q (signal_20340) ) ;
    buf_clk cell_15458 ( .C (clk), .D (signal_20345), .Q (signal_20346) ) ;
    buf_clk cell_15464 ( .C (clk), .D (signal_20351), .Q (signal_20352) ) ;
    buf_clk cell_15470 ( .C (clk), .D (signal_20357), .Q (signal_20358) ) ;
    buf_clk cell_15476 ( .C (clk), .D (signal_20363), .Q (signal_20364) ) ;
    buf_clk cell_15482 ( .C (clk), .D (signal_20369), .Q (signal_20370) ) ;
    buf_clk cell_15488 ( .C (clk), .D (signal_20375), .Q (signal_20376) ) ;
    buf_clk cell_15494 ( .C (clk), .D (signal_20381), .Q (signal_20382) ) ;
    buf_clk cell_15500 ( .C (clk), .D (signal_20387), .Q (signal_20388) ) ;
    buf_clk cell_15506 ( .C (clk), .D (signal_20393), .Q (signal_20394) ) ;
    buf_clk cell_15512 ( .C (clk), .D (signal_20399), .Q (signal_20400) ) ;
    buf_clk cell_15518 ( .C (clk), .D (signal_20405), .Q (signal_20406) ) ;
    buf_clk cell_15524 ( .C (clk), .D (signal_20411), .Q (signal_20412) ) ;
    buf_clk cell_15530 ( .C (clk), .D (signal_20417), .Q (signal_20418) ) ;
    buf_clk cell_15536 ( .C (clk), .D (signal_20423), .Q (signal_20424) ) ;
    buf_clk cell_15542 ( .C (clk), .D (signal_20429), .Q (signal_20430) ) ;
    buf_clk cell_15548 ( .C (clk), .D (signal_20435), .Q (signal_20436) ) ;
    buf_clk cell_15554 ( .C (clk), .D (signal_20441), .Q (signal_20442) ) ;
    buf_clk cell_15560 ( .C (clk), .D (signal_20447), .Q (signal_20448) ) ;
    buf_clk cell_15566 ( .C (clk), .D (signal_20453), .Q (signal_20454) ) ;
    buf_clk cell_15572 ( .C (clk), .D (signal_20459), .Q (signal_20460) ) ;
    buf_clk cell_15578 ( .C (clk), .D (signal_20465), .Q (signal_20466) ) ;
    buf_clk cell_15584 ( .C (clk), .D (signal_20471), .Q (signal_20472) ) ;
    buf_clk cell_15590 ( .C (clk), .D (signal_20477), .Q (signal_20478) ) ;
    buf_clk cell_15596 ( .C (clk), .D (signal_20483), .Q (signal_20484) ) ;
    buf_clk cell_15602 ( .C (clk), .D (signal_20489), .Q (signal_20490) ) ;
    buf_clk cell_15608 ( .C (clk), .D (signal_20495), .Q (signal_20496) ) ;
    buf_clk cell_15614 ( .C (clk), .D (signal_20501), .Q (signal_20502) ) ;
    buf_clk cell_15620 ( .C (clk), .D (signal_20507), .Q (signal_20508) ) ;
    buf_clk cell_15626 ( .C (clk), .D (signal_20513), .Q (signal_20514) ) ;
    buf_clk cell_15632 ( .C (clk), .D (signal_20519), .Q (signal_20520) ) ;
    buf_clk cell_15638 ( .C (clk), .D (signal_20525), .Q (signal_20526) ) ;
    buf_clk cell_15644 ( .C (clk), .D (signal_20531), .Q (signal_20532) ) ;
    buf_clk cell_15650 ( .C (clk), .D (signal_20537), .Q (signal_20538) ) ;
    buf_clk cell_15656 ( .C (clk), .D (signal_20543), .Q (signal_20544) ) ;
    buf_clk cell_15662 ( .C (clk), .D (signal_20549), .Q (signal_20550) ) ;
    buf_clk cell_15668 ( .C (clk), .D (signal_20555), .Q (signal_20556) ) ;
    buf_clk cell_15674 ( .C (clk), .D (signal_20561), .Q (signal_20562) ) ;
    buf_clk cell_15680 ( .C (clk), .D (signal_20567), .Q (signal_20568) ) ;
    buf_clk cell_15686 ( .C (clk), .D (signal_20573), .Q (signal_20574) ) ;
    buf_clk cell_15692 ( .C (clk), .D (signal_20579), .Q (signal_20580) ) ;
    buf_clk cell_15698 ( .C (clk), .D (signal_20585), .Q (signal_20586) ) ;
    buf_clk cell_15704 ( .C (clk), .D (signal_20591), .Q (signal_20592) ) ;
    buf_clk cell_15710 ( .C (clk), .D (signal_20597), .Q (signal_20598) ) ;
    buf_clk cell_15716 ( .C (clk), .D (signal_20603), .Q (signal_20604) ) ;
    buf_clk cell_15722 ( .C (clk), .D (signal_20609), .Q (signal_20610) ) ;
    buf_clk cell_15728 ( .C (clk), .D (signal_20615), .Q (signal_20616) ) ;
    buf_clk cell_15734 ( .C (clk), .D (signal_20621), .Q (signal_20622) ) ;
    buf_clk cell_15740 ( .C (clk), .D (signal_20627), .Q (signal_20628) ) ;
    buf_clk cell_15746 ( .C (clk), .D (signal_20633), .Q (signal_20634) ) ;
    buf_clk cell_15752 ( .C (clk), .D (signal_20639), .Q (signal_20640) ) ;
    buf_clk cell_15758 ( .C (clk), .D (signal_20645), .Q (signal_20646) ) ;
    buf_clk cell_15764 ( .C (clk), .D (signal_20651), .Q (signal_20652) ) ;
    buf_clk cell_15770 ( .C (clk), .D (signal_20657), .Q (signal_20658) ) ;
    buf_clk cell_15776 ( .C (clk), .D (signal_20663), .Q (signal_20664) ) ;
    buf_clk cell_15782 ( .C (clk), .D (signal_20669), .Q (signal_20670) ) ;
    buf_clk cell_15788 ( .C (clk), .D (signal_20675), .Q (signal_20676) ) ;
    buf_clk cell_15794 ( .C (clk), .D (signal_20681), .Q (signal_20682) ) ;
    buf_clk cell_15800 ( .C (clk), .D (signal_20687), .Q (signal_20688) ) ;
    buf_clk cell_15806 ( .C (clk), .D (signal_20693), .Q (signal_20694) ) ;
    buf_clk cell_15812 ( .C (clk), .D (signal_20699), .Q (signal_20700) ) ;
    buf_clk cell_15818 ( .C (clk), .D (signal_20705), .Q (signal_20706) ) ;
    buf_clk cell_15824 ( .C (clk), .D (signal_20711), .Q (signal_20712) ) ;
    buf_clk cell_15830 ( .C (clk), .D (signal_20717), .Q (signal_20718) ) ;
    buf_clk cell_15836 ( .C (clk), .D (signal_20723), .Q (signal_20724) ) ;
    buf_clk cell_15842 ( .C (clk), .D (signal_20729), .Q (signal_20730) ) ;
    buf_clk cell_15848 ( .C (clk), .D (signal_20735), .Q (signal_20736) ) ;
    buf_clk cell_15854 ( .C (clk), .D (signal_20741), .Q (signal_20742) ) ;
    buf_clk cell_15860 ( .C (clk), .D (signal_20747), .Q (signal_20748) ) ;
    buf_clk cell_15866 ( .C (clk), .D (signal_20753), .Q (signal_20754) ) ;
    buf_clk cell_15872 ( .C (clk), .D (signal_20759), .Q (signal_20760) ) ;
    buf_clk cell_15878 ( .C (clk), .D (signal_20765), .Q (signal_20766) ) ;
    buf_clk cell_15884 ( .C (clk), .D (signal_20771), .Q (signal_20772) ) ;
    buf_clk cell_15890 ( .C (clk), .D (signal_20777), .Q (signal_20778) ) ;
    buf_clk cell_15896 ( .C (clk), .D (signal_20783), .Q (signal_20784) ) ;
    buf_clk cell_15902 ( .C (clk), .D (signal_20789), .Q (signal_20790) ) ;
    buf_clk cell_15908 ( .C (clk), .D (signal_20795), .Q (signal_20796) ) ;
    buf_clk cell_15914 ( .C (clk), .D (signal_20801), .Q (signal_20802) ) ;
    buf_clk cell_15920 ( .C (clk), .D (signal_20807), .Q (signal_20808) ) ;
    buf_clk cell_15926 ( .C (clk), .D (signal_20813), .Q (signal_20814) ) ;
    buf_clk cell_15932 ( .C (clk), .D (signal_20819), .Q (signal_20820) ) ;
    buf_clk cell_15938 ( .C (clk), .D (signal_20825), .Q (signal_20826) ) ;
    buf_clk cell_15944 ( .C (clk), .D (signal_20831), .Q (signal_20832) ) ;
    buf_clk cell_15950 ( .C (clk), .D (signal_20837), .Q (signal_20838) ) ;
    buf_clk cell_15956 ( .C (clk), .D (signal_20843), .Q (signal_20844) ) ;
    buf_clk cell_15962 ( .C (clk), .D (signal_20849), .Q (signal_20850) ) ;
    buf_clk cell_15968 ( .C (clk), .D (signal_20855), .Q (signal_20856) ) ;
    buf_clk cell_15974 ( .C (clk), .D (signal_20861), .Q (signal_20862) ) ;
    buf_clk cell_15980 ( .C (clk), .D (signal_20867), .Q (signal_20868) ) ;
    buf_clk cell_15986 ( .C (clk), .D (signal_20873), .Q (signal_20874) ) ;
    buf_clk cell_15992 ( .C (clk), .D (signal_20879), .Q (signal_20880) ) ;
    buf_clk cell_15998 ( .C (clk), .D (signal_20885), .Q (signal_20886) ) ;
    buf_clk cell_16004 ( .C (clk), .D (signal_20891), .Q (signal_20892) ) ;
    buf_clk cell_16010 ( .C (clk), .D (signal_20897), .Q (signal_20898) ) ;
    buf_clk cell_16016 ( .C (clk), .D (signal_20903), .Q (signal_20904) ) ;
    buf_clk cell_16022 ( .C (clk), .D (signal_20909), .Q (signal_20910) ) ;
    buf_clk cell_16028 ( .C (clk), .D (signal_20915), .Q (signal_20916) ) ;
    buf_clk cell_16034 ( .C (clk), .D (signal_20921), .Q (signal_20922) ) ;
    buf_clk cell_16040 ( .C (clk), .D (signal_20927), .Q (signal_20928) ) ;
    buf_clk cell_16046 ( .C (clk), .D (signal_20933), .Q (signal_20934) ) ;
    buf_clk cell_16052 ( .C (clk), .D (signal_20939), .Q (signal_20940) ) ;
    buf_clk cell_16058 ( .C (clk), .D (signal_20945), .Q (signal_20946) ) ;
    buf_clk cell_16064 ( .C (clk), .D (signal_20951), .Q (signal_20952) ) ;
    buf_clk cell_16070 ( .C (clk), .D (signal_20957), .Q (signal_20958) ) ;
    buf_clk cell_16076 ( .C (clk), .D (signal_20963), .Q (signal_20964) ) ;
    buf_clk cell_16082 ( .C (clk), .D (signal_20969), .Q (signal_20970) ) ;
    buf_clk cell_16088 ( .C (clk), .D (signal_20975), .Q (signal_20976) ) ;
    buf_clk cell_16094 ( .C (clk), .D (signal_20981), .Q (signal_20982) ) ;
    buf_clk cell_16100 ( .C (clk), .D (signal_20987), .Q (signal_20988) ) ;
    buf_clk cell_16106 ( .C (clk), .D (signal_20993), .Q (signal_20994) ) ;
    buf_clk cell_16112 ( .C (clk), .D (signal_20999), .Q (signal_21000) ) ;
    buf_clk cell_16118 ( .C (clk), .D (signal_21005), .Q (signal_21006) ) ;
    buf_clk cell_16124 ( .C (clk), .D (signal_21011), .Q (signal_21012) ) ;
    buf_clk cell_16130 ( .C (clk), .D (signal_21017), .Q (signal_21018) ) ;
    buf_clk cell_16136 ( .C (clk), .D (signal_21023), .Q (signal_21024) ) ;
    buf_clk cell_16142 ( .C (clk), .D (signal_21029), .Q (signal_21030) ) ;
    buf_clk cell_16148 ( .C (clk), .D (signal_21035), .Q (signal_21036) ) ;
    buf_clk cell_16154 ( .C (clk), .D (signal_21041), .Q (signal_21042) ) ;
    buf_clk cell_16160 ( .C (clk), .D (signal_21047), .Q (signal_21048) ) ;
    buf_clk cell_16166 ( .C (clk), .D (signal_21053), .Q (signal_21054) ) ;
    buf_clk cell_16172 ( .C (clk), .D (signal_21059), .Q (signal_21060) ) ;
    buf_clk cell_16178 ( .C (clk), .D (signal_21065), .Q (signal_21066) ) ;
    buf_clk cell_16184 ( .C (clk), .D (signal_21071), .Q (signal_21072) ) ;
    buf_clk cell_16190 ( .C (clk), .D (signal_21077), .Q (signal_21078) ) ;
    buf_clk cell_16196 ( .C (clk), .D (signal_21083), .Q (signal_21084) ) ;
    buf_clk cell_16202 ( .C (clk), .D (signal_21089), .Q (signal_21090) ) ;
    buf_clk cell_16208 ( .C (clk), .D (signal_21095), .Q (signal_21096) ) ;
    buf_clk cell_16214 ( .C (clk), .D (signal_21101), .Q (signal_21102) ) ;
    buf_clk cell_16220 ( .C (clk), .D (signal_21107), .Q (signal_21108) ) ;
    buf_clk cell_16226 ( .C (clk), .D (signal_21113), .Q (signal_21114) ) ;
    buf_clk cell_16232 ( .C (clk), .D (signal_21119), .Q (signal_21120) ) ;
    buf_clk cell_16238 ( .C (clk), .D (signal_21125), .Q (signal_21126) ) ;
    buf_clk cell_16244 ( .C (clk), .D (signal_21131), .Q (signal_21132) ) ;
    buf_clk cell_16250 ( .C (clk), .D (signal_21137), .Q (signal_21138) ) ;
    buf_clk cell_16256 ( .C (clk), .D (signal_21143), .Q (signal_21144) ) ;
    buf_clk cell_16262 ( .C (clk), .D (signal_21149), .Q (signal_21150) ) ;
    buf_clk cell_16268 ( .C (clk), .D (signal_21155), .Q (signal_21156) ) ;
    buf_clk cell_16274 ( .C (clk), .D (signal_21161), .Q (signal_21162) ) ;
    buf_clk cell_16280 ( .C (clk), .D (signal_21167), .Q (signal_21168) ) ;
    buf_clk cell_16286 ( .C (clk), .D (signal_21173), .Q (signal_21174) ) ;
    buf_clk cell_16292 ( .C (clk), .D (signal_21179), .Q (signal_21180) ) ;
    buf_clk cell_16298 ( .C (clk), .D (signal_21185), .Q (signal_21186) ) ;
    buf_clk cell_16304 ( .C (clk), .D (signal_21191), .Q (signal_21192) ) ;
    buf_clk cell_16310 ( .C (clk), .D (signal_21197), .Q (signal_21198) ) ;
    buf_clk cell_16316 ( .C (clk), .D (signal_21203), .Q (signal_21204) ) ;
    buf_clk cell_16322 ( .C (clk), .D (signal_21209), .Q (signal_21210) ) ;
    buf_clk cell_16328 ( .C (clk), .D (signal_21215), .Q (signal_21216) ) ;
    buf_clk cell_16334 ( .C (clk), .D (signal_21221), .Q (signal_21222) ) ;
    buf_clk cell_16340 ( .C (clk), .D (signal_21227), .Q (signal_21228) ) ;
    buf_clk cell_16346 ( .C (clk), .D (signal_21233), .Q (signal_21234) ) ;
    buf_clk cell_16352 ( .C (clk), .D (signal_21239), .Q (signal_21240) ) ;
    buf_clk cell_16358 ( .C (clk), .D (signal_21245), .Q (signal_21246) ) ;
    buf_clk cell_16364 ( .C (clk), .D (signal_21251), .Q (signal_21252) ) ;
    buf_clk cell_16370 ( .C (clk), .D (signal_21257), .Q (signal_21258) ) ;
    buf_clk cell_16376 ( .C (clk), .D (signal_21263), .Q (signal_21264) ) ;
    buf_clk cell_16382 ( .C (clk), .D (signal_21269), .Q (signal_21270) ) ;
    buf_clk cell_16388 ( .C (clk), .D (signal_21275), .Q (signal_21276) ) ;
    buf_clk cell_16394 ( .C (clk), .D (signal_21281), .Q (signal_21282) ) ;
    buf_clk cell_16400 ( .C (clk), .D (signal_21287), .Q (signal_21288) ) ;
    buf_clk cell_16406 ( .C (clk), .D (signal_21293), .Q (signal_21294) ) ;
    buf_clk cell_16412 ( .C (clk), .D (signal_21299), .Q (signal_21300) ) ;
    buf_clk cell_16418 ( .C (clk), .D (signal_21305), .Q (signal_21306) ) ;
    buf_clk cell_16424 ( .C (clk), .D (signal_21311), .Q (signal_21312) ) ;
    buf_clk cell_16430 ( .C (clk), .D (signal_21317), .Q (signal_21318) ) ;
    buf_clk cell_16436 ( .C (clk), .D (signal_21323), .Q (signal_21324) ) ;
    buf_clk cell_16442 ( .C (clk), .D (signal_21329), .Q (signal_21330) ) ;
    buf_clk cell_16448 ( .C (clk), .D (signal_21335), .Q (signal_21336) ) ;
    buf_clk cell_16454 ( .C (clk), .D (signal_21341), .Q (signal_21342) ) ;
    buf_clk cell_16460 ( .C (clk), .D (signal_21347), .Q (signal_21348) ) ;
    buf_clk cell_16466 ( .C (clk), .D (signal_21353), .Q (signal_21354) ) ;
    buf_clk cell_16472 ( .C (clk), .D (signal_21359), .Q (signal_21360) ) ;
    buf_clk cell_16478 ( .C (clk), .D (signal_21365), .Q (signal_21366) ) ;
    buf_clk cell_16484 ( .C (clk), .D (signal_21371), .Q (signal_21372) ) ;
    buf_clk cell_16490 ( .C (clk), .D (signal_21377), .Q (signal_21378) ) ;
    buf_clk cell_16496 ( .C (clk), .D (signal_21383), .Q (signal_21384) ) ;
    buf_clk cell_16502 ( .C (clk), .D (signal_21389), .Q (signal_21390) ) ;
    buf_clk cell_16508 ( .C (clk), .D (signal_21395), .Q (signal_21396) ) ;
    buf_clk cell_16514 ( .C (clk), .D (signal_21401), .Q (signal_21402) ) ;
    buf_clk cell_16520 ( .C (clk), .D (signal_21407), .Q (signal_21408) ) ;
    buf_clk cell_16526 ( .C (clk), .D (signal_21413), .Q (signal_21414) ) ;
    buf_clk cell_16532 ( .C (clk), .D (signal_21419), .Q (signal_21420) ) ;
    buf_clk cell_16538 ( .C (clk), .D (signal_21425), .Q (signal_21426) ) ;
    buf_clk cell_16544 ( .C (clk), .D (signal_21431), .Q (signal_21432) ) ;
    buf_clk cell_16550 ( .C (clk), .D (signal_21437), .Q (signal_21438) ) ;
    buf_clk cell_16556 ( .C (clk), .D (signal_21443), .Q (signal_21444) ) ;
    buf_clk cell_16562 ( .C (clk), .D (signal_21449), .Q (signal_21450) ) ;
    buf_clk cell_16568 ( .C (clk), .D (signal_21455), .Q (signal_21456) ) ;
    buf_clk cell_16574 ( .C (clk), .D (signal_21461), .Q (signal_21462) ) ;
    buf_clk cell_16580 ( .C (clk), .D (signal_21467), .Q (signal_21468) ) ;
    buf_clk cell_16586 ( .C (clk), .D (signal_21473), .Q (signal_21474) ) ;
    buf_clk cell_16592 ( .C (clk), .D (signal_21479), .Q (signal_21480) ) ;
    buf_clk cell_16598 ( .C (clk), .D (signal_21485), .Q (signal_21486) ) ;
    buf_clk cell_16604 ( .C (clk), .D (signal_21491), .Q (signal_21492) ) ;
    buf_clk cell_16610 ( .C (clk), .D (signal_21497), .Q (signal_21498) ) ;
    buf_clk cell_16616 ( .C (clk), .D (signal_21503), .Q (signal_21504) ) ;
    buf_clk cell_16622 ( .C (clk), .D (signal_21509), .Q (signal_21510) ) ;
    buf_clk cell_16628 ( .C (clk), .D (signal_21515), .Q (signal_21516) ) ;
    buf_clk cell_16634 ( .C (clk), .D (signal_21521), .Q (signal_21522) ) ;
    buf_clk cell_16640 ( .C (clk), .D (signal_21527), .Q (signal_21528) ) ;
    buf_clk cell_16646 ( .C (clk), .D (signal_21533), .Q (signal_21534) ) ;
    buf_clk cell_16652 ( .C (clk), .D (signal_21539), .Q (signal_21540) ) ;
    buf_clk cell_16658 ( .C (clk), .D (signal_21545), .Q (signal_21546) ) ;
    buf_clk cell_16664 ( .C (clk), .D (signal_21551), .Q (signal_21552) ) ;
    buf_clk cell_16670 ( .C (clk), .D (signal_21557), .Q (signal_21558) ) ;
    buf_clk cell_16676 ( .C (clk), .D (signal_21563), .Q (signal_21564) ) ;
    buf_clk cell_16682 ( .C (clk), .D (signal_21569), .Q (signal_21570) ) ;
    buf_clk cell_16688 ( .C (clk), .D (signal_21575), .Q (signal_21576) ) ;
    buf_clk cell_16694 ( .C (clk), .D (signal_21581), .Q (signal_21582) ) ;
    buf_clk cell_16700 ( .C (clk), .D (signal_21587), .Q (signal_21588) ) ;
    buf_clk cell_16706 ( .C (clk), .D (signal_21593), .Q (signal_21594) ) ;
    buf_clk cell_16712 ( .C (clk), .D (signal_21599), .Q (signal_21600) ) ;
    buf_clk cell_16718 ( .C (clk), .D (signal_21605), .Q (signal_21606) ) ;
    buf_clk cell_16724 ( .C (clk), .D (signal_21611), .Q (signal_21612) ) ;
    buf_clk cell_16730 ( .C (clk), .D (signal_21617), .Q (signal_21618) ) ;
    buf_clk cell_16736 ( .C (clk), .D (signal_21623), .Q (signal_21624) ) ;
    buf_clk cell_16742 ( .C (clk), .D (signal_21629), .Q (signal_21630) ) ;
    buf_clk cell_16748 ( .C (clk), .D (signal_21635), .Q (signal_21636) ) ;
    buf_clk cell_16754 ( .C (clk), .D (signal_21641), .Q (signal_21642) ) ;
    buf_clk cell_16760 ( .C (clk), .D (signal_21647), .Q (signal_21648) ) ;
    buf_clk cell_16766 ( .C (clk), .D (signal_21653), .Q (signal_21654) ) ;
    buf_clk cell_16772 ( .C (clk), .D (signal_21659), .Q (signal_21660) ) ;
    buf_clk cell_16778 ( .C (clk), .D (signal_21665), .Q (signal_21666) ) ;
    buf_clk cell_16784 ( .C (clk), .D (signal_21671), .Q (signal_21672) ) ;
    buf_clk cell_16790 ( .C (clk), .D (signal_21677), .Q (signal_21678) ) ;
    buf_clk cell_16796 ( .C (clk), .D (signal_21683), .Q (signal_21684) ) ;
    buf_clk cell_16802 ( .C (clk), .D (signal_21689), .Q (signal_21690) ) ;
    buf_clk cell_16808 ( .C (clk), .D (signal_21695), .Q (signal_21696) ) ;
    buf_clk cell_16814 ( .C (clk), .D (signal_21701), .Q (signal_21702) ) ;
    buf_clk cell_16820 ( .C (clk), .D (signal_21707), .Q (signal_21708) ) ;
    buf_clk cell_16826 ( .C (clk), .D (signal_21713), .Q (signal_21714) ) ;
    buf_clk cell_16832 ( .C (clk), .D (signal_21719), .Q (signal_21720) ) ;
    buf_clk cell_16838 ( .C (clk), .D (signal_21725), .Q (signal_21726) ) ;
    buf_clk cell_16844 ( .C (clk), .D (signal_21731), .Q (signal_21732) ) ;
    buf_clk cell_16850 ( .C (clk), .D (signal_21737), .Q (signal_21738) ) ;
    buf_clk cell_16856 ( .C (clk), .D (signal_21743), .Q (signal_21744) ) ;
    buf_clk cell_16862 ( .C (clk), .D (signal_21749), .Q (signal_21750) ) ;
    buf_clk cell_16868 ( .C (clk), .D (signal_21755), .Q (signal_21756) ) ;
    buf_clk cell_16874 ( .C (clk), .D (signal_21761), .Q (signal_21762) ) ;
    buf_clk cell_16880 ( .C (clk), .D (signal_21767), .Q (signal_21768) ) ;
    buf_clk cell_16886 ( .C (clk), .D (signal_21773), .Q (signal_21774) ) ;
    buf_clk cell_16892 ( .C (clk), .D (signal_21779), .Q (signal_21780) ) ;
    buf_clk cell_16898 ( .C (clk), .D (signal_21785), .Q (signal_21786) ) ;
    buf_clk cell_16904 ( .C (clk), .D (signal_21791), .Q (signal_21792) ) ;
    buf_clk cell_16910 ( .C (clk), .D (signal_21797), .Q (signal_21798) ) ;
    buf_clk cell_16916 ( .C (clk), .D (signal_21803), .Q (signal_21804) ) ;
    buf_clk cell_16922 ( .C (clk), .D (signal_21809), .Q (signal_21810) ) ;
    buf_clk cell_16928 ( .C (clk), .D (signal_21815), .Q (signal_21816) ) ;
    buf_clk cell_16934 ( .C (clk), .D (signal_21821), .Q (signal_21822) ) ;
    buf_clk cell_16940 ( .C (clk), .D (signal_21827), .Q (signal_21828) ) ;
    buf_clk cell_16946 ( .C (clk), .D (signal_21833), .Q (signal_21834) ) ;
    buf_clk cell_16952 ( .C (clk), .D (signal_21839), .Q (signal_21840) ) ;
    buf_clk cell_16958 ( .C (clk), .D (signal_21845), .Q (signal_21846) ) ;
    buf_clk cell_16964 ( .C (clk), .D (signal_21851), .Q (signal_21852) ) ;
    buf_clk cell_16970 ( .C (clk), .D (signal_21857), .Q (signal_21858) ) ;
    buf_clk cell_16976 ( .C (clk), .D (signal_21863), .Q (signal_21864) ) ;
    buf_clk cell_16982 ( .C (clk), .D (signal_21869), .Q (signal_21870) ) ;
    buf_clk cell_16988 ( .C (clk), .D (signal_21875), .Q (signal_21876) ) ;
    buf_clk cell_16994 ( .C (clk), .D (signal_21881), .Q (signal_21882) ) ;
    buf_clk cell_17000 ( .C (clk), .D (signal_21887), .Q (signal_21888) ) ;
    buf_clk cell_17006 ( .C (clk), .D (signal_21893), .Q (signal_21894) ) ;
    buf_clk cell_17012 ( .C (clk), .D (signal_21899), .Q (signal_21900) ) ;
    buf_clk cell_17018 ( .C (clk), .D (signal_21905), .Q (signal_21906) ) ;
    buf_clk cell_17024 ( .C (clk), .D (signal_21911), .Q (signal_21912) ) ;
    buf_clk cell_17030 ( .C (clk), .D (signal_21917), .Q (signal_21918) ) ;
    buf_clk cell_17036 ( .C (clk), .D (signal_21923), .Q (signal_21924) ) ;
    buf_clk cell_17042 ( .C (clk), .D (signal_21929), .Q (signal_21930) ) ;
    buf_clk cell_17048 ( .C (clk), .D (signal_21935), .Q (signal_21936) ) ;
    buf_clk cell_17054 ( .C (clk), .D (signal_21941), .Q (signal_21942) ) ;
    buf_clk cell_17060 ( .C (clk), .D (signal_21947), .Q (signal_21948) ) ;
    buf_clk cell_17066 ( .C (clk), .D (signal_21953), .Q (signal_21954) ) ;
    buf_clk cell_17072 ( .C (clk), .D (signal_21959), .Q (signal_21960) ) ;
    buf_clk cell_17078 ( .C (clk), .D (signal_21965), .Q (signal_21966) ) ;
    buf_clk cell_17084 ( .C (clk), .D (signal_21971), .Q (signal_21972) ) ;
    buf_clk cell_17090 ( .C (clk), .D (signal_21977), .Q (signal_21978) ) ;
    buf_clk cell_17096 ( .C (clk), .D (signal_21983), .Q (signal_21984) ) ;
    buf_clk cell_17102 ( .C (clk), .D (signal_21989), .Q (signal_21990) ) ;
    buf_clk cell_17108 ( .C (clk), .D (signal_21995), .Q (signal_21996) ) ;
    buf_clk cell_17114 ( .C (clk), .D (signal_22001), .Q (signal_22002) ) ;
    buf_clk cell_17120 ( .C (clk), .D (signal_22007), .Q (signal_22008) ) ;
    buf_clk cell_17126 ( .C (clk), .D (signal_22013), .Q (signal_22014) ) ;
    buf_clk cell_17132 ( .C (clk), .D (signal_22019), .Q (signal_22020) ) ;
    buf_clk cell_17138 ( .C (clk), .D (signal_22025), .Q (signal_22026) ) ;
    buf_clk cell_17144 ( .C (clk), .D (signal_22031), .Q (signal_22032) ) ;
    buf_clk cell_17150 ( .C (clk), .D (signal_22037), .Q (signal_22038) ) ;
    buf_clk cell_17156 ( .C (clk), .D (signal_22043), .Q (signal_22044) ) ;
    buf_clk cell_17162 ( .C (clk), .D (signal_22049), .Q (signal_22050) ) ;
    buf_clk cell_17168 ( .C (clk), .D (signal_22055), .Q (signal_22056) ) ;
    buf_clk cell_17174 ( .C (clk), .D (signal_22061), .Q (signal_22062) ) ;
    buf_clk cell_17180 ( .C (clk), .D (signal_22067), .Q (signal_22068) ) ;
    buf_clk cell_17186 ( .C (clk), .D (signal_22073), .Q (signal_22074) ) ;
    buf_clk cell_17192 ( .C (clk), .D (signal_22079), .Q (signal_22080) ) ;
    buf_clk cell_17198 ( .C (clk), .D (signal_22085), .Q (signal_22086) ) ;
    buf_clk cell_17204 ( .C (clk), .D (signal_22091), .Q (signal_22092) ) ;
    buf_clk cell_17210 ( .C (clk), .D (signal_22097), .Q (signal_22098) ) ;
    buf_clk cell_17216 ( .C (clk), .D (signal_22103), .Q (signal_22104) ) ;
    buf_clk cell_17222 ( .C (clk), .D (signal_22109), .Q (signal_22110) ) ;
    buf_clk cell_17228 ( .C (clk), .D (signal_22115), .Q (signal_22116) ) ;
    buf_clk cell_17234 ( .C (clk), .D (signal_22121), .Q (signal_22122) ) ;
    buf_clk cell_17240 ( .C (clk), .D (signal_22127), .Q (signal_22128) ) ;
    buf_clk cell_17246 ( .C (clk), .D (signal_22133), .Q (signal_22134) ) ;
    buf_clk cell_17252 ( .C (clk), .D (signal_22139), .Q (signal_22140) ) ;
    buf_clk cell_17258 ( .C (clk), .D (signal_22145), .Q (signal_22146) ) ;
    buf_clk cell_17264 ( .C (clk), .D (signal_22151), .Q (signal_22152) ) ;
    buf_clk cell_17270 ( .C (clk), .D (signal_22157), .Q (signal_22158) ) ;
    buf_clk cell_17276 ( .C (clk), .D (signal_22163), .Q (signal_22164) ) ;
    buf_clk cell_17282 ( .C (clk), .D (signal_22169), .Q (signal_22170) ) ;
    buf_clk cell_17288 ( .C (clk), .D (signal_22175), .Q (signal_22176) ) ;
    buf_clk cell_17294 ( .C (clk), .D (signal_22181), .Q (signal_22182) ) ;
    buf_clk cell_17300 ( .C (clk), .D (signal_22187), .Q (signal_22188) ) ;
    buf_clk cell_17306 ( .C (clk), .D (signal_22193), .Q (signal_22194) ) ;
    buf_clk cell_17312 ( .C (clk), .D (signal_22199), .Q (signal_22200) ) ;
    buf_clk cell_17318 ( .C (clk), .D (signal_22205), .Q (signal_22206) ) ;
    buf_clk cell_17324 ( .C (clk), .D (signal_22211), .Q (signal_22212) ) ;
    buf_clk cell_17330 ( .C (clk), .D (signal_22217), .Q (signal_22218) ) ;
    buf_clk cell_17336 ( .C (clk), .D (signal_22223), .Q (signal_22224) ) ;
    buf_clk cell_17342 ( .C (clk), .D (signal_22229), .Q (signal_22230) ) ;
    buf_clk cell_17348 ( .C (clk), .D (signal_22235), .Q (signal_22236) ) ;
    buf_clk cell_17354 ( .C (clk), .D (signal_22241), .Q (signal_22242) ) ;
    buf_clk cell_17360 ( .C (clk), .D (signal_22247), .Q (signal_22248) ) ;
    buf_clk cell_17366 ( .C (clk), .D (signal_22253), .Q (signal_22254) ) ;
    buf_clk cell_17372 ( .C (clk), .D (signal_22259), .Q (signal_22260) ) ;
    buf_clk cell_17378 ( .C (clk), .D (signal_22265), .Q (signal_22266) ) ;
    buf_clk cell_17384 ( .C (clk), .D (signal_22271), .Q (signal_22272) ) ;
    buf_clk cell_17390 ( .C (clk), .D (signal_22277), .Q (signal_22278) ) ;
    buf_clk cell_17396 ( .C (clk), .D (signal_22283), .Q (signal_22284) ) ;
    buf_clk cell_17402 ( .C (clk), .D (signal_22289), .Q (signal_22290) ) ;
    buf_clk cell_17408 ( .C (clk), .D (signal_22295), .Q (signal_22296) ) ;
    buf_clk cell_17414 ( .C (clk), .D (signal_22301), .Q (signal_22302) ) ;
    buf_clk cell_17420 ( .C (clk), .D (signal_22307), .Q (signal_22308) ) ;
    buf_clk cell_17426 ( .C (clk), .D (signal_22313), .Q (signal_22314) ) ;
    buf_clk cell_17432 ( .C (clk), .D (signal_22319), .Q (signal_22320) ) ;
    buf_clk cell_17438 ( .C (clk), .D (signal_22325), .Q (signal_22326) ) ;
    buf_clk cell_17444 ( .C (clk), .D (signal_22331), .Q (signal_22332) ) ;
    buf_clk cell_17450 ( .C (clk), .D (signal_22337), .Q (signal_22338) ) ;
    buf_clk cell_17456 ( .C (clk), .D (signal_22343), .Q (signal_22344) ) ;
    buf_clk cell_17462 ( .C (clk), .D (signal_22349), .Q (signal_22350) ) ;
    buf_clk cell_17468 ( .C (clk), .D (signal_22355), .Q (signal_22356) ) ;
    buf_clk cell_17474 ( .C (clk), .D (signal_22361), .Q (signal_22362) ) ;
    buf_clk cell_17480 ( .C (clk), .D (signal_22367), .Q (signal_22368) ) ;
    buf_clk cell_17486 ( .C (clk), .D (signal_22373), .Q (signal_22374) ) ;
    buf_clk cell_17492 ( .C (clk), .D (signal_22379), .Q (signal_22380) ) ;
    buf_clk cell_17498 ( .C (clk), .D (signal_22385), .Q (signal_22386) ) ;
    buf_clk cell_17504 ( .C (clk), .D (signal_22391), .Q (signal_22392) ) ;
    buf_clk cell_17510 ( .C (clk), .D (signal_22397), .Q (signal_22398) ) ;
    buf_clk cell_17516 ( .C (clk), .D (signal_22403), .Q (signal_22404) ) ;
    buf_clk cell_17522 ( .C (clk), .D (signal_22409), .Q (signal_22410) ) ;
    buf_clk cell_17528 ( .C (clk), .D (signal_22415), .Q (signal_22416) ) ;
    buf_clk cell_17534 ( .C (clk), .D (signal_22421), .Q (signal_22422) ) ;
    buf_clk cell_17540 ( .C (clk), .D (signal_22427), .Q (signal_22428) ) ;
    buf_clk cell_17546 ( .C (clk), .D (signal_22433), .Q (signal_22434) ) ;
    buf_clk cell_17552 ( .C (clk), .D (signal_22439), .Q (signal_22440) ) ;
    buf_clk cell_17558 ( .C (clk), .D (signal_22445), .Q (signal_22446) ) ;
    buf_clk cell_17564 ( .C (clk), .D (signal_22451), .Q (signal_22452) ) ;
    buf_clk cell_17570 ( .C (clk), .D (signal_22457), .Q (signal_22458) ) ;
    buf_clk cell_17576 ( .C (clk), .D (signal_22463), .Q (signal_22464) ) ;
    buf_clk cell_17582 ( .C (clk), .D (signal_22469), .Q (signal_22470) ) ;
    buf_clk cell_17588 ( .C (clk), .D (signal_22475), .Q (signal_22476) ) ;
    buf_clk cell_17596 ( .C (clk), .D (signal_22483), .Q (signal_22484) ) ;
    buf_clk cell_17604 ( .C (clk), .D (signal_22491), .Q (signal_22492) ) ;
    buf_clk cell_17612 ( .C (clk), .D (signal_22499), .Q (signal_22500) ) ;
    buf_clk cell_17620 ( .C (clk), .D (signal_22507), .Q (signal_22508) ) ;
    buf_clk cell_17628 ( .C (clk), .D (signal_22515), .Q (signal_22516) ) ;
    buf_clk cell_17636 ( .C (clk), .D (signal_22523), .Q (signal_22524) ) ;
    buf_clk cell_17644 ( .C (clk), .D (signal_22531), .Q (signal_22532) ) ;
    buf_clk cell_17652 ( .C (clk), .D (signal_22539), .Q (signal_22540) ) ;
    buf_clk cell_17660 ( .C (clk), .D (signal_22547), .Q (signal_22548) ) ;
    buf_clk cell_17668 ( .C (clk), .D (signal_22555), .Q (signal_22556) ) ;
    buf_clk cell_17676 ( .C (clk), .D (signal_22563), .Q (signal_22564) ) ;
    buf_clk cell_17684 ( .C (clk), .D (signal_22571), .Q (signal_22572) ) ;
    buf_clk cell_17692 ( .C (clk), .D (signal_22579), .Q (signal_22580) ) ;
    buf_clk cell_17700 ( .C (clk), .D (signal_22587), .Q (signal_22588) ) ;
    buf_clk cell_17708 ( .C (clk), .D (signal_22595), .Q (signal_22596) ) ;
    buf_clk cell_17716 ( .C (clk), .D (signal_22603), .Q (signal_22604) ) ;
    buf_clk cell_17724 ( .C (clk), .D (signal_22611), .Q (signal_22612) ) ;
    buf_clk cell_17732 ( .C (clk), .D (signal_22619), .Q (signal_22620) ) ;
    buf_clk cell_17740 ( .C (clk), .D (signal_22627), .Q (signal_22628) ) ;
    buf_clk cell_17748 ( .C (clk), .D (signal_22635), .Q (signal_22636) ) ;
    buf_clk cell_17756 ( .C (clk), .D (signal_22643), .Q (signal_22644) ) ;
    buf_clk cell_17764 ( .C (clk), .D (signal_22651), .Q (signal_22652) ) ;
    buf_clk cell_17772 ( .C (clk), .D (signal_22659), .Q (signal_22660) ) ;
    buf_clk cell_17780 ( .C (clk), .D (signal_22667), .Q (signal_22668) ) ;
    buf_clk cell_17788 ( .C (clk), .D (signal_22675), .Q (signal_22676) ) ;
    buf_clk cell_17796 ( .C (clk), .D (signal_22683), .Q (signal_22684) ) ;
    buf_clk cell_17804 ( .C (clk), .D (signal_22691), .Q (signal_22692) ) ;
    buf_clk cell_17812 ( .C (clk), .D (signal_22699), .Q (signal_22700) ) ;
    buf_clk cell_17820 ( .C (clk), .D (signal_22707), .Q (signal_22708) ) ;
    buf_clk cell_17828 ( .C (clk), .D (signal_22715), .Q (signal_22716) ) ;
    buf_clk cell_17836 ( .C (clk), .D (signal_22723), .Q (signal_22724) ) ;
    buf_clk cell_17844 ( .C (clk), .D (signal_22731), .Q (signal_22732) ) ;
    buf_clk cell_17852 ( .C (clk), .D (signal_22739), .Q (signal_22740) ) ;
    buf_clk cell_17860 ( .C (clk), .D (signal_22747), .Q (signal_22748) ) ;
    buf_clk cell_17868 ( .C (clk), .D (signal_22755), .Q (signal_22756) ) ;
    buf_clk cell_17876 ( .C (clk), .D (signal_22763), .Q (signal_22764) ) ;
    buf_clk cell_17884 ( .C (clk), .D (signal_22771), .Q (signal_22772) ) ;
    buf_clk cell_17892 ( .C (clk), .D (signal_22779), .Q (signal_22780) ) ;
    buf_clk cell_17900 ( .C (clk), .D (signal_22787), .Q (signal_22788) ) ;
    buf_clk cell_17908 ( .C (clk), .D (signal_22795), .Q (signal_22796) ) ;
    buf_clk cell_17916 ( .C (clk), .D (signal_22803), .Q (signal_22804) ) ;
    buf_clk cell_17924 ( .C (clk), .D (signal_22811), .Q (signal_22812) ) ;
    buf_clk cell_17932 ( .C (clk), .D (signal_22819), .Q (signal_22820) ) ;
    buf_clk cell_17940 ( .C (clk), .D (signal_22827), .Q (signal_22828) ) ;
    buf_clk cell_17948 ( .C (clk), .D (signal_22835), .Q (signal_22836) ) ;
    buf_clk cell_17956 ( .C (clk), .D (signal_22843), .Q (signal_22844) ) ;
    buf_clk cell_17964 ( .C (clk), .D (signal_22851), .Q (signal_22852) ) ;
    buf_clk cell_17972 ( .C (clk), .D (signal_22859), .Q (signal_22860) ) ;
    buf_clk cell_17980 ( .C (clk), .D (signal_22867), .Q (signal_22868) ) ;
    buf_clk cell_17988 ( .C (clk), .D (signal_22875), .Q (signal_22876) ) ;
    buf_clk cell_17996 ( .C (clk), .D (signal_22883), .Q (signal_22884) ) ;
    buf_clk cell_18004 ( .C (clk), .D (signal_22891), .Q (signal_22892) ) ;
    buf_clk cell_18012 ( .C (clk), .D (signal_22899), .Q (signal_22900) ) ;
    buf_clk cell_18020 ( .C (clk), .D (signal_22907), .Q (signal_22908) ) ;
    buf_clk cell_18028 ( .C (clk), .D (signal_22915), .Q (signal_22916) ) ;
    buf_clk cell_18036 ( .C (clk), .D (signal_22923), .Q (signal_22924) ) ;
    buf_clk cell_18044 ( .C (clk), .D (signal_22931), .Q (signal_22932) ) ;
    buf_clk cell_18052 ( .C (clk), .D (signal_22939), .Q (signal_22940) ) ;
    buf_clk cell_18060 ( .C (clk), .D (signal_22947), .Q (signal_22948) ) ;
    buf_clk cell_18068 ( .C (clk), .D (signal_22955), .Q (signal_22956) ) ;
    buf_clk cell_18076 ( .C (clk), .D (signal_22963), .Q (signal_22964) ) ;
    buf_clk cell_18084 ( .C (clk), .D (signal_22971), .Q (signal_22972) ) ;
    buf_clk cell_18092 ( .C (clk), .D (signal_22979), .Q (signal_22980) ) ;
    buf_clk cell_18100 ( .C (clk), .D (signal_22987), .Q (signal_22988) ) ;
    buf_clk cell_18108 ( .C (clk), .D (signal_22995), .Q (signal_22996) ) ;
    buf_clk cell_18116 ( .C (clk), .D (signal_23003), .Q (signal_23004) ) ;
    buf_clk cell_18124 ( .C (clk), .D (signal_23011), .Q (signal_23012) ) ;
    buf_clk cell_18132 ( .C (clk), .D (signal_23019), .Q (signal_23020) ) ;
    buf_clk cell_18140 ( .C (clk), .D (signal_23027), .Q (signal_23028) ) ;
    buf_clk cell_18148 ( .C (clk), .D (signal_23035), .Q (signal_23036) ) ;
    buf_clk cell_18156 ( .C (clk), .D (signal_23043), .Q (signal_23044) ) ;
    buf_clk cell_18164 ( .C (clk), .D (signal_23051), .Q (signal_23052) ) ;
    buf_clk cell_18172 ( .C (clk), .D (signal_23059), .Q (signal_23060) ) ;
    buf_clk cell_18180 ( .C (clk), .D (signal_23067), .Q (signal_23068) ) ;
    buf_clk cell_18188 ( .C (clk), .D (signal_23075), .Q (signal_23076) ) ;
    buf_clk cell_18196 ( .C (clk), .D (signal_23083), .Q (signal_23084) ) ;
    buf_clk cell_18204 ( .C (clk), .D (signal_23091), .Q (signal_23092) ) ;
    buf_clk cell_18212 ( .C (clk), .D (signal_23099), .Q (signal_23100) ) ;
    buf_clk cell_18220 ( .C (clk), .D (signal_23107), .Q (signal_23108) ) ;
    buf_clk cell_18228 ( .C (clk), .D (signal_23115), .Q (signal_23116) ) ;
    buf_clk cell_18236 ( .C (clk), .D (signal_23123), .Q (signal_23124) ) ;
    buf_clk cell_18244 ( .C (clk), .D (signal_23131), .Q (signal_23132) ) ;
    buf_clk cell_18252 ( .C (clk), .D (signal_23139), .Q (signal_23140) ) ;
    buf_clk cell_18260 ( .C (clk), .D (signal_23147), .Q (signal_23148) ) ;
    buf_clk cell_18268 ( .C (clk), .D (signal_23155), .Q (signal_23156) ) ;
    buf_clk cell_18276 ( .C (clk), .D (signal_23163), .Q (signal_23164) ) ;
    buf_clk cell_18284 ( .C (clk), .D (signal_23171), .Q (signal_23172) ) ;
    buf_clk cell_18292 ( .C (clk), .D (signal_23179), .Q (signal_23180) ) ;
    buf_clk cell_18300 ( .C (clk), .D (signal_23187), .Q (signal_23188) ) ;
    buf_clk cell_18308 ( .C (clk), .D (signal_23195), .Q (signal_23196) ) ;
    buf_clk cell_18316 ( .C (clk), .D (signal_23203), .Q (signal_23204) ) ;
    buf_clk cell_18324 ( .C (clk), .D (signal_23211), .Q (signal_23212) ) ;
    buf_clk cell_18332 ( .C (clk), .D (signal_23219), .Q (signal_23220) ) ;
    buf_clk cell_18340 ( .C (clk), .D (signal_23227), .Q (signal_23228) ) ;
    buf_clk cell_18348 ( .C (clk), .D (signal_23235), .Q (signal_23236) ) ;
    buf_clk cell_18356 ( .C (clk), .D (signal_23243), .Q (signal_23244) ) ;
    buf_clk cell_18364 ( .C (clk), .D (signal_23251), .Q (signal_23252) ) ;
    buf_clk cell_18372 ( .C (clk), .D (signal_23259), .Q (signal_23260) ) ;
    buf_clk cell_18380 ( .C (clk), .D (signal_23267), .Q (signal_23268) ) ;
    buf_clk cell_18388 ( .C (clk), .D (signal_23275), .Q (signal_23276) ) ;
    buf_clk cell_18396 ( .C (clk), .D (signal_23283), .Q (signal_23284) ) ;
    buf_clk cell_18408 ( .C (clk), .D (signal_23295), .Q (signal_23296) ) ;
    buf_clk cell_18416 ( .C (clk), .D (signal_23303), .Q (signal_23304) ) ;
    buf_clk cell_18424 ( .C (clk), .D (signal_23311), .Q (signal_23312) ) ;
    buf_clk cell_18432 ( .C (clk), .D (signal_23319), .Q (signal_23320) ) ;
    buf_clk cell_18440 ( .C (clk), .D (signal_23327), .Q (signal_23328) ) ;
    buf_clk cell_18448 ( .C (clk), .D (signal_23335), .Q (signal_23336) ) ;
    buf_clk cell_18456 ( .C (clk), .D (signal_23343), .Q (signal_23344) ) ;
    buf_clk cell_18464 ( .C (clk), .D (signal_23351), .Q (signal_23352) ) ;
    buf_clk cell_18472 ( .C (clk), .D (signal_23359), .Q (signal_23360) ) ;
    buf_clk cell_18480 ( .C (clk), .D (signal_23367), .Q (signal_23368) ) ;
    buf_clk cell_18488 ( .C (clk), .D (signal_23375), .Q (signal_23376) ) ;
    buf_clk cell_18496 ( .C (clk), .D (signal_23383), .Q (signal_23384) ) ;
    buf_clk cell_18504 ( .C (clk), .D (signal_23391), .Q (signal_23392) ) ;
    buf_clk cell_18512 ( .C (clk), .D (signal_23399), .Q (signal_23400) ) ;
    buf_clk cell_18520 ( .C (clk), .D (signal_23407), .Q (signal_23408) ) ;
    buf_clk cell_18528 ( .C (clk), .D (signal_23415), .Q (signal_23416) ) ;
    buf_clk cell_18536 ( .C (clk), .D (signal_23423), .Q (signal_23424) ) ;
    buf_clk cell_18544 ( .C (clk), .D (signal_23431), .Q (signal_23432) ) ;
    buf_clk cell_18552 ( .C (clk), .D (signal_23439), .Q (signal_23440) ) ;
    buf_clk cell_18560 ( .C (clk), .D (signal_23447), .Q (signal_23448) ) ;
    buf_clk cell_18568 ( .C (clk), .D (signal_23455), .Q (signal_23456) ) ;
    buf_clk cell_18576 ( .C (clk), .D (signal_23463), .Q (signal_23464) ) ;
    buf_clk cell_18584 ( .C (clk), .D (signal_23471), .Q (signal_23472) ) ;
    buf_clk cell_18592 ( .C (clk), .D (signal_23479), .Q (signal_23480) ) ;
    buf_clk cell_18600 ( .C (clk), .D (signal_23487), .Q (signal_23488) ) ;
    buf_clk cell_18608 ( .C (clk), .D (signal_23495), .Q (signal_23496) ) ;
    buf_clk cell_18616 ( .C (clk), .D (signal_23503), .Q (signal_23504) ) ;
    buf_clk cell_18624 ( .C (clk), .D (signal_23511), .Q (signal_23512) ) ;
    buf_clk cell_18632 ( .C (clk), .D (signal_23519), .Q (signal_23520) ) ;
    buf_clk cell_18640 ( .C (clk), .D (signal_23527), .Q (signal_23528) ) ;
    buf_clk cell_18652 ( .C (clk), .D (signal_23539), .Q (signal_23540) ) ;
    buf_clk cell_18660 ( .C (clk), .D (signal_23547), .Q (signal_23548) ) ;
    buf_clk cell_18668 ( .C (clk), .D (signal_23555), .Q (signal_23556) ) ;
    buf_clk cell_18676 ( .C (clk), .D (signal_23563), .Q (signal_23564) ) ;
    buf_clk cell_18684 ( .C (clk), .D (signal_23571), .Q (signal_23572) ) ;
    buf_clk cell_18692 ( .C (clk), .D (signal_23579), .Q (signal_23580) ) ;
    buf_clk cell_18700 ( .C (clk), .D (signal_23587), .Q (signal_23588) ) ;
    buf_clk cell_18708 ( .C (clk), .D (signal_23595), .Q (signal_23596) ) ;
    buf_clk cell_18716 ( .C (clk), .D (signal_23603), .Q (signal_23604) ) ;
    buf_clk cell_18724 ( .C (clk), .D (signal_23611), .Q (signal_23612) ) ;
    buf_clk cell_18732 ( .C (clk), .D (signal_23619), .Q (signal_23620) ) ;
    buf_clk cell_18740 ( .C (clk), .D (signal_23627), .Q (signal_23628) ) ;
    buf_clk cell_18752 ( .C (clk), .D (signal_23639), .Q (signal_23640) ) ;
    buf_clk cell_18760 ( .C (clk), .D (signal_23647), .Q (signal_23648) ) ;
    buf_clk cell_18768 ( .C (clk), .D (signal_23655), .Q (signal_23656) ) ;
    buf_clk cell_18776 ( .C (clk), .D (signal_23663), .Q (signal_23664) ) ;
    buf_clk cell_18784 ( .C (clk), .D (signal_23671), .Q (signal_23672) ) ;
    buf_clk cell_18792 ( .C (clk), .D (signal_23679), .Q (signal_23680) ) ;
    buf_clk cell_18800 ( .C (clk), .D (signal_23687), .Q (signal_23688) ) ;
    buf_clk cell_18808 ( .C (clk), .D (signal_23695), .Q (signal_23696) ) ;
    buf_clk cell_18816 ( .C (clk), .D (signal_23703), .Q (signal_23704) ) ;
    buf_clk cell_18824 ( .C (clk), .D (signal_23711), .Q (signal_23712) ) ;
    buf_clk cell_18832 ( .C (clk), .D (signal_23719), .Q (signal_23720) ) ;
    buf_clk cell_18840 ( .C (clk), .D (signal_23727), .Q (signal_23728) ) ;
    buf_clk cell_18848 ( .C (clk), .D (signal_23735), .Q (signal_23736) ) ;
    buf_clk cell_18856 ( .C (clk), .D (signal_23743), .Q (signal_23744) ) ;
    buf_clk cell_18864 ( .C (clk), .D (signal_23751), .Q (signal_23752) ) ;
    buf_clk cell_18872 ( .C (clk), .D (signal_23759), .Q (signal_23760) ) ;
    buf_clk cell_18880 ( .C (clk), .D (signal_23767), .Q (signal_23768) ) ;
    buf_clk cell_18888 ( .C (clk), .D (signal_23775), .Q (signal_23776) ) ;
    buf_clk cell_18896 ( .C (clk), .D (signal_23783), .Q (signal_23784) ) ;
    buf_clk cell_18904 ( .C (clk), .D (signal_23791), .Q (signal_23792) ) ;
    buf_clk cell_18912 ( .C (clk), .D (signal_23799), .Q (signal_23800) ) ;
    buf_clk cell_18920 ( .C (clk), .D (signal_23807), .Q (signal_23808) ) ;
    buf_clk cell_18928 ( .C (clk), .D (signal_23815), .Q (signal_23816) ) ;
    buf_clk cell_18936 ( .C (clk), .D (signal_23823), .Q (signal_23824) ) ;
    buf_clk cell_18944 ( .C (clk), .D (signal_23831), .Q (signal_23832) ) ;
    buf_clk cell_18952 ( .C (clk), .D (signal_23839), .Q (signal_23840) ) ;
    buf_clk cell_18960 ( .C (clk), .D (signal_23847), .Q (signal_23848) ) ;
    buf_clk cell_18968 ( .C (clk), .D (signal_23855), .Q (signal_23856) ) ;
    buf_clk cell_18976 ( .C (clk), .D (signal_23863), .Q (signal_23864) ) ;
    buf_clk cell_18984 ( .C (clk), .D (signal_23871), .Q (signal_23872) ) ;
    buf_clk cell_18992 ( .C (clk), .D (signal_23879), .Q (signal_23880) ) ;
    buf_clk cell_19000 ( .C (clk), .D (signal_23887), .Q (signal_23888) ) ;
    buf_clk cell_19008 ( .C (clk), .D (signal_23895), .Q (signal_23896) ) ;
    buf_clk cell_19016 ( .C (clk), .D (signal_23903), .Q (signal_23904) ) ;
    buf_clk cell_19024 ( .C (clk), .D (signal_23911), .Q (signal_23912) ) ;
    buf_clk cell_19032 ( .C (clk), .D (signal_23919), .Q (signal_23920) ) ;
    buf_clk cell_19040 ( .C (clk), .D (signal_23927), .Q (signal_23928) ) ;
    buf_clk cell_19048 ( .C (clk), .D (signal_23935), .Q (signal_23936) ) ;
    buf_clk cell_19056 ( .C (clk), .D (signal_23943), .Q (signal_23944) ) ;
    buf_clk cell_19064 ( .C (clk), .D (signal_23951), .Q (signal_23952) ) ;
    buf_clk cell_19072 ( .C (clk), .D (signal_23959), .Q (signal_23960) ) ;
    buf_clk cell_19080 ( .C (clk), .D (signal_23967), .Q (signal_23968) ) ;
    buf_clk cell_19088 ( .C (clk), .D (signal_23975), .Q (signal_23976) ) ;
    buf_clk cell_19096 ( .C (clk), .D (signal_23983), .Q (signal_23984) ) ;
    buf_clk cell_19104 ( .C (clk), .D (signal_23991), .Q (signal_23992) ) ;
    buf_clk cell_19112 ( .C (clk), .D (signal_23999), .Q (signal_24000) ) ;

    /* cells in depth 5 */
    buf_clk cell_8221 ( .C (clk), .D (signal_12790), .Q (signal_13109) ) ;
    buf_clk cell_8223 ( .C (clk), .D (signal_12792), .Q (signal_13111) ) ;
    buf_clk cell_8225 ( .C (clk), .D (signal_5607), .Q (signal_13113) ) ;
    buf_clk cell_8227 ( .C (clk), .D (signal_8927), .Q (signal_13115) ) ;
    buf_clk cell_8229 ( .C (clk), .D (signal_12794), .Q (signal_13117) ) ;
    buf_clk cell_8231 ( .C (clk), .D (signal_12796), .Q (signal_13119) ) ;
    buf_clk cell_8233 ( .C (clk), .D (signal_5713), .Q (signal_13121) ) ;
    buf_clk cell_8235 ( .C (clk), .D (signal_9033), .Q (signal_13123) ) ;
    buf_clk cell_8237 ( .C (clk), .D (signal_12802), .Q (signal_13125) ) ;
    buf_clk cell_8239 ( .C (clk), .D (signal_12804), .Q (signal_13127) ) ;
    buf_clk cell_8241 ( .C (clk), .D (signal_5617), .Q (signal_13129) ) ;
    buf_clk cell_8243 ( .C (clk), .D (signal_8931), .Q (signal_13131) ) ;
    buf_clk cell_8245 ( .C (clk), .D (signal_12806), .Q (signal_13133) ) ;
    buf_clk cell_8247 ( .C (clk), .D (signal_12808), .Q (signal_13135) ) ;
    buf_clk cell_8249 ( .C (clk), .D (signal_5726), .Q (signal_13137) ) ;
    buf_clk cell_8251 ( .C (clk), .D (signal_9034), .Q (signal_13139) ) ;
    buf_clk cell_8253 ( .C (clk), .D (signal_12814), .Q (signal_13141) ) ;
    buf_clk cell_8255 ( .C (clk), .D (signal_12816), .Q (signal_13143) ) ;
    buf_clk cell_8257 ( .C (clk), .D (signal_5627), .Q (signal_13145) ) ;
    buf_clk cell_8259 ( .C (clk), .D (signal_8935), .Q (signal_13147) ) ;
    buf_clk cell_8261 ( .C (clk), .D (signal_12818), .Q (signal_13149) ) ;
    buf_clk cell_8263 ( .C (clk), .D (signal_12820), .Q (signal_13151) ) ;
    buf_clk cell_8265 ( .C (clk), .D (signal_5739), .Q (signal_13153) ) ;
    buf_clk cell_8267 ( .C (clk), .D (signal_9035), .Q (signal_13155) ) ;
    buf_clk cell_8269 ( .C (clk), .D (signal_12826), .Q (signal_13157) ) ;
    buf_clk cell_8271 ( .C (clk), .D (signal_12828), .Q (signal_13159) ) ;
    buf_clk cell_8273 ( .C (clk), .D (signal_5631), .Q (signal_13161) ) ;
    buf_clk cell_8275 ( .C (clk), .D (signal_8908), .Q (signal_13163) ) ;
    buf_clk cell_8277 ( .C (clk), .D (signal_12830), .Q (signal_13165) ) ;
    buf_clk cell_8279 ( .C (clk), .D (signal_12832), .Q (signal_13167) ) ;
    buf_clk cell_8281 ( .C (clk), .D (signal_5740), .Q (signal_13169) ) ;
    buf_clk cell_8283 ( .C (clk), .D (signal_9017), .Q (signal_13171) ) ;
    buf_clk cell_8285 ( .C (clk), .D (signal_12838), .Q (signal_13173) ) ;
    buf_clk cell_8287 ( .C (clk), .D (signal_12840), .Q (signal_13175) ) ;
    buf_clk cell_8289 ( .C (clk), .D (signal_5635), .Q (signal_13177) ) ;
    buf_clk cell_8291 ( .C (clk), .D (signal_8912), .Q (signal_13179) ) ;
    buf_clk cell_8293 ( .C (clk), .D (signal_12842), .Q (signal_13181) ) ;
    buf_clk cell_8295 ( .C (clk), .D (signal_12844), .Q (signal_13183) ) ;
    buf_clk cell_8297 ( .C (clk), .D (signal_5741), .Q (signal_13185) ) ;
    buf_clk cell_8299 ( .C (clk), .D (signal_9018), .Q (signal_13187) ) ;
    buf_clk cell_8301 ( .C (clk), .D (signal_12850), .Q (signal_13189) ) ;
    buf_clk cell_8303 ( .C (clk), .D (signal_12852), .Q (signal_13191) ) ;
    buf_clk cell_8305 ( .C (clk), .D (signal_5639), .Q (signal_13193) ) ;
    buf_clk cell_8307 ( .C (clk), .D (signal_8916), .Q (signal_13195) ) ;
    buf_clk cell_8309 ( .C (clk), .D (signal_12854), .Q (signal_13197) ) ;
    buf_clk cell_8311 ( .C (clk), .D (signal_12856), .Q (signal_13199) ) ;
    buf_clk cell_8313 ( .C (clk), .D (signal_5742), .Q (signal_13201) ) ;
    buf_clk cell_8315 ( .C (clk), .D (signal_9019), .Q (signal_13203) ) ;
    buf_clk cell_8317 ( .C (clk), .D (signal_12862), .Q (signal_13205) ) ;
    buf_clk cell_8319 ( .C (clk), .D (signal_12864), .Q (signal_13207) ) ;
    buf_clk cell_8321 ( .C (clk), .D (signal_5643), .Q (signal_13209) ) ;
    buf_clk cell_8323 ( .C (clk), .D (signal_8920), .Q (signal_13211) ) ;
    buf_clk cell_8325 ( .C (clk), .D (signal_12866), .Q (signal_13213) ) ;
    buf_clk cell_8327 ( .C (clk), .D (signal_12868), .Q (signal_13215) ) ;
    buf_clk cell_8329 ( .C (clk), .D (signal_5743), .Q (signal_13217) ) ;
    buf_clk cell_8331 ( .C (clk), .D (signal_9020), .Q (signal_13219) ) ;
    buf_clk cell_8333 ( .C (clk), .D (signal_12874), .Q (signal_13221) ) ;
    buf_clk cell_8335 ( .C (clk), .D (signal_12876), .Q (signal_13223) ) ;
    buf_clk cell_8337 ( .C (clk), .D (signal_5688), .Q (signal_13225) ) ;
    buf_clk cell_8339 ( .C (clk), .D (signal_8968), .Q (signal_13227) ) ;
    buf_clk cell_8341 ( .C (clk), .D (signal_12878), .Q (signal_13229) ) ;
    buf_clk cell_8343 ( .C (clk), .D (signal_12880), .Q (signal_13231) ) ;
    buf_clk cell_8345 ( .C (clk), .D (signal_5796), .Q (signal_13233) ) ;
    buf_clk cell_8347 ( .C (clk), .D (signal_9088), .Q (signal_13235) ) ;
    buf_clk cell_8349 ( .C (clk), .D (signal_12886), .Q (signal_13237) ) ;
    buf_clk cell_8351 ( .C (clk), .D (signal_12888), .Q (signal_13239) ) ;
    buf_clk cell_8353 ( .C (clk), .D (signal_5692), .Q (signal_13241) ) ;
    buf_clk cell_8355 ( .C (clk), .D (signal_8972), .Q (signal_13243) ) ;
    buf_clk cell_8357 ( .C (clk), .D (signal_12890), .Q (signal_13245) ) ;
    buf_clk cell_8359 ( .C (clk), .D (signal_12892), .Q (signal_13247) ) ;
    buf_clk cell_8361 ( .C (clk), .D (signal_5797), .Q (signal_13249) ) ;
    buf_clk cell_8363 ( .C (clk), .D (signal_9089), .Q (signal_13251) ) ;
    buf_clk cell_8365 ( .C (clk), .D (signal_12898), .Q (signal_13253) ) ;
    buf_clk cell_8367 ( .C (clk), .D (signal_12900), .Q (signal_13255) ) ;
    buf_clk cell_8369 ( .C (clk), .D (signal_5696), .Q (signal_13257) ) ;
    buf_clk cell_8371 ( .C (clk), .D (signal_8976), .Q (signal_13259) ) ;
    buf_clk cell_8373 ( .C (clk), .D (signal_12902), .Q (signal_13261) ) ;
    buf_clk cell_8375 ( .C (clk), .D (signal_12904), .Q (signal_13263) ) ;
    buf_clk cell_8377 ( .C (clk), .D (signal_5798), .Q (signal_13265) ) ;
    buf_clk cell_8379 ( .C (clk), .D (signal_9090), .Q (signal_13267) ) ;
    buf_clk cell_8381 ( .C (clk), .D (signal_12910), .Q (signal_13269) ) ;
    buf_clk cell_8383 ( .C (clk), .D (signal_12912), .Q (signal_13271) ) ;
    buf_clk cell_8385 ( .C (clk), .D (signal_5700), .Q (signal_13273) ) ;
    buf_clk cell_8387 ( .C (clk), .D (signal_8980), .Q (signal_13275) ) ;
    buf_clk cell_8389 ( .C (clk), .D (signal_12914), .Q (signal_13277) ) ;
    buf_clk cell_8391 ( .C (clk), .D (signal_12916), .Q (signal_13279) ) ;
    buf_clk cell_8393 ( .C (clk), .D (signal_5799), .Q (signal_13281) ) ;
    buf_clk cell_8395 ( .C (clk), .D (signal_9091), .Q (signal_13283) ) ;
    buf_clk cell_8397 ( .C (clk), .D (signal_12922), .Q (signal_13285) ) ;
    buf_clk cell_8399 ( .C (clk), .D (signal_12924), .Q (signal_13287) ) ;
    buf_clk cell_8401 ( .C (clk), .D (signal_5704), .Q (signal_13289) ) ;
    buf_clk cell_8403 ( .C (clk), .D (signal_8984), .Q (signal_13291) ) ;
    buf_clk cell_8405 ( .C (clk), .D (signal_12926), .Q (signal_13293) ) ;
    buf_clk cell_8407 ( .C (clk), .D (signal_12928), .Q (signal_13295) ) ;
    buf_clk cell_8409 ( .C (clk), .D (signal_5800), .Q (signal_13297) ) ;
    buf_clk cell_8411 ( .C (clk), .D (signal_9092), .Q (signal_13299) ) ;
    buf_clk cell_8413 ( .C (clk), .D (signal_12934), .Q (signal_13301) ) ;
    buf_clk cell_8415 ( .C (clk), .D (signal_12936), .Q (signal_13303) ) ;
    buf_clk cell_8417 ( .C (clk), .D (signal_5708), .Q (signal_13305) ) ;
    buf_clk cell_8419 ( .C (clk), .D (signal_8988), .Q (signal_13307) ) ;
    buf_clk cell_8421 ( .C (clk), .D (signal_12938), .Q (signal_13309) ) ;
    buf_clk cell_8423 ( .C (clk), .D (signal_12940), .Q (signal_13311) ) ;
    buf_clk cell_8425 ( .C (clk), .D (signal_5801), .Q (signal_13313) ) ;
    buf_clk cell_8427 ( .C (clk), .D (signal_9093), .Q (signal_13315) ) ;
    buf_clk cell_8429 ( .C (clk), .D (signal_12946), .Q (signal_13317) ) ;
    buf_clk cell_8431 ( .C (clk), .D (signal_12948), .Q (signal_13319) ) ;
    buf_clk cell_8433 ( .C (clk), .D (signal_5712), .Q (signal_13321) ) ;
    buf_clk cell_8435 ( .C (clk), .D (signal_8992), .Q (signal_13323) ) ;
    buf_clk cell_8437 ( .C (clk), .D (signal_12950), .Q (signal_13325) ) ;
    buf_clk cell_8439 ( .C (clk), .D (signal_12952), .Q (signal_13327) ) ;
    buf_clk cell_8441 ( .C (clk), .D (signal_5802), .Q (signal_13329) ) ;
    buf_clk cell_8443 ( .C (clk), .D (signal_9094), .Q (signal_13331) ) ;
    buf_clk cell_8445 ( .C (clk), .D (signal_12962), .Q (signal_13333) ) ;
    buf_clk cell_8447 ( .C (clk), .D (signal_12964), .Q (signal_13335) ) ;
    buf_clk cell_8449 ( .C (clk), .D (signal_5717), .Q (signal_13337) ) ;
    buf_clk cell_8451 ( .C (clk), .D (signal_8996), .Q (signal_13339) ) ;
    buf_clk cell_8453 ( .C (clk), .D (signal_12966), .Q (signal_13341) ) ;
    buf_clk cell_8455 ( .C (clk), .D (signal_12968), .Q (signal_13343) ) ;
    buf_clk cell_8457 ( .C (clk), .D (signal_5807), .Q (signal_13345) ) ;
    buf_clk cell_8459 ( .C (clk), .D (signal_9095), .Q (signal_13347) ) ;
    buf_clk cell_8461 ( .C (clk), .D (signal_12974), .Q (signal_13349) ) ;
    buf_clk cell_8463 ( .C (clk), .D (signal_12976), .Q (signal_13351) ) ;
    buf_clk cell_8465 ( .C (clk), .D (signal_5721), .Q (signal_13353) ) ;
    buf_clk cell_8467 ( .C (clk), .D (signal_9000), .Q (signal_13355) ) ;
    buf_clk cell_8469 ( .C (clk), .D (signal_12978), .Q (signal_13357) ) ;
    buf_clk cell_8471 ( .C (clk), .D (signal_12980), .Q (signal_13359) ) ;
    buf_clk cell_8473 ( .C (clk), .D (signal_5808), .Q (signal_13361) ) ;
    buf_clk cell_8475 ( .C (clk), .D (signal_9096), .Q (signal_13363) ) ;
    buf_clk cell_8477 ( .C (clk), .D (signal_12986), .Q (signal_13365) ) ;
    buf_clk cell_8479 ( .C (clk), .D (signal_12988), .Q (signal_13367) ) ;
    buf_clk cell_8481 ( .C (clk), .D (signal_5725), .Q (signal_13369) ) ;
    buf_clk cell_8483 ( .C (clk), .D (signal_9004), .Q (signal_13371) ) ;
    buf_clk cell_8485 ( .C (clk), .D (signal_12990), .Q (signal_13373) ) ;
    buf_clk cell_8487 ( .C (clk), .D (signal_12992), .Q (signal_13375) ) ;
    buf_clk cell_8489 ( .C (clk), .D (signal_5809), .Q (signal_13377) ) ;
    buf_clk cell_8491 ( .C (clk), .D (signal_9097), .Q (signal_13379) ) ;
    buf_clk cell_8493 ( .C (clk), .D (signal_13002), .Q (signal_13381) ) ;
    buf_clk cell_8495 ( .C (clk), .D (signal_13004), .Q (signal_13383) ) ;
    buf_clk cell_8497 ( .C (clk), .D (signal_5730), .Q (signal_13385) ) ;
    buf_clk cell_8499 ( .C (clk), .D (signal_9008), .Q (signal_13387) ) ;
    buf_clk cell_8501 ( .C (clk), .D (signal_13006), .Q (signal_13389) ) ;
    buf_clk cell_8503 ( .C (clk), .D (signal_13008), .Q (signal_13391) ) ;
    buf_clk cell_8505 ( .C (clk), .D (signal_5814), .Q (signal_13393) ) ;
    buf_clk cell_8507 ( .C (clk), .D (signal_9098), .Q (signal_13395) ) ;
    buf_clk cell_8509 ( .C (clk), .D (signal_13014), .Q (signal_13397) ) ;
    buf_clk cell_8511 ( .C (clk), .D (signal_13016), .Q (signal_13399) ) ;
    buf_clk cell_8513 ( .C (clk), .D (signal_5734), .Q (signal_13401) ) ;
    buf_clk cell_8515 ( .C (clk), .D (signal_9012), .Q (signal_13403) ) ;
    buf_clk cell_8517 ( .C (clk), .D (signal_13018), .Q (signal_13405) ) ;
    buf_clk cell_8519 ( .C (clk), .D (signal_13020), .Q (signal_13407) ) ;
    buf_clk cell_8521 ( .C (clk), .D (signal_5815), .Q (signal_13409) ) ;
    buf_clk cell_8523 ( .C (clk), .D (signal_9099), .Q (signal_13411) ) ;
    buf_clk cell_8525 ( .C (clk), .D (signal_13026), .Q (signal_13413) ) ;
    buf_clk cell_8527 ( .C (clk), .D (signal_13028), .Q (signal_13415) ) ;
    buf_clk cell_8529 ( .C (clk), .D (signal_5738), .Q (signal_13417) ) ;
    buf_clk cell_8531 ( .C (clk), .D (signal_9016), .Q (signal_13419) ) ;
    buf_clk cell_8533 ( .C (clk), .D (signal_13030), .Q (signal_13421) ) ;
    buf_clk cell_8535 ( .C (clk), .D (signal_13032), .Q (signal_13423) ) ;
    buf_clk cell_8537 ( .C (clk), .D (signal_5816), .Q (signal_13425) ) ;
    buf_clk cell_8539 ( .C (clk), .D (signal_9100), .Q (signal_13427) ) ;
    buf_clk cell_8545 ( .C (clk), .D (signal_13432), .Q (signal_13433) ) ;
    buf_clk cell_8553 ( .C (clk), .D (signal_13440), .Q (signal_13441) ) ;
    buf_clk cell_8561 ( .C (clk), .D (signal_13448), .Q (signal_13449) ) ;
    buf_clk cell_8569 ( .C (clk), .D (signal_13456), .Q (signal_13457) ) ;
    buf_clk cell_8577 ( .C (clk), .D (signal_13464), .Q (signal_13465) ) ;
    buf_clk cell_8585 ( .C (clk), .D (signal_13472), .Q (signal_13473) ) ;
    buf_clk cell_8593 ( .C (clk), .D (signal_13480), .Q (signal_13481) ) ;
    buf_clk cell_8601 ( .C (clk), .D (signal_13488), .Q (signal_13489) ) ;
    buf_clk cell_8609 ( .C (clk), .D (signal_13496), .Q (signal_13497) ) ;
    buf_clk cell_8617 ( .C (clk), .D (signal_13504), .Q (signal_13505) ) ;
    buf_clk cell_8625 ( .C (clk), .D (signal_13512), .Q (signal_13513) ) ;
    buf_clk cell_8633 ( .C (clk), .D (signal_13520), .Q (signal_13521) ) ;
    buf_clk cell_8641 ( .C (clk), .D (signal_13528), .Q (signal_13529) ) ;
    buf_clk cell_8649 ( .C (clk), .D (signal_13536), .Q (signal_13537) ) ;
    buf_clk cell_8657 ( .C (clk), .D (signal_13544), .Q (signal_13545) ) ;
    buf_clk cell_8665 ( .C (clk), .D (signal_13552), .Q (signal_13553) ) ;
    buf_clk cell_8673 ( .C (clk), .D (signal_13560), .Q (signal_13561) ) ;
    buf_clk cell_8681 ( .C (clk), .D (signal_13568), .Q (signal_13569) ) ;
    buf_clk cell_8689 ( .C (clk), .D (signal_13576), .Q (signal_13577) ) ;
    buf_clk cell_8697 ( .C (clk), .D (signal_13584), .Q (signal_13585) ) ;
    buf_clk cell_8705 ( .C (clk), .D (signal_13592), .Q (signal_13593) ) ;
    buf_clk cell_8713 ( .C (clk), .D (signal_13600), .Q (signal_13601) ) ;
    buf_clk cell_8721 ( .C (clk), .D (signal_13608), .Q (signal_13609) ) ;
    buf_clk cell_8729 ( .C (clk), .D (signal_13616), .Q (signal_13617) ) ;
    buf_clk cell_8737 ( .C (clk), .D (signal_13624), .Q (signal_13625) ) ;
    buf_clk cell_8745 ( .C (clk), .D (signal_13632), .Q (signal_13633) ) ;
    buf_clk cell_8753 ( .C (clk), .D (signal_13640), .Q (signal_13641) ) ;
    buf_clk cell_8761 ( .C (clk), .D (signal_13648), .Q (signal_13649) ) ;
    buf_clk cell_8769 ( .C (clk), .D (signal_13656), .Q (signal_13657) ) ;
    buf_clk cell_8777 ( .C (clk), .D (signal_13664), .Q (signal_13665) ) ;
    buf_clk cell_8785 ( .C (clk), .D (signal_13672), .Q (signal_13673) ) ;
    buf_clk cell_8793 ( .C (clk), .D (signal_13680), .Q (signal_13681) ) ;
    buf_clk cell_8801 ( .C (clk), .D (signal_13688), .Q (signal_13689) ) ;
    buf_clk cell_8809 ( .C (clk), .D (signal_13696), .Q (signal_13697) ) ;
    buf_clk cell_8817 ( .C (clk), .D (signal_13704), .Q (signal_13705) ) ;
    buf_clk cell_8825 ( .C (clk), .D (signal_13712), .Q (signal_13713) ) ;
    buf_clk cell_8833 ( .C (clk), .D (signal_13720), .Q (signal_13721) ) ;
    buf_clk cell_8841 ( .C (clk), .D (signal_13728), .Q (signal_13729) ) ;
    buf_clk cell_8849 ( .C (clk), .D (signal_13736), .Q (signal_13737) ) ;
    buf_clk cell_8857 ( .C (clk), .D (signal_13744), .Q (signal_13745) ) ;
    buf_clk cell_8865 ( .C (clk), .D (signal_13752), .Q (signal_13753) ) ;
    buf_clk cell_8873 ( .C (clk), .D (signal_13760), .Q (signal_13761) ) ;
    buf_clk cell_8881 ( .C (clk), .D (signal_13768), .Q (signal_13769) ) ;
    buf_clk cell_8889 ( .C (clk), .D (signal_13776), .Q (signal_13777) ) ;
    buf_clk cell_8897 ( .C (clk), .D (signal_13784), .Q (signal_13785) ) ;
    buf_clk cell_8905 ( .C (clk), .D (signal_13792), .Q (signal_13793) ) ;
    buf_clk cell_8913 ( .C (clk), .D (signal_13800), .Q (signal_13801) ) ;
    buf_clk cell_8921 ( .C (clk), .D (signal_13808), .Q (signal_13809) ) ;
    buf_clk cell_8929 ( .C (clk), .D (signal_13816), .Q (signal_13817) ) ;
    buf_clk cell_8937 ( .C (clk), .D (signal_13824), .Q (signal_13825) ) ;
    buf_clk cell_8945 ( .C (clk), .D (signal_13832), .Q (signal_13833) ) ;
    buf_clk cell_8953 ( .C (clk), .D (signal_13840), .Q (signal_13841) ) ;
    buf_clk cell_8961 ( .C (clk), .D (signal_13848), .Q (signal_13849) ) ;
    buf_clk cell_8969 ( .C (clk), .D (signal_13856), .Q (signal_13857) ) ;
    buf_clk cell_8977 ( .C (clk), .D (signal_13864), .Q (signal_13865) ) ;
    buf_clk cell_8985 ( .C (clk), .D (signal_13872), .Q (signal_13873) ) ;
    buf_clk cell_8993 ( .C (clk), .D (signal_13880), .Q (signal_13881) ) ;
    buf_clk cell_9001 ( .C (clk), .D (signal_13888), .Q (signal_13889) ) ;
    buf_clk cell_9009 ( .C (clk), .D (signal_13896), .Q (signal_13897) ) ;
    buf_clk cell_9017 ( .C (clk), .D (signal_13904), .Q (signal_13905) ) ;
    buf_clk cell_9025 ( .C (clk), .D (signal_13912), .Q (signal_13913) ) ;
    buf_clk cell_9033 ( .C (clk), .D (signal_13920), .Q (signal_13921) ) ;
    buf_clk cell_9041 ( .C (clk), .D (signal_13928), .Q (signal_13929) ) ;
    buf_clk cell_9049 ( .C (clk), .D (signal_13936), .Q (signal_13937) ) ;
    buf_clk cell_9057 ( .C (clk), .D (signal_13944), .Q (signal_13945) ) ;
    buf_clk cell_9065 ( .C (clk), .D (signal_13952), .Q (signal_13953) ) ;
    buf_clk cell_9073 ( .C (clk), .D (signal_13960), .Q (signal_13961) ) ;
    buf_clk cell_9081 ( .C (clk), .D (signal_13968), .Q (signal_13969) ) ;
    buf_clk cell_9089 ( .C (clk), .D (signal_13976), .Q (signal_13977) ) ;
    buf_clk cell_9097 ( .C (clk), .D (signal_13984), .Q (signal_13985) ) ;
    buf_clk cell_9105 ( .C (clk), .D (signal_13992), .Q (signal_13993) ) ;
    buf_clk cell_9113 ( .C (clk), .D (signal_14000), .Q (signal_14001) ) ;
    buf_clk cell_9121 ( .C (clk), .D (signal_14008), .Q (signal_14009) ) ;
    buf_clk cell_9129 ( .C (clk), .D (signal_14016), .Q (signal_14017) ) ;
    buf_clk cell_9137 ( .C (clk), .D (signal_14024), .Q (signal_14025) ) ;
    buf_clk cell_9145 ( .C (clk), .D (signal_14032), .Q (signal_14033) ) ;
    buf_clk cell_9153 ( .C (clk), .D (signal_14040), .Q (signal_14041) ) ;
    buf_clk cell_9161 ( .C (clk), .D (signal_14048), .Q (signal_14049) ) ;
    buf_clk cell_9169 ( .C (clk), .D (signal_14056), .Q (signal_14057) ) ;
    buf_clk cell_9177 ( .C (clk), .D (signal_14064), .Q (signal_14065) ) ;
    buf_clk cell_9185 ( .C (clk), .D (signal_14072), .Q (signal_14073) ) ;
    buf_clk cell_9193 ( .C (clk), .D (signal_14080), .Q (signal_14081) ) ;
    buf_clk cell_9201 ( .C (clk), .D (signal_14088), .Q (signal_14089) ) ;
    buf_clk cell_9209 ( .C (clk), .D (signal_14096), .Q (signal_14097) ) ;
    buf_clk cell_9217 ( .C (clk), .D (signal_14104), .Q (signal_14105) ) ;
    buf_clk cell_9225 ( .C (clk), .D (signal_14112), .Q (signal_14113) ) ;
    buf_clk cell_9233 ( .C (clk), .D (signal_14120), .Q (signal_14121) ) ;
    buf_clk cell_9241 ( .C (clk), .D (signal_14128), .Q (signal_14129) ) ;
    buf_clk cell_9249 ( .C (clk), .D (signal_14136), .Q (signal_14137) ) ;
    buf_clk cell_9257 ( .C (clk), .D (signal_14144), .Q (signal_14145) ) ;
    buf_clk cell_9265 ( .C (clk), .D (signal_14152), .Q (signal_14153) ) ;
    buf_clk cell_9273 ( .C (clk), .D (signal_14160), .Q (signal_14161) ) ;
    buf_clk cell_9281 ( .C (clk), .D (signal_14168), .Q (signal_14169) ) ;
    buf_clk cell_9289 ( .C (clk), .D (signal_14176), .Q (signal_14177) ) ;
    buf_clk cell_9297 ( .C (clk), .D (signal_14184), .Q (signal_14185) ) ;
    buf_clk cell_9305 ( .C (clk), .D (signal_14192), .Q (signal_14193) ) ;
    buf_clk cell_9313 ( .C (clk), .D (signal_14200), .Q (signal_14201) ) ;
    buf_clk cell_9321 ( .C (clk), .D (signal_14208), .Q (signal_14209) ) ;
    buf_clk cell_9329 ( .C (clk), .D (signal_14216), .Q (signal_14217) ) ;
    buf_clk cell_9337 ( .C (clk), .D (signal_14224), .Q (signal_14225) ) ;
    buf_clk cell_9345 ( .C (clk), .D (signal_14232), .Q (signal_14233) ) ;
    buf_clk cell_9353 ( .C (clk), .D (signal_14240), .Q (signal_14241) ) ;
    buf_clk cell_9361 ( .C (clk), .D (signal_14248), .Q (signal_14249) ) ;
    buf_clk cell_9369 ( .C (clk), .D (signal_14256), .Q (signal_14257) ) ;
    buf_clk cell_9377 ( .C (clk), .D (signal_14264), .Q (signal_14265) ) ;
    buf_clk cell_9385 ( .C (clk), .D (signal_14272), .Q (signal_14273) ) ;
    buf_clk cell_9393 ( .C (clk), .D (signal_14280), .Q (signal_14281) ) ;
    buf_clk cell_9401 ( .C (clk), .D (signal_14288), .Q (signal_14289) ) ;
    buf_clk cell_9409 ( .C (clk), .D (signal_14296), .Q (signal_14297) ) ;
    buf_clk cell_9417 ( .C (clk), .D (signal_14304), .Q (signal_14305) ) ;
    buf_clk cell_9425 ( .C (clk), .D (signal_14312), .Q (signal_14313) ) ;
    buf_clk cell_9433 ( .C (clk), .D (signal_14320), .Q (signal_14321) ) ;
    buf_clk cell_9441 ( .C (clk), .D (signal_14328), .Q (signal_14329) ) ;
    buf_clk cell_9449 ( .C (clk), .D (signal_14336), .Q (signal_14337) ) ;
    buf_clk cell_9457 ( .C (clk), .D (signal_14344), .Q (signal_14345) ) ;
    buf_clk cell_9465 ( .C (clk), .D (signal_14352), .Q (signal_14353) ) ;
    buf_clk cell_9473 ( .C (clk), .D (signal_14360), .Q (signal_14361) ) ;
    buf_clk cell_9481 ( .C (clk), .D (signal_14368), .Q (signal_14369) ) ;
    buf_clk cell_9489 ( .C (clk), .D (signal_14376), .Q (signal_14377) ) ;
    buf_clk cell_9497 ( .C (clk), .D (signal_14384), .Q (signal_14385) ) ;
    buf_clk cell_9505 ( .C (clk), .D (signal_14392), .Q (signal_14393) ) ;
    buf_clk cell_9513 ( .C (clk), .D (signal_14400), .Q (signal_14401) ) ;
    buf_clk cell_9521 ( .C (clk), .D (signal_14408), .Q (signal_14409) ) ;
    buf_clk cell_9529 ( .C (clk), .D (signal_14416), .Q (signal_14417) ) ;
    buf_clk cell_9537 ( .C (clk), .D (signal_14424), .Q (signal_14425) ) ;
    buf_clk cell_9545 ( .C (clk), .D (signal_14432), .Q (signal_14433) ) ;
    buf_clk cell_9553 ( .C (clk), .D (signal_14440), .Q (signal_14441) ) ;
    buf_clk cell_9561 ( .C (clk), .D (signal_14448), .Q (signal_14449) ) ;
    buf_clk cell_9569 ( .C (clk), .D (signal_14456), .Q (signal_14457) ) ;
    buf_clk cell_9577 ( .C (clk), .D (signal_14464), .Q (signal_14465) ) ;
    buf_clk cell_9585 ( .C (clk), .D (signal_14472), .Q (signal_14473) ) ;
    buf_clk cell_9593 ( .C (clk), .D (signal_14480), .Q (signal_14481) ) ;
    buf_clk cell_9601 ( .C (clk), .D (signal_14488), .Q (signal_14489) ) ;
    buf_clk cell_9609 ( .C (clk), .D (signal_14496), .Q (signal_14497) ) ;
    buf_clk cell_9617 ( .C (clk), .D (signal_14504), .Q (signal_14505) ) ;
    buf_clk cell_9625 ( .C (clk), .D (signal_14512), .Q (signal_14513) ) ;
    buf_clk cell_9633 ( .C (clk), .D (signal_14520), .Q (signal_14521) ) ;
    buf_clk cell_9641 ( .C (clk), .D (signal_14528), .Q (signal_14529) ) ;
    buf_clk cell_9649 ( .C (clk), .D (signal_14536), .Q (signal_14537) ) ;
    buf_clk cell_9657 ( .C (clk), .D (signal_14544), .Q (signal_14545) ) ;
    buf_clk cell_9665 ( .C (clk), .D (signal_14552), .Q (signal_14553) ) ;
    buf_clk cell_9673 ( .C (clk), .D (signal_14560), .Q (signal_14561) ) ;
    buf_clk cell_9681 ( .C (clk), .D (signal_14568), .Q (signal_14569) ) ;
    buf_clk cell_9689 ( .C (clk), .D (signal_14576), .Q (signal_14577) ) ;
    buf_clk cell_9697 ( .C (clk), .D (signal_14584), .Q (signal_14585) ) ;
    buf_clk cell_9705 ( .C (clk), .D (signal_14592), .Q (signal_14593) ) ;
    buf_clk cell_9713 ( .C (clk), .D (signal_14600), .Q (signal_14601) ) ;
    buf_clk cell_9721 ( .C (clk), .D (signal_14608), .Q (signal_14609) ) ;
    buf_clk cell_9729 ( .C (clk), .D (signal_14616), .Q (signal_14617) ) ;
    buf_clk cell_9737 ( .C (clk), .D (signal_14624), .Q (signal_14625) ) ;
    buf_clk cell_9745 ( .C (clk), .D (signal_14632), .Q (signal_14633) ) ;
    buf_clk cell_9753 ( .C (clk), .D (signal_14640), .Q (signal_14641) ) ;
    buf_clk cell_9761 ( .C (clk), .D (signal_14648), .Q (signal_14649) ) ;
    buf_clk cell_9769 ( .C (clk), .D (signal_14656), .Q (signal_14657) ) ;
    buf_clk cell_9777 ( .C (clk), .D (signal_14664), .Q (signal_14665) ) ;
    buf_clk cell_9785 ( .C (clk), .D (signal_14672), .Q (signal_14673) ) ;
    buf_clk cell_9793 ( .C (clk), .D (signal_14680), .Q (signal_14681) ) ;
    buf_clk cell_9801 ( .C (clk), .D (signal_14688), .Q (signal_14689) ) ;
    buf_clk cell_9809 ( .C (clk), .D (signal_14696), .Q (signal_14697) ) ;
    buf_clk cell_9817 ( .C (clk), .D (signal_14704), .Q (signal_14705) ) ;
    buf_clk cell_9825 ( .C (clk), .D (signal_14712), .Q (signal_14713) ) ;
    buf_clk cell_9833 ( .C (clk), .D (signal_14720), .Q (signal_14721) ) ;
    buf_clk cell_9841 ( .C (clk), .D (signal_14728), .Q (signal_14729) ) ;
    buf_clk cell_9849 ( .C (clk), .D (signal_14736), .Q (signal_14737) ) ;
    buf_clk cell_9857 ( .C (clk), .D (signal_14744), .Q (signal_14745) ) ;
    buf_clk cell_9865 ( .C (clk), .D (signal_14752), .Q (signal_14753) ) ;
    buf_clk cell_9873 ( .C (clk), .D (signal_14760), .Q (signal_14761) ) ;
    buf_clk cell_9881 ( .C (clk), .D (signal_14768), .Q (signal_14769) ) ;
    buf_clk cell_9889 ( .C (clk), .D (signal_14776), .Q (signal_14777) ) ;
    buf_clk cell_9897 ( .C (clk), .D (signal_14784), .Q (signal_14785) ) ;
    buf_clk cell_9905 ( .C (clk), .D (signal_14792), .Q (signal_14793) ) ;
    buf_clk cell_9913 ( .C (clk), .D (signal_14800), .Q (signal_14801) ) ;
    buf_clk cell_9921 ( .C (clk), .D (signal_14808), .Q (signal_14809) ) ;
    buf_clk cell_9929 ( .C (clk), .D (signal_14816), .Q (signal_14817) ) ;
    buf_clk cell_9937 ( .C (clk), .D (signal_14824), .Q (signal_14825) ) ;
    buf_clk cell_9945 ( .C (clk), .D (signal_14832), .Q (signal_14833) ) ;
    buf_clk cell_9953 ( .C (clk), .D (signal_14840), .Q (signal_14841) ) ;
    buf_clk cell_9961 ( .C (clk), .D (signal_14848), .Q (signal_14849) ) ;
    buf_clk cell_9969 ( .C (clk), .D (signal_14856), .Q (signal_14857) ) ;
    buf_clk cell_9977 ( .C (clk), .D (signal_14864), .Q (signal_14865) ) ;
    buf_clk cell_9985 ( .C (clk), .D (signal_14872), .Q (signal_14873) ) ;
    buf_clk cell_9993 ( .C (clk), .D (signal_14880), .Q (signal_14881) ) ;
    buf_clk cell_10001 ( .C (clk), .D (signal_14888), .Q (signal_14889) ) ;
    buf_clk cell_10009 ( .C (clk), .D (signal_14896), .Q (signal_14897) ) ;
    buf_clk cell_10017 ( .C (clk), .D (signal_14904), .Q (signal_14905) ) ;
    buf_clk cell_10025 ( .C (clk), .D (signal_14912), .Q (signal_14913) ) ;
    buf_clk cell_10033 ( .C (clk), .D (signal_14920), .Q (signal_14921) ) ;
    buf_clk cell_10041 ( .C (clk), .D (signal_14928), .Q (signal_14929) ) ;
    buf_clk cell_10049 ( .C (clk), .D (signal_14936), .Q (signal_14937) ) ;
    buf_clk cell_10057 ( .C (clk), .D (signal_14944), .Q (signal_14945) ) ;
    buf_clk cell_10065 ( .C (clk), .D (signal_14952), .Q (signal_14953) ) ;
    buf_clk cell_10073 ( .C (clk), .D (signal_14960), .Q (signal_14961) ) ;
    buf_clk cell_10081 ( .C (clk), .D (signal_14968), .Q (signal_14969) ) ;
    buf_clk cell_10089 ( .C (clk), .D (signal_14976), .Q (signal_14977) ) ;
    buf_clk cell_10097 ( .C (clk), .D (signal_14984), .Q (signal_14985) ) ;
    buf_clk cell_10105 ( .C (clk), .D (signal_14992), .Q (signal_14993) ) ;
    buf_clk cell_10113 ( .C (clk), .D (signal_15000), .Q (signal_15001) ) ;
    buf_clk cell_10121 ( .C (clk), .D (signal_15008), .Q (signal_15009) ) ;
    buf_clk cell_10129 ( .C (clk), .D (signal_15016), .Q (signal_15017) ) ;
    buf_clk cell_10137 ( .C (clk), .D (signal_15024), .Q (signal_15025) ) ;
    buf_clk cell_10145 ( .C (clk), .D (signal_15032), .Q (signal_15033) ) ;
    buf_clk cell_10153 ( .C (clk), .D (signal_15040), .Q (signal_15041) ) ;
    buf_clk cell_10161 ( .C (clk), .D (signal_15048), .Q (signal_15049) ) ;
    buf_clk cell_10169 ( .C (clk), .D (signal_15056), .Q (signal_15057) ) ;
    buf_clk cell_10177 ( .C (clk), .D (signal_15064), .Q (signal_15065) ) ;
    buf_clk cell_10185 ( .C (clk), .D (signal_15072), .Q (signal_15073) ) ;
    buf_clk cell_10193 ( .C (clk), .D (signal_15080), .Q (signal_15081) ) ;
    buf_clk cell_10201 ( .C (clk), .D (signal_15088), .Q (signal_15089) ) ;
    buf_clk cell_10209 ( .C (clk), .D (signal_15096), .Q (signal_15097) ) ;
    buf_clk cell_10217 ( .C (clk), .D (signal_15104), .Q (signal_15105) ) ;
    buf_clk cell_10225 ( .C (clk), .D (signal_15112), .Q (signal_15113) ) ;
    buf_clk cell_10233 ( .C (clk), .D (signal_15120), .Q (signal_15121) ) ;
    buf_clk cell_10241 ( .C (clk), .D (signal_15128), .Q (signal_15129) ) ;
    buf_clk cell_10249 ( .C (clk), .D (signal_15136), .Q (signal_15137) ) ;
    buf_clk cell_10257 ( .C (clk), .D (signal_15144), .Q (signal_15145) ) ;
    buf_clk cell_10265 ( .C (clk), .D (signal_15152), .Q (signal_15153) ) ;
    buf_clk cell_10273 ( .C (clk), .D (signal_15160), .Q (signal_15161) ) ;
    buf_clk cell_10281 ( .C (clk), .D (signal_15168), .Q (signal_15169) ) ;
    buf_clk cell_10289 ( .C (clk), .D (signal_15176), .Q (signal_15177) ) ;
    buf_clk cell_10297 ( .C (clk), .D (signal_15184), .Q (signal_15185) ) ;
    buf_clk cell_10305 ( .C (clk), .D (signal_15192), .Q (signal_15193) ) ;
    buf_clk cell_10313 ( .C (clk), .D (signal_15200), .Q (signal_15201) ) ;
    buf_clk cell_10321 ( .C (clk), .D (signal_15208), .Q (signal_15209) ) ;
    buf_clk cell_10329 ( .C (clk), .D (signal_15216), .Q (signal_15217) ) ;
    buf_clk cell_10337 ( .C (clk), .D (signal_15224), .Q (signal_15225) ) ;
    buf_clk cell_10345 ( .C (clk), .D (signal_15232), .Q (signal_15233) ) ;
    buf_clk cell_10353 ( .C (clk), .D (signal_15240), .Q (signal_15241) ) ;
    buf_clk cell_10361 ( .C (clk), .D (signal_15248), .Q (signal_15249) ) ;
    buf_clk cell_10369 ( .C (clk), .D (signal_15256), .Q (signal_15257) ) ;
    buf_clk cell_10377 ( .C (clk), .D (signal_15264), .Q (signal_15265) ) ;
    buf_clk cell_10385 ( .C (clk), .D (signal_15272), .Q (signal_15273) ) ;
    buf_clk cell_10393 ( .C (clk), .D (signal_15280), .Q (signal_15281) ) ;
    buf_clk cell_10401 ( .C (clk), .D (signal_15288), .Q (signal_15289) ) ;
    buf_clk cell_10409 ( .C (clk), .D (signal_15296), .Q (signal_15297) ) ;
    buf_clk cell_10417 ( .C (clk), .D (signal_15304), .Q (signal_15305) ) ;
    buf_clk cell_10425 ( .C (clk), .D (signal_15312), .Q (signal_15313) ) ;
    buf_clk cell_10433 ( .C (clk), .D (signal_15320), .Q (signal_15321) ) ;
    buf_clk cell_10441 ( .C (clk), .D (signal_15328), .Q (signal_15329) ) ;
    buf_clk cell_10449 ( .C (clk), .D (signal_15336), .Q (signal_15337) ) ;
    buf_clk cell_10457 ( .C (clk), .D (signal_15344), .Q (signal_15345) ) ;
    buf_clk cell_10465 ( .C (clk), .D (signal_15352), .Q (signal_15353) ) ;
    buf_clk cell_10473 ( .C (clk), .D (signal_15360), .Q (signal_15361) ) ;
    buf_clk cell_10481 ( .C (clk), .D (signal_15368), .Q (signal_15369) ) ;
    buf_clk cell_10489 ( .C (clk), .D (signal_15376), .Q (signal_15377) ) ;
    buf_clk cell_10497 ( .C (clk), .D (signal_15384), .Q (signal_15385) ) ;
    buf_clk cell_10505 ( .C (clk), .D (signal_15392), .Q (signal_15393) ) ;
    buf_clk cell_10513 ( .C (clk), .D (signal_15400), .Q (signal_15401) ) ;
    buf_clk cell_10521 ( .C (clk), .D (signal_15408), .Q (signal_15409) ) ;
    buf_clk cell_10529 ( .C (clk), .D (signal_15416), .Q (signal_15417) ) ;
    buf_clk cell_10537 ( .C (clk), .D (signal_15424), .Q (signal_15425) ) ;
    buf_clk cell_10545 ( .C (clk), .D (signal_15432), .Q (signal_15433) ) ;
    buf_clk cell_10553 ( .C (clk), .D (signal_15440), .Q (signal_15441) ) ;
    buf_clk cell_10561 ( .C (clk), .D (signal_15448), .Q (signal_15449) ) ;
    buf_clk cell_10569 ( .C (clk), .D (signal_15456), .Q (signal_15457) ) ;
    buf_clk cell_10577 ( .C (clk), .D (signal_15464), .Q (signal_15465) ) ;
    buf_clk cell_10585 ( .C (clk), .D (signal_15472), .Q (signal_15473) ) ;
    buf_clk cell_10593 ( .C (clk), .D (signal_15480), .Q (signal_15481) ) ;
    buf_clk cell_10601 ( .C (clk), .D (signal_15488), .Q (signal_15489) ) ;
    buf_clk cell_10609 ( .C (clk), .D (signal_15496), .Q (signal_15497) ) ;
    buf_clk cell_10617 ( .C (clk), .D (signal_15504), .Q (signal_15505) ) ;
    buf_clk cell_10625 ( .C (clk), .D (signal_15512), .Q (signal_15513) ) ;
    buf_clk cell_10633 ( .C (clk), .D (signal_15520), .Q (signal_15521) ) ;
    buf_clk cell_10641 ( .C (clk), .D (signal_15528), .Q (signal_15529) ) ;
    buf_clk cell_10649 ( .C (clk), .D (signal_15536), .Q (signal_15537) ) ;
    buf_clk cell_10657 ( .C (clk), .D (signal_15544), .Q (signal_15545) ) ;
    buf_clk cell_10665 ( .C (clk), .D (signal_15552), .Q (signal_15553) ) ;
    buf_clk cell_10673 ( .C (clk), .D (signal_15560), .Q (signal_15561) ) ;
    buf_clk cell_10681 ( .C (clk), .D (signal_15568), .Q (signal_15569) ) ;
    buf_clk cell_10689 ( .C (clk), .D (signal_15576), .Q (signal_15577) ) ;
    buf_clk cell_10697 ( .C (clk), .D (signal_15584), .Q (signal_15585) ) ;
    buf_clk cell_10705 ( .C (clk), .D (signal_15592), .Q (signal_15593) ) ;
    buf_clk cell_10713 ( .C (clk), .D (signal_15600), .Q (signal_15601) ) ;
    buf_clk cell_10721 ( .C (clk), .D (signal_15608), .Q (signal_15609) ) ;
    buf_clk cell_10729 ( .C (clk), .D (signal_15616), .Q (signal_15617) ) ;
    buf_clk cell_10737 ( .C (clk), .D (signal_15624), .Q (signal_15625) ) ;
    buf_clk cell_10745 ( .C (clk), .D (signal_15632), .Q (signal_15633) ) ;
    buf_clk cell_10753 ( .C (clk), .D (signal_15640), .Q (signal_15641) ) ;
    buf_clk cell_10761 ( .C (clk), .D (signal_15648), .Q (signal_15649) ) ;
    buf_clk cell_10769 ( .C (clk), .D (signal_15656), .Q (signal_15657) ) ;
    buf_clk cell_10777 ( .C (clk), .D (signal_15664), .Q (signal_15665) ) ;
    buf_clk cell_10785 ( .C (clk), .D (signal_15672), .Q (signal_15673) ) ;
    buf_clk cell_10793 ( .C (clk), .D (signal_15680), .Q (signal_15681) ) ;
    buf_clk cell_10801 ( .C (clk), .D (signal_15688), .Q (signal_15689) ) ;
    buf_clk cell_10809 ( .C (clk), .D (signal_15696), .Q (signal_15697) ) ;
    buf_clk cell_10817 ( .C (clk), .D (signal_15704), .Q (signal_15705) ) ;
    buf_clk cell_10825 ( .C (clk), .D (signal_15712), .Q (signal_15713) ) ;
    buf_clk cell_10833 ( .C (clk), .D (signal_15720), .Q (signal_15721) ) ;
    buf_clk cell_10841 ( .C (clk), .D (signal_15728), .Q (signal_15729) ) ;
    buf_clk cell_10849 ( .C (clk), .D (signal_15736), .Q (signal_15737) ) ;
    buf_clk cell_10857 ( .C (clk), .D (signal_15744), .Q (signal_15745) ) ;
    buf_clk cell_10865 ( .C (clk), .D (signal_15752), .Q (signal_15753) ) ;
    buf_clk cell_10873 ( .C (clk), .D (signal_15760), .Q (signal_15761) ) ;
    buf_clk cell_10881 ( .C (clk), .D (signal_15768), .Q (signal_15769) ) ;
    buf_clk cell_10889 ( .C (clk), .D (signal_15776), .Q (signal_15777) ) ;
    buf_clk cell_10897 ( .C (clk), .D (signal_15784), .Q (signal_15785) ) ;
    buf_clk cell_10905 ( .C (clk), .D (signal_15792), .Q (signal_15793) ) ;
    buf_clk cell_10913 ( .C (clk), .D (signal_15800), .Q (signal_15801) ) ;
    buf_clk cell_10921 ( .C (clk), .D (signal_15808), .Q (signal_15809) ) ;
    buf_clk cell_10929 ( .C (clk), .D (signal_15816), .Q (signal_15817) ) ;
    buf_clk cell_10937 ( .C (clk), .D (signal_15824), .Q (signal_15825) ) ;
    buf_clk cell_10945 ( .C (clk), .D (signal_15832), .Q (signal_15833) ) ;
    buf_clk cell_10953 ( .C (clk), .D (signal_15840), .Q (signal_15841) ) ;
    buf_clk cell_10961 ( .C (clk), .D (signal_15848), .Q (signal_15849) ) ;
    buf_clk cell_10969 ( .C (clk), .D (signal_15856), .Q (signal_15857) ) ;
    buf_clk cell_10977 ( .C (clk), .D (signal_15864), .Q (signal_15865) ) ;
    buf_clk cell_10985 ( .C (clk), .D (signal_15872), .Q (signal_15873) ) ;
    buf_clk cell_10993 ( .C (clk), .D (signal_15880), .Q (signal_15881) ) ;
    buf_clk cell_11001 ( .C (clk), .D (signal_15888), .Q (signal_15889) ) ;
    buf_clk cell_11009 ( .C (clk), .D (signal_15896), .Q (signal_15897) ) ;
    buf_clk cell_11017 ( .C (clk), .D (signal_15904), .Q (signal_15905) ) ;
    buf_clk cell_11025 ( .C (clk), .D (signal_15912), .Q (signal_15913) ) ;
    buf_clk cell_11033 ( .C (clk), .D (signal_15920), .Q (signal_15921) ) ;
    buf_clk cell_11041 ( .C (clk), .D (signal_15928), .Q (signal_15929) ) ;
    buf_clk cell_11049 ( .C (clk), .D (signal_15936), .Q (signal_15937) ) ;
    buf_clk cell_11057 ( .C (clk), .D (signal_15944), .Q (signal_15945) ) ;
    buf_clk cell_11065 ( .C (clk), .D (signal_15952), .Q (signal_15953) ) ;
    buf_clk cell_11073 ( .C (clk), .D (signal_15960), .Q (signal_15961) ) ;
    buf_clk cell_11081 ( .C (clk), .D (signal_15968), .Q (signal_15969) ) ;
    buf_clk cell_11089 ( .C (clk), .D (signal_15976), .Q (signal_15977) ) ;
    buf_clk cell_11097 ( .C (clk), .D (signal_15984), .Q (signal_15985) ) ;
    buf_clk cell_11105 ( .C (clk), .D (signal_15992), .Q (signal_15993) ) ;
    buf_clk cell_11113 ( .C (clk), .D (signal_16000), .Q (signal_16001) ) ;
    buf_clk cell_11121 ( .C (clk), .D (signal_16008), .Q (signal_16009) ) ;
    buf_clk cell_11129 ( .C (clk), .D (signal_16016), .Q (signal_16017) ) ;
    buf_clk cell_11137 ( .C (clk), .D (signal_16024), .Q (signal_16025) ) ;
    buf_clk cell_11145 ( .C (clk), .D (signal_16032), .Q (signal_16033) ) ;
    buf_clk cell_11153 ( .C (clk), .D (signal_16040), .Q (signal_16041) ) ;
    buf_clk cell_11161 ( .C (clk), .D (signal_16048), .Q (signal_16049) ) ;
    buf_clk cell_11169 ( .C (clk), .D (signal_16056), .Q (signal_16057) ) ;
    buf_clk cell_11177 ( .C (clk), .D (signal_16064), .Q (signal_16065) ) ;
    buf_clk cell_11185 ( .C (clk), .D (signal_16072), .Q (signal_16073) ) ;
    buf_clk cell_11193 ( .C (clk), .D (signal_16080), .Q (signal_16081) ) ;
    buf_clk cell_11201 ( .C (clk), .D (signal_16088), .Q (signal_16089) ) ;
    buf_clk cell_11209 ( .C (clk), .D (signal_16096), .Q (signal_16097) ) ;
    buf_clk cell_11217 ( .C (clk), .D (signal_16104), .Q (signal_16105) ) ;
    buf_clk cell_11225 ( .C (clk), .D (signal_16112), .Q (signal_16113) ) ;
    buf_clk cell_11233 ( .C (clk), .D (signal_16120), .Q (signal_16121) ) ;
    buf_clk cell_11241 ( .C (clk), .D (signal_16128), .Q (signal_16129) ) ;
    buf_clk cell_11249 ( .C (clk), .D (signal_16136), .Q (signal_16137) ) ;
    buf_clk cell_11257 ( .C (clk), .D (signal_16144), .Q (signal_16145) ) ;
    buf_clk cell_11265 ( .C (clk), .D (signal_16152), .Q (signal_16153) ) ;
    buf_clk cell_11273 ( .C (clk), .D (signal_16160), .Q (signal_16161) ) ;
    buf_clk cell_11281 ( .C (clk), .D (signal_16168), .Q (signal_16169) ) ;
    buf_clk cell_11289 ( .C (clk), .D (signal_16176), .Q (signal_16177) ) ;
    buf_clk cell_11297 ( .C (clk), .D (signal_16184), .Q (signal_16185) ) ;
    buf_clk cell_11305 ( .C (clk), .D (signal_16192), .Q (signal_16193) ) ;
    buf_clk cell_11313 ( .C (clk), .D (signal_16200), .Q (signal_16201) ) ;
    buf_clk cell_11321 ( .C (clk), .D (signal_16208), .Q (signal_16209) ) ;
    buf_clk cell_11329 ( .C (clk), .D (signal_16216), .Q (signal_16217) ) ;
    buf_clk cell_11337 ( .C (clk), .D (signal_16224), .Q (signal_16225) ) ;
    buf_clk cell_11345 ( .C (clk), .D (signal_16232), .Q (signal_16233) ) ;
    buf_clk cell_11353 ( .C (clk), .D (signal_16240), .Q (signal_16241) ) ;
    buf_clk cell_11361 ( .C (clk), .D (signal_16248), .Q (signal_16249) ) ;
    buf_clk cell_11369 ( .C (clk), .D (signal_16256), .Q (signal_16257) ) ;
    buf_clk cell_11377 ( .C (clk), .D (signal_16264), .Q (signal_16265) ) ;
    buf_clk cell_11385 ( .C (clk), .D (signal_16272), .Q (signal_16273) ) ;
    buf_clk cell_11393 ( .C (clk), .D (signal_16280), .Q (signal_16281) ) ;
    buf_clk cell_11401 ( .C (clk), .D (signal_16288), .Q (signal_16289) ) ;
    buf_clk cell_11409 ( .C (clk), .D (signal_16296), .Q (signal_16297) ) ;
    buf_clk cell_11417 ( .C (clk), .D (signal_16304), .Q (signal_16305) ) ;
    buf_clk cell_11425 ( .C (clk), .D (signal_16312), .Q (signal_16313) ) ;
    buf_clk cell_11433 ( .C (clk), .D (signal_16320), .Q (signal_16321) ) ;
    buf_clk cell_11441 ( .C (clk), .D (signal_16328), .Q (signal_16329) ) ;
    buf_clk cell_11449 ( .C (clk), .D (signal_16336), .Q (signal_16337) ) ;
    buf_clk cell_11457 ( .C (clk), .D (signal_16344), .Q (signal_16345) ) ;
    buf_clk cell_11465 ( .C (clk), .D (signal_16352), .Q (signal_16353) ) ;
    buf_clk cell_11473 ( .C (clk), .D (signal_16360), .Q (signal_16361) ) ;
    buf_clk cell_11481 ( .C (clk), .D (signal_16368), .Q (signal_16369) ) ;
    buf_clk cell_11489 ( .C (clk), .D (signal_16376), .Q (signal_16377) ) ;
    buf_clk cell_11497 ( .C (clk), .D (signal_16384), .Q (signal_16385) ) ;
    buf_clk cell_11505 ( .C (clk), .D (signal_16392), .Q (signal_16393) ) ;
    buf_clk cell_11513 ( .C (clk), .D (signal_16400), .Q (signal_16401) ) ;
    buf_clk cell_11521 ( .C (clk), .D (signal_16408), .Q (signal_16409) ) ;
    buf_clk cell_11529 ( .C (clk), .D (signal_16416), .Q (signal_16417) ) ;
    buf_clk cell_11537 ( .C (clk), .D (signal_16424), .Q (signal_16425) ) ;
    buf_clk cell_11545 ( .C (clk), .D (signal_16432), .Q (signal_16433) ) ;
    buf_clk cell_11553 ( .C (clk), .D (signal_16440), .Q (signal_16441) ) ;
    buf_clk cell_11561 ( .C (clk), .D (signal_16448), .Q (signal_16449) ) ;
    buf_clk cell_11569 ( .C (clk), .D (signal_16456), .Q (signal_16457) ) ;
    buf_clk cell_11577 ( .C (clk), .D (signal_16464), .Q (signal_16465) ) ;
    buf_clk cell_11585 ( .C (clk), .D (signal_16472), .Q (signal_16473) ) ;
    buf_clk cell_11593 ( .C (clk), .D (signal_16480), .Q (signal_16481) ) ;
    buf_clk cell_11601 ( .C (clk), .D (signal_16488), .Q (signal_16489) ) ;
    buf_clk cell_11609 ( .C (clk), .D (signal_16496), .Q (signal_16497) ) ;
    buf_clk cell_11617 ( .C (clk), .D (signal_16504), .Q (signal_16505) ) ;
    buf_clk cell_11625 ( .C (clk), .D (signal_16512), .Q (signal_16513) ) ;
    buf_clk cell_11633 ( .C (clk), .D (signal_16520), .Q (signal_16521) ) ;
    buf_clk cell_11641 ( .C (clk), .D (signal_16528), .Q (signal_16529) ) ;
    buf_clk cell_11649 ( .C (clk), .D (signal_16536), .Q (signal_16537) ) ;
    buf_clk cell_11657 ( .C (clk), .D (signal_16544), .Q (signal_16545) ) ;
    buf_clk cell_11665 ( .C (clk), .D (signal_16552), .Q (signal_16553) ) ;
    buf_clk cell_11673 ( .C (clk), .D (signal_16560), .Q (signal_16561) ) ;
    buf_clk cell_11681 ( .C (clk), .D (signal_16568), .Q (signal_16569) ) ;
    buf_clk cell_11689 ( .C (clk), .D (signal_16576), .Q (signal_16577) ) ;
    buf_clk cell_11697 ( .C (clk), .D (signal_16584), .Q (signal_16585) ) ;
    buf_clk cell_11705 ( .C (clk), .D (signal_16592), .Q (signal_16593) ) ;
    buf_clk cell_11713 ( .C (clk), .D (signal_16600), .Q (signal_16601) ) ;
    buf_clk cell_11721 ( .C (clk), .D (signal_16608), .Q (signal_16609) ) ;
    buf_clk cell_11729 ( .C (clk), .D (signal_16616), .Q (signal_16617) ) ;
    buf_clk cell_11737 ( .C (clk), .D (signal_16624), .Q (signal_16625) ) ;
    buf_clk cell_11745 ( .C (clk), .D (signal_16632), .Q (signal_16633) ) ;
    buf_clk cell_11753 ( .C (clk), .D (signal_16640), .Q (signal_16641) ) ;
    buf_clk cell_11761 ( .C (clk), .D (signal_16648), .Q (signal_16649) ) ;
    buf_clk cell_11769 ( .C (clk), .D (signal_16656), .Q (signal_16657) ) ;
    buf_clk cell_11777 ( .C (clk), .D (signal_16664), .Q (signal_16665) ) ;
    buf_clk cell_11785 ( .C (clk), .D (signal_16672), .Q (signal_16673) ) ;
    buf_clk cell_11793 ( .C (clk), .D (signal_16680), .Q (signal_16681) ) ;
    buf_clk cell_11801 ( .C (clk), .D (signal_16688), .Q (signal_16689) ) ;
    buf_clk cell_11809 ( .C (clk), .D (signal_16696), .Q (signal_16697) ) ;
    buf_clk cell_11817 ( .C (clk), .D (signal_16704), .Q (signal_16705) ) ;
    buf_clk cell_11825 ( .C (clk), .D (signal_16712), .Q (signal_16713) ) ;
    buf_clk cell_11833 ( .C (clk), .D (signal_16720), .Q (signal_16721) ) ;
    buf_clk cell_11841 ( .C (clk), .D (signal_16728), .Q (signal_16729) ) ;
    buf_clk cell_11849 ( .C (clk), .D (signal_16736), .Q (signal_16737) ) ;
    buf_clk cell_11857 ( .C (clk), .D (signal_16744), .Q (signal_16745) ) ;
    buf_clk cell_11865 ( .C (clk), .D (signal_16752), .Q (signal_16753) ) ;
    buf_clk cell_11873 ( .C (clk), .D (signal_16760), .Q (signal_16761) ) ;
    buf_clk cell_11881 ( .C (clk), .D (signal_16768), .Q (signal_16769) ) ;
    buf_clk cell_11889 ( .C (clk), .D (signal_16776), .Q (signal_16777) ) ;
    buf_clk cell_11897 ( .C (clk), .D (signal_16784), .Q (signal_16785) ) ;
    buf_clk cell_11905 ( .C (clk), .D (signal_16792), .Q (signal_16793) ) ;
    buf_clk cell_11913 ( .C (clk), .D (signal_16800), .Q (signal_16801) ) ;
    buf_clk cell_11921 ( .C (clk), .D (signal_16808), .Q (signal_16809) ) ;
    buf_clk cell_11929 ( .C (clk), .D (signal_16816), .Q (signal_16817) ) ;
    buf_clk cell_11937 ( .C (clk), .D (signal_16824), .Q (signal_16825) ) ;
    buf_clk cell_11945 ( .C (clk), .D (signal_16832), .Q (signal_16833) ) ;
    buf_clk cell_11953 ( .C (clk), .D (signal_16840), .Q (signal_16841) ) ;
    buf_clk cell_11961 ( .C (clk), .D (signal_16848), .Q (signal_16849) ) ;
    buf_clk cell_11969 ( .C (clk), .D (signal_16856), .Q (signal_16857) ) ;
    buf_clk cell_11977 ( .C (clk), .D (signal_16864), .Q (signal_16865) ) ;
    buf_clk cell_11985 ( .C (clk), .D (signal_16872), .Q (signal_16873) ) ;
    buf_clk cell_11993 ( .C (clk), .D (signal_16880), .Q (signal_16881) ) ;
    buf_clk cell_12001 ( .C (clk), .D (signal_16888), .Q (signal_16889) ) ;
    buf_clk cell_12009 ( .C (clk), .D (signal_16896), .Q (signal_16897) ) ;
    buf_clk cell_12017 ( .C (clk), .D (signal_16904), .Q (signal_16905) ) ;
    buf_clk cell_12025 ( .C (clk), .D (signal_16912), .Q (signal_16913) ) ;
    buf_clk cell_12033 ( .C (clk), .D (signal_16920), .Q (signal_16921) ) ;
    buf_clk cell_12041 ( .C (clk), .D (signal_16928), .Q (signal_16929) ) ;
    buf_clk cell_12049 ( .C (clk), .D (signal_16936), .Q (signal_16937) ) ;
    buf_clk cell_12057 ( .C (clk), .D (signal_16944), .Q (signal_16945) ) ;
    buf_clk cell_12065 ( .C (clk), .D (signal_16952), .Q (signal_16953) ) ;
    buf_clk cell_12073 ( .C (clk), .D (signal_16960), .Q (signal_16961) ) ;
    buf_clk cell_12081 ( .C (clk), .D (signal_16968), .Q (signal_16969) ) ;
    buf_clk cell_12089 ( .C (clk), .D (signal_16976), .Q (signal_16977) ) ;
    buf_clk cell_12097 ( .C (clk), .D (signal_16984), .Q (signal_16985) ) ;
    buf_clk cell_12105 ( .C (clk), .D (signal_16992), .Q (signal_16993) ) ;
    buf_clk cell_12113 ( .C (clk), .D (signal_17000), .Q (signal_17001) ) ;
    buf_clk cell_12121 ( .C (clk), .D (signal_17008), .Q (signal_17009) ) ;
    buf_clk cell_12129 ( .C (clk), .D (signal_17016), .Q (signal_17017) ) ;
    buf_clk cell_12137 ( .C (clk), .D (signal_17024), .Q (signal_17025) ) ;
    buf_clk cell_12145 ( .C (clk), .D (signal_17032), .Q (signal_17033) ) ;
    buf_clk cell_12153 ( .C (clk), .D (signal_17040), .Q (signal_17041) ) ;
    buf_clk cell_12161 ( .C (clk), .D (signal_17048), .Q (signal_17049) ) ;
    buf_clk cell_12169 ( .C (clk), .D (signal_17056), .Q (signal_17057) ) ;
    buf_clk cell_12177 ( .C (clk), .D (signal_17064), .Q (signal_17065) ) ;
    buf_clk cell_12185 ( .C (clk), .D (signal_17072), .Q (signal_17073) ) ;
    buf_clk cell_12193 ( .C (clk), .D (signal_17080), .Q (signal_17081) ) ;
    buf_clk cell_12201 ( .C (clk), .D (signal_17088), .Q (signal_17089) ) ;
    buf_clk cell_12209 ( .C (clk), .D (signal_17096), .Q (signal_17097) ) ;
    buf_clk cell_12217 ( .C (clk), .D (signal_17104), .Q (signal_17105) ) ;
    buf_clk cell_12225 ( .C (clk), .D (signal_17112), .Q (signal_17113) ) ;
    buf_clk cell_12233 ( .C (clk), .D (signal_17120), .Q (signal_17121) ) ;
    buf_clk cell_12241 ( .C (clk), .D (signal_17128), .Q (signal_17129) ) ;
    buf_clk cell_12249 ( .C (clk), .D (signal_17136), .Q (signal_17137) ) ;
    buf_clk cell_12257 ( .C (clk), .D (signal_17144), .Q (signal_17145) ) ;
    buf_clk cell_12265 ( .C (clk), .D (signal_17152), .Q (signal_17153) ) ;
    buf_clk cell_12273 ( .C (clk), .D (signal_17160), .Q (signal_17161) ) ;
    buf_clk cell_12281 ( .C (clk), .D (signal_17168), .Q (signal_17169) ) ;
    buf_clk cell_12289 ( .C (clk), .D (signal_17176), .Q (signal_17177) ) ;
    buf_clk cell_12297 ( .C (clk), .D (signal_17184), .Q (signal_17185) ) ;
    buf_clk cell_12305 ( .C (clk), .D (signal_17192), .Q (signal_17193) ) ;
    buf_clk cell_12313 ( .C (clk), .D (signal_17200), .Q (signal_17201) ) ;
    buf_clk cell_12321 ( .C (clk), .D (signal_17208), .Q (signal_17209) ) ;
    buf_clk cell_12329 ( .C (clk), .D (signal_17216), .Q (signal_17217) ) ;
    buf_clk cell_12337 ( .C (clk), .D (signal_17224), .Q (signal_17225) ) ;
    buf_clk cell_12345 ( .C (clk), .D (signal_17232), .Q (signal_17233) ) ;
    buf_clk cell_12353 ( .C (clk), .D (signal_17240), .Q (signal_17241) ) ;
    buf_clk cell_12361 ( .C (clk), .D (signal_17248), .Q (signal_17249) ) ;
    buf_clk cell_12369 ( .C (clk), .D (signal_17256), .Q (signal_17257) ) ;
    buf_clk cell_12377 ( .C (clk), .D (signal_17264), .Q (signal_17265) ) ;
    buf_clk cell_12385 ( .C (clk), .D (signal_17272), .Q (signal_17273) ) ;
    buf_clk cell_12393 ( .C (clk), .D (signal_17280), .Q (signal_17281) ) ;
    buf_clk cell_12401 ( .C (clk), .D (signal_17288), .Q (signal_17289) ) ;
    buf_clk cell_12409 ( .C (clk), .D (signal_17296), .Q (signal_17297) ) ;
    buf_clk cell_12417 ( .C (clk), .D (signal_17304), .Q (signal_17305) ) ;
    buf_clk cell_12425 ( .C (clk), .D (signal_17312), .Q (signal_17313) ) ;
    buf_clk cell_12433 ( .C (clk), .D (signal_17320), .Q (signal_17321) ) ;
    buf_clk cell_12441 ( .C (clk), .D (signal_17328), .Q (signal_17329) ) ;
    buf_clk cell_12449 ( .C (clk), .D (signal_17336), .Q (signal_17337) ) ;
    buf_clk cell_12457 ( .C (clk), .D (signal_17344), .Q (signal_17345) ) ;
    buf_clk cell_12465 ( .C (clk), .D (signal_17352), .Q (signal_17353) ) ;
    buf_clk cell_12473 ( .C (clk), .D (signal_17360), .Q (signal_17361) ) ;
    buf_clk cell_12481 ( .C (clk), .D (signal_17368), .Q (signal_17369) ) ;
    buf_clk cell_12489 ( .C (clk), .D (signal_17376), .Q (signal_17377) ) ;
    buf_clk cell_12497 ( .C (clk), .D (signal_17384), .Q (signal_17385) ) ;
    buf_clk cell_12505 ( .C (clk), .D (signal_17392), .Q (signal_17393) ) ;
    buf_clk cell_12513 ( .C (clk), .D (signal_17400), .Q (signal_17401) ) ;
    buf_clk cell_12521 ( .C (clk), .D (signal_17408), .Q (signal_17409) ) ;
    buf_clk cell_12529 ( .C (clk), .D (signal_17416), .Q (signal_17417) ) ;
    buf_clk cell_12537 ( .C (clk), .D (signal_17424), .Q (signal_17425) ) ;
    buf_clk cell_12545 ( .C (clk), .D (signal_17432), .Q (signal_17433) ) ;
    buf_clk cell_12553 ( .C (clk), .D (signal_17440), .Q (signal_17441) ) ;
    buf_clk cell_12561 ( .C (clk), .D (signal_17448), .Q (signal_17449) ) ;
    buf_clk cell_12569 ( .C (clk), .D (signal_17456), .Q (signal_17457) ) ;
    buf_clk cell_12577 ( .C (clk), .D (signal_17464), .Q (signal_17465) ) ;
    buf_clk cell_12585 ( .C (clk), .D (signal_17472), .Q (signal_17473) ) ;
    buf_clk cell_12593 ( .C (clk), .D (signal_17480), .Q (signal_17481) ) ;
    buf_clk cell_12601 ( .C (clk), .D (signal_17488), .Q (signal_17489) ) ;
    buf_clk cell_12609 ( .C (clk), .D (signal_17496), .Q (signal_17497) ) ;
    buf_clk cell_12617 ( .C (clk), .D (signal_17504), .Q (signal_17505) ) ;
    buf_clk cell_12625 ( .C (clk), .D (signal_17512), .Q (signal_17513) ) ;
    buf_clk cell_12633 ( .C (clk), .D (signal_17520), .Q (signal_17521) ) ;
    buf_clk cell_12641 ( .C (clk), .D (signal_17528), .Q (signal_17529) ) ;
    buf_clk cell_12649 ( .C (clk), .D (signal_17536), .Q (signal_17537) ) ;
    buf_clk cell_12657 ( .C (clk), .D (signal_17544), .Q (signal_17545) ) ;
    buf_clk cell_12665 ( .C (clk), .D (signal_17552), .Q (signal_17553) ) ;
    buf_clk cell_12673 ( .C (clk), .D (signal_17560), .Q (signal_17561) ) ;
    buf_clk cell_12681 ( .C (clk), .D (signal_17568), .Q (signal_17569) ) ;
    buf_clk cell_12689 ( .C (clk), .D (signal_17576), .Q (signal_17577) ) ;
    buf_clk cell_12697 ( .C (clk), .D (signal_17584), .Q (signal_17585) ) ;
    buf_clk cell_12705 ( .C (clk), .D (signal_17592), .Q (signal_17593) ) ;
    buf_clk cell_12713 ( .C (clk), .D (signal_17600), .Q (signal_17601) ) ;
    buf_clk cell_12721 ( .C (clk), .D (signal_17608), .Q (signal_17609) ) ;
    buf_clk cell_12729 ( .C (clk), .D (signal_17616), .Q (signal_17617) ) ;
    buf_clk cell_12737 ( .C (clk), .D (signal_17624), .Q (signal_17625) ) ;
    buf_clk cell_12745 ( .C (clk), .D (signal_17632), .Q (signal_17633) ) ;
    buf_clk cell_12753 ( .C (clk), .D (signal_17640), .Q (signal_17641) ) ;
    buf_clk cell_12761 ( .C (clk), .D (signal_17648), .Q (signal_17649) ) ;
    buf_clk cell_12769 ( .C (clk), .D (signal_17656), .Q (signal_17657) ) ;
    buf_clk cell_12777 ( .C (clk), .D (signal_17664), .Q (signal_17665) ) ;
    buf_clk cell_12785 ( .C (clk), .D (signal_17672), .Q (signal_17673) ) ;
    buf_clk cell_12793 ( .C (clk), .D (signal_17680), .Q (signal_17681) ) ;
    buf_clk cell_12801 ( .C (clk), .D (signal_17688), .Q (signal_17689) ) ;
    buf_clk cell_12809 ( .C (clk), .D (signal_17696), .Q (signal_17697) ) ;
    buf_clk cell_12817 ( .C (clk), .D (signal_17704), .Q (signal_17705) ) ;
    buf_clk cell_12825 ( .C (clk), .D (signal_17712), .Q (signal_17713) ) ;
    buf_clk cell_12833 ( .C (clk), .D (signal_17720), .Q (signal_17721) ) ;
    buf_clk cell_12841 ( .C (clk), .D (signal_17728), .Q (signal_17729) ) ;
    buf_clk cell_12849 ( .C (clk), .D (signal_17736), .Q (signal_17737) ) ;
    buf_clk cell_12857 ( .C (clk), .D (signal_17744), .Q (signal_17745) ) ;
    buf_clk cell_12865 ( .C (clk), .D (signal_17752), .Q (signal_17753) ) ;
    buf_clk cell_12873 ( .C (clk), .D (signal_17760), .Q (signal_17761) ) ;
    buf_clk cell_12881 ( .C (clk), .D (signal_17768), .Q (signal_17769) ) ;
    buf_clk cell_12889 ( .C (clk), .D (signal_17776), .Q (signal_17777) ) ;
    buf_clk cell_12897 ( .C (clk), .D (signal_17784), .Q (signal_17785) ) ;
    buf_clk cell_12905 ( .C (clk), .D (signal_17792), .Q (signal_17793) ) ;
    buf_clk cell_12913 ( .C (clk), .D (signal_17800), .Q (signal_17801) ) ;
    buf_clk cell_12921 ( .C (clk), .D (signal_17808), .Q (signal_17809) ) ;
    buf_clk cell_12929 ( .C (clk), .D (signal_17816), .Q (signal_17817) ) ;
    buf_clk cell_12937 ( .C (clk), .D (signal_17824), .Q (signal_17825) ) ;
    buf_clk cell_12945 ( .C (clk), .D (signal_17832), .Q (signal_17833) ) ;
    buf_clk cell_12953 ( .C (clk), .D (signal_17840), .Q (signal_17841) ) ;
    buf_clk cell_12961 ( .C (clk), .D (signal_17848), .Q (signal_17849) ) ;
    buf_clk cell_12969 ( .C (clk), .D (signal_17856), .Q (signal_17857) ) ;
    buf_clk cell_12977 ( .C (clk), .D (signal_17864), .Q (signal_17865) ) ;
    buf_clk cell_12985 ( .C (clk), .D (signal_17872), .Q (signal_17873) ) ;
    buf_clk cell_12993 ( .C (clk), .D (signal_17880), .Q (signal_17881) ) ;
    buf_clk cell_13001 ( .C (clk), .D (signal_17888), .Q (signal_17889) ) ;
    buf_clk cell_13009 ( .C (clk), .D (signal_17896), .Q (signal_17897) ) ;
    buf_clk cell_13017 ( .C (clk), .D (signal_17904), .Q (signal_17905) ) ;
    buf_clk cell_13025 ( .C (clk), .D (signal_17912), .Q (signal_17913) ) ;
    buf_clk cell_13033 ( .C (clk), .D (signal_17920), .Q (signal_17921) ) ;
    buf_clk cell_13041 ( .C (clk), .D (signal_17928), .Q (signal_17929) ) ;
    buf_clk cell_13049 ( .C (clk), .D (signal_17936), .Q (signal_17937) ) ;
    buf_clk cell_13057 ( .C (clk), .D (signal_17944), .Q (signal_17945) ) ;
    buf_clk cell_13065 ( .C (clk), .D (signal_17952), .Q (signal_17953) ) ;
    buf_clk cell_13073 ( .C (clk), .D (signal_17960), .Q (signal_17961) ) ;
    buf_clk cell_13081 ( .C (clk), .D (signal_17968), .Q (signal_17969) ) ;
    buf_clk cell_13089 ( .C (clk), .D (signal_17976), .Q (signal_17977) ) ;
    buf_clk cell_13097 ( .C (clk), .D (signal_17984), .Q (signal_17985) ) ;
    buf_clk cell_13105 ( .C (clk), .D (signal_17992), .Q (signal_17993) ) ;
    buf_clk cell_13113 ( .C (clk), .D (signal_18000), .Q (signal_18001) ) ;
    buf_clk cell_13121 ( .C (clk), .D (signal_18008), .Q (signal_18009) ) ;
    buf_clk cell_13129 ( .C (clk), .D (signal_18016), .Q (signal_18017) ) ;
    buf_clk cell_13137 ( .C (clk), .D (signal_18024), .Q (signal_18025) ) ;
    buf_clk cell_13145 ( .C (clk), .D (signal_18032), .Q (signal_18033) ) ;
    buf_clk cell_13153 ( .C (clk), .D (signal_18040), .Q (signal_18041) ) ;
    buf_clk cell_13161 ( .C (clk), .D (signal_18048), .Q (signal_18049) ) ;
    buf_clk cell_13169 ( .C (clk), .D (signal_18056), .Q (signal_18057) ) ;
    buf_clk cell_13177 ( .C (clk), .D (signal_18064), .Q (signal_18065) ) ;
    buf_clk cell_13185 ( .C (clk), .D (signal_18072), .Q (signal_18073) ) ;
    buf_clk cell_13193 ( .C (clk), .D (signal_18080), .Q (signal_18081) ) ;
    buf_clk cell_13201 ( .C (clk), .D (signal_18088), .Q (signal_18089) ) ;
    buf_clk cell_13209 ( .C (clk), .D (signal_18096), .Q (signal_18097) ) ;
    buf_clk cell_13217 ( .C (clk), .D (signal_18104), .Q (signal_18105) ) ;
    buf_clk cell_13225 ( .C (clk), .D (signal_18112), .Q (signal_18113) ) ;
    buf_clk cell_13233 ( .C (clk), .D (signal_18120), .Q (signal_18121) ) ;
    buf_clk cell_13241 ( .C (clk), .D (signal_18128), .Q (signal_18129) ) ;
    buf_clk cell_13249 ( .C (clk), .D (signal_18136), .Q (signal_18137) ) ;
    buf_clk cell_13257 ( .C (clk), .D (signal_18144), .Q (signal_18145) ) ;
    buf_clk cell_13265 ( .C (clk), .D (signal_18152), .Q (signal_18153) ) ;
    buf_clk cell_13273 ( .C (clk), .D (signal_18160), .Q (signal_18161) ) ;
    buf_clk cell_13281 ( .C (clk), .D (signal_18168), .Q (signal_18169) ) ;
    buf_clk cell_13287 ( .C (clk), .D (signal_18174), .Q (signal_18175) ) ;
    buf_clk cell_13293 ( .C (clk), .D (signal_18180), .Q (signal_18181) ) ;
    buf_clk cell_13299 ( .C (clk), .D (signal_18186), .Q (signal_18187) ) ;
    buf_clk cell_13305 ( .C (clk), .D (signal_18192), .Q (signal_18193) ) ;
    buf_clk cell_13311 ( .C (clk), .D (signal_18198), .Q (signal_18199) ) ;
    buf_clk cell_13317 ( .C (clk), .D (signal_18204), .Q (signal_18205) ) ;
    buf_clk cell_13323 ( .C (clk), .D (signal_18210), .Q (signal_18211) ) ;
    buf_clk cell_13329 ( .C (clk), .D (signal_18216), .Q (signal_18217) ) ;
    buf_clk cell_13335 ( .C (clk), .D (signal_18222), .Q (signal_18223) ) ;
    buf_clk cell_13341 ( .C (clk), .D (signal_18228), .Q (signal_18229) ) ;
    buf_clk cell_13347 ( .C (clk), .D (signal_18234), .Q (signal_18235) ) ;
    buf_clk cell_13353 ( .C (clk), .D (signal_18240), .Q (signal_18241) ) ;
    buf_clk cell_13359 ( .C (clk), .D (signal_18246), .Q (signal_18247) ) ;
    buf_clk cell_13365 ( .C (clk), .D (signal_18252), .Q (signal_18253) ) ;
    buf_clk cell_13371 ( .C (clk), .D (signal_18258), .Q (signal_18259) ) ;
    buf_clk cell_13377 ( .C (clk), .D (signal_18264), .Q (signal_18265) ) ;
    buf_clk cell_13383 ( .C (clk), .D (signal_18270), .Q (signal_18271) ) ;
    buf_clk cell_13389 ( .C (clk), .D (signal_18276), .Q (signal_18277) ) ;
    buf_clk cell_13395 ( .C (clk), .D (signal_18282), .Q (signal_18283) ) ;
    buf_clk cell_13401 ( .C (clk), .D (signal_18288), .Q (signal_18289) ) ;
    buf_clk cell_13407 ( .C (clk), .D (signal_18294), .Q (signal_18295) ) ;
    buf_clk cell_13413 ( .C (clk), .D (signal_18300), .Q (signal_18301) ) ;
    buf_clk cell_13419 ( .C (clk), .D (signal_18306), .Q (signal_18307) ) ;
    buf_clk cell_13425 ( .C (clk), .D (signal_18312), .Q (signal_18313) ) ;
    buf_clk cell_13431 ( .C (clk), .D (signal_18318), .Q (signal_18319) ) ;
    buf_clk cell_13437 ( .C (clk), .D (signal_18324), .Q (signal_18325) ) ;
    buf_clk cell_13443 ( .C (clk), .D (signal_18330), .Q (signal_18331) ) ;
    buf_clk cell_13449 ( .C (clk), .D (signal_18336), .Q (signal_18337) ) ;
    buf_clk cell_13455 ( .C (clk), .D (signal_18342), .Q (signal_18343) ) ;
    buf_clk cell_13461 ( .C (clk), .D (signal_18348), .Q (signal_18349) ) ;
    buf_clk cell_13467 ( .C (clk), .D (signal_18354), .Q (signal_18355) ) ;
    buf_clk cell_13473 ( .C (clk), .D (signal_18360), .Q (signal_18361) ) ;
    buf_clk cell_13479 ( .C (clk), .D (signal_18366), .Q (signal_18367) ) ;
    buf_clk cell_13485 ( .C (clk), .D (signal_18372), .Q (signal_18373) ) ;
    buf_clk cell_13491 ( .C (clk), .D (signal_18378), .Q (signal_18379) ) ;
    buf_clk cell_13497 ( .C (clk), .D (signal_18384), .Q (signal_18385) ) ;
    buf_clk cell_13503 ( .C (clk), .D (signal_18390), .Q (signal_18391) ) ;
    buf_clk cell_13509 ( .C (clk), .D (signal_18396), .Q (signal_18397) ) ;
    buf_clk cell_13515 ( .C (clk), .D (signal_18402), .Q (signal_18403) ) ;
    buf_clk cell_13521 ( .C (clk), .D (signal_18408), .Q (signal_18409) ) ;
    buf_clk cell_13527 ( .C (clk), .D (signal_18414), .Q (signal_18415) ) ;
    buf_clk cell_13533 ( .C (clk), .D (signal_18420), .Q (signal_18421) ) ;
    buf_clk cell_13539 ( .C (clk), .D (signal_18426), .Q (signal_18427) ) ;
    buf_clk cell_13545 ( .C (clk), .D (signal_18432), .Q (signal_18433) ) ;
    buf_clk cell_13551 ( .C (clk), .D (signal_18438), .Q (signal_18439) ) ;
    buf_clk cell_13557 ( .C (clk), .D (signal_18444), .Q (signal_18445) ) ;
    buf_clk cell_13563 ( .C (clk), .D (signal_18450), .Q (signal_18451) ) ;
    buf_clk cell_13569 ( .C (clk), .D (signal_18456), .Q (signal_18457) ) ;
    buf_clk cell_13575 ( .C (clk), .D (signal_18462), .Q (signal_18463) ) ;
    buf_clk cell_13581 ( .C (clk), .D (signal_18468), .Q (signal_18469) ) ;
    buf_clk cell_13587 ( .C (clk), .D (signal_18474), .Q (signal_18475) ) ;
    buf_clk cell_13593 ( .C (clk), .D (signal_18480), .Q (signal_18481) ) ;
    buf_clk cell_13599 ( .C (clk), .D (signal_18486), .Q (signal_18487) ) ;
    buf_clk cell_13605 ( .C (clk), .D (signal_18492), .Q (signal_18493) ) ;
    buf_clk cell_13611 ( .C (clk), .D (signal_18498), .Q (signal_18499) ) ;
    buf_clk cell_13617 ( .C (clk), .D (signal_18504), .Q (signal_18505) ) ;
    buf_clk cell_13623 ( .C (clk), .D (signal_18510), .Q (signal_18511) ) ;
    buf_clk cell_13629 ( .C (clk), .D (signal_18516), .Q (signal_18517) ) ;
    buf_clk cell_13635 ( .C (clk), .D (signal_18522), .Q (signal_18523) ) ;
    buf_clk cell_13641 ( .C (clk), .D (signal_18528), .Q (signal_18529) ) ;
    buf_clk cell_13647 ( .C (clk), .D (signal_18534), .Q (signal_18535) ) ;
    buf_clk cell_13653 ( .C (clk), .D (signal_18540), .Q (signal_18541) ) ;
    buf_clk cell_13659 ( .C (clk), .D (signal_18546), .Q (signal_18547) ) ;
    buf_clk cell_13665 ( .C (clk), .D (signal_18552), .Q (signal_18553) ) ;
    buf_clk cell_13671 ( .C (clk), .D (signal_18558), .Q (signal_18559) ) ;
    buf_clk cell_13677 ( .C (clk), .D (signal_18564), .Q (signal_18565) ) ;
    buf_clk cell_13683 ( .C (clk), .D (signal_18570), .Q (signal_18571) ) ;
    buf_clk cell_13689 ( .C (clk), .D (signal_18576), .Q (signal_18577) ) ;
    buf_clk cell_13695 ( .C (clk), .D (signal_18582), .Q (signal_18583) ) ;
    buf_clk cell_13701 ( .C (clk), .D (signal_18588), .Q (signal_18589) ) ;
    buf_clk cell_13707 ( .C (clk), .D (signal_18594), .Q (signal_18595) ) ;
    buf_clk cell_13713 ( .C (clk), .D (signal_18600), .Q (signal_18601) ) ;
    buf_clk cell_13719 ( .C (clk), .D (signal_18606), .Q (signal_18607) ) ;
    buf_clk cell_13725 ( .C (clk), .D (signal_18612), .Q (signal_18613) ) ;
    buf_clk cell_13731 ( .C (clk), .D (signal_18618), .Q (signal_18619) ) ;
    buf_clk cell_13737 ( .C (clk), .D (signal_18624), .Q (signal_18625) ) ;
    buf_clk cell_13743 ( .C (clk), .D (signal_18630), .Q (signal_18631) ) ;
    buf_clk cell_13749 ( .C (clk), .D (signal_18636), .Q (signal_18637) ) ;
    buf_clk cell_13755 ( .C (clk), .D (signal_18642), .Q (signal_18643) ) ;
    buf_clk cell_13761 ( .C (clk), .D (signal_18648), .Q (signal_18649) ) ;
    buf_clk cell_13767 ( .C (clk), .D (signal_18654), .Q (signal_18655) ) ;
    buf_clk cell_13773 ( .C (clk), .D (signal_18660), .Q (signal_18661) ) ;
    buf_clk cell_13779 ( .C (clk), .D (signal_18666), .Q (signal_18667) ) ;
    buf_clk cell_13785 ( .C (clk), .D (signal_18672), .Q (signal_18673) ) ;
    buf_clk cell_13791 ( .C (clk), .D (signal_18678), .Q (signal_18679) ) ;
    buf_clk cell_13797 ( .C (clk), .D (signal_18684), .Q (signal_18685) ) ;
    buf_clk cell_13803 ( .C (clk), .D (signal_18690), .Q (signal_18691) ) ;
    buf_clk cell_13809 ( .C (clk), .D (signal_18696), .Q (signal_18697) ) ;
    buf_clk cell_13815 ( .C (clk), .D (signal_18702), .Q (signal_18703) ) ;
    buf_clk cell_13821 ( .C (clk), .D (signal_18708), .Q (signal_18709) ) ;
    buf_clk cell_13827 ( .C (clk), .D (signal_18714), .Q (signal_18715) ) ;
    buf_clk cell_13833 ( .C (clk), .D (signal_18720), .Q (signal_18721) ) ;
    buf_clk cell_13839 ( .C (clk), .D (signal_18726), .Q (signal_18727) ) ;
    buf_clk cell_13845 ( .C (clk), .D (signal_18732), .Q (signal_18733) ) ;
    buf_clk cell_13851 ( .C (clk), .D (signal_18738), .Q (signal_18739) ) ;
    buf_clk cell_13857 ( .C (clk), .D (signal_18744), .Q (signal_18745) ) ;
    buf_clk cell_13863 ( .C (clk), .D (signal_18750), .Q (signal_18751) ) ;
    buf_clk cell_13869 ( .C (clk), .D (signal_18756), .Q (signal_18757) ) ;
    buf_clk cell_13875 ( .C (clk), .D (signal_18762), .Q (signal_18763) ) ;
    buf_clk cell_13881 ( .C (clk), .D (signal_18768), .Q (signal_18769) ) ;
    buf_clk cell_13887 ( .C (clk), .D (signal_18774), .Q (signal_18775) ) ;
    buf_clk cell_13893 ( .C (clk), .D (signal_18780), .Q (signal_18781) ) ;
    buf_clk cell_13899 ( .C (clk), .D (signal_18786), .Q (signal_18787) ) ;
    buf_clk cell_13905 ( .C (clk), .D (signal_18792), .Q (signal_18793) ) ;
    buf_clk cell_13911 ( .C (clk), .D (signal_18798), .Q (signal_18799) ) ;
    buf_clk cell_13917 ( .C (clk), .D (signal_18804), .Q (signal_18805) ) ;
    buf_clk cell_13923 ( .C (clk), .D (signal_18810), .Q (signal_18811) ) ;
    buf_clk cell_13929 ( .C (clk), .D (signal_18816), .Q (signal_18817) ) ;
    buf_clk cell_13935 ( .C (clk), .D (signal_18822), .Q (signal_18823) ) ;
    buf_clk cell_13941 ( .C (clk), .D (signal_18828), .Q (signal_18829) ) ;
    buf_clk cell_13947 ( .C (clk), .D (signal_18834), .Q (signal_18835) ) ;
    buf_clk cell_13953 ( .C (clk), .D (signal_18840), .Q (signal_18841) ) ;
    buf_clk cell_13959 ( .C (clk), .D (signal_18846), .Q (signal_18847) ) ;
    buf_clk cell_13965 ( .C (clk), .D (signal_18852), .Q (signal_18853) ) ;
    buf_clk cell_13971 ( .C (clk), .D (signal_18858), .Q (signal_18859) ) ;
    buf_clk cell_13977 ( .C (clk), .D (signal_18864), .Q (signal_18865) ) ;
    buf_clk cell_13983 ( .C (clk), .D (signal_18870), .Q (signal_18871) ) ;
    buf_clk cell_13989 ( .C (clk), .D (signal_18876), .Q (signal_18877) ) ;
    buf_clk cell_13995 ( .C (clk), .D (signal_18882), .Q (signal_18883) ) ;
    buf_clk cell_14001 ( .C (clk), .D (signal_18888), .Q (signal_18889) ) ;
    buf_clk cell_14007 ( .C (clk), .D (signal_18894), .Q (signal_18895) ) ;
    buf_clk cell_14013 ( .C (clk), .D (signal_18900), .Q (signal_18901) ) ;
    buf_clk cell_14019 ( .C (clk), .D (signal_18906), .Q (signal_18907) ) ;
    buf_clk cell_14025 ( .C (clk), .D (signal_18912), .Q (signal_18913) ) ;
    buf_clk cell_14031 ( .C (clk), .D (signal_18918), .Q (signal_18919) ) ;
    buf_clk cell_14037 ( .C (clk), .D (signal_18924), .Q (signal_18925) ) ;
    buf_clk cell_14043 ( .C (clk), .D (signal_18930), .Q (signal_18931) ) ;
    buf_clk cell_14049 ( .C (clk), .D (signal_18936), .Q (signal_18937) ) ;
    buf_clk cell_14055 ( .C (clk), .D (signal_18942), .Q (signal_18943) ) ;
    buf_clk cell_14061 ( .C (clk), .D (signal_18948), .Q (signal_18949) ) ;
    buf_clk cell_14067 ( .C (clk), .D (signal_18954), .Q (signal_18955) ) ;
    buf_clk cell_14073 ( .C (clk), .D (signal_18960), .Q (signal_18961) ) ;
    buf_clk cell_14079 ( .C (clk), .D (signal_18966), .Q (signal_18967) ) ;
    buf_clk cell_14085 ( .C (clk), .D (signal_18972), .Q (signal_18973) ) ;
    buf_clk cell_14091 ( .C (clk), .D (signal_18978), .Q (signal_18979) ) ;
    buf_clk cell_14097 ( .C (clk), .D (signal_18984), .Q (signal_18985) ) ;
    buf_clk cell_14103 ( .C (clk), .D (signal_18990), .Q (signal_18991) ) ;
    buf_clk cell_14109 ( .C (clk), .D (signal_18996), .Q (signal_18997) ) ;
    buf_clk cell_14115 ( .C (clk), .D (signal_19002), .Q (signal_19003) ) ;
    buf_clk cell_14121 ( .C (clk), .D (signal_19008), .Q (signal_19009) ) ;
    buf_clk cell_14127 ( .C (clk), .D (signal_19014), .Q (signal_19015) ) ;
    buf_clk cell_14133 ( .C (clk), .D (signal_19020), .Q (signal_19021) ) ;
    buf_clk cell_14139 ( .C (clk), .D (signal_19026), .Q (signal_19027) ) ;
    buf_clk cell_14145 ( .C (clk), .D (signal_19032), .Q (signal_19033) ) ;
    buf_clk cell_14151 ( .C (clk), .D (signal_19038), .Q (signal_19039) ) ;
    buf_clk cell_14157 ( .C (clk), .D (signal_19044), .Q (signal_19045) ) ;
    buf_clk cell_14163 ( .C (clk), .D (signal_19050), .Q (signal_19051) ) ;
    buf_clk cell_14169 ( .C (clk), .D (signal_19056), .Q (signal_19057) ) ;
    buf_clk cell_14175 ( .C (clk), .D (signal_19062), .Q (signal_19063) ) ;
    buf_clk cell_14181 ( .C (clk), .D (signal_19068), .Q (signal_19069) ) ;
    buf_clk cell_14187 ( .C (clk), .D (signal_19074), .Q (signal_19075) ) ;
    buf_clk cell_14193 ( .C (clk), .D (signal_19080), .Q (signal_19081) ) ;
    buf_clk cell_14199 ( .C (clk), .D (signal_19086), .Q (signal_19087) ) ;
    buf_clk cell_14205 ( .C (clk), .D (signal_19092), .Q (signal_19093) ) ;
    buf_clk cell_14211 ( .C (clk), .D (signal_19098), .Q (signal_19099) ) ;
    buf_clk cell_14217 ( .C (clk), .D (signal_19104), .Q (signal_19105) ) ;
    buf_clk cell_14223 ( .C (clk), .D (signal_19110), .Q (signal_19111) ) ;
    buf_clk cell_14229 ( .C (clk), .D (signal_19116), .Q (signal_19117) ) ;
    buf_clk cell_14235 ( .C (clk), .D (signal_19122), .Q (signal_19123) ) ;
    buf_clk cell_14241 ( .C (clk), .D (signal_19128), .Q (signal_19129) ) ;
    buf_clk cell_14247 ( .C (clk), .D (signal_19134), .Q (signal_19135) ) ;
    buf_clk cell_14253 ( .C (clk), .D (signal_19140), .Q (signal_19141) ) ;
    buf_clk cell_14259 ( .C (clk), .D (signal_19146), .Q (signal_19147) ) ;
    buf_clk cell_14265 ( .C (clk), .D (signal_19152), .Q (signal_19153) ) ;
    buf_clk cell_14271 ( .C (clk), .D (signal_19158), .Q (signal_19159) ) ;
    buf_clk cell_14277 ( .C (clk), .D (signal_19164), .Q (signal_19165) ) ;
    buf_clk cell_14283 ( .C (clk), .D (signal_19170), .Q (signal_19171) ) ;
    buf_clk cell_14289 ( .C (clk), .D (signal_19176), .Q (signal_19177) ) ;
    buf_clk cell_14295 ( .C (clk), .D (signal_19182), .Q (signal_19183) ) ;
    buf_clk cell_14301 ( .C (clk), .D (signal_19188), .Q (signal_19189) ) ;
    buf_clk cell_14307 ( .C (clk), .D (signal_19194), .Q (signal_19195) ) ;
    buf_clk cell_14313 ( .C (clk), .D (signal_19200), .Q (signal_19201) ) ;
    buf_clk cell_14319 ( .C (clk), .D (signal_19206), .Q (signal_19207) ) ;
    buf_clk cell_14325 ( .C (clk), .D (signal_19212), .Q (signal_19213) ) ;
    buf_clk cell_14331 ( .C (clk), .D (signal_19218), .Q (signal_19219) ) ;
    buf_clk cell_14337 ( .C (clk), .D (signal_19224), .Q (signal_19225) ) ;
    buf_clk cell_14343 ( .C (clk), .D (signal_19230), .Q (signal_19231) ) ;
    buf_clk cell_14349 ( .C (clk), .D (signal_19236), .Q (signal_19237) ) ;
    buf_clk cell_14355 ( .C (clk), .D (signal_19242), .Q (signal_19243) ) ;
    buf_clk cell_14361 ( .C (clk), .D (signal_19248), .Q (signal_19249) ) ;
    buf_clk cell_14367 ( .C (clk), .D (signal_19254), .Q (signal_19255) ) ;
    buf_clk cell_14373 ( .C (clk), .D (signal_19260), .Q (signal_19261) ) ;
    buf_clk cell_14379 ( .C (clk), .D (signal_19266), .Q (signal_19267) ) ;
    buf_clk cell_14385 ( .C (clk), .D (signal_19272), .Q (signal_19273) ) ;
    buf_clk cell_14391 ( .C (clk), .D (signal_19278), .Q (signal_19279) ) ;
    buf_clk cell_14397 ( .C (clk), .D (signal_19284), .Q (signal_19285) ) ;
    buf_clk cell_14403 ( .C (clk), .D (signal_19290), .Q (signal_19291) ) ;
    buf_clk cell_14409 ( .C (clk), .D (signal_19296), .Q (signal_19297) ) ;
    buf_clk cell_14415 ( .C (clk), .D (signal_19302), .Q (signal_19303) ) ;
    buf_clk cell_14421 ( .C (clk), .D (signal_19308), .Q (signal_19309) ) ;
    buf_clk cell_14427 ( .C (clk), .D (signal_19314), .Q (signal_19315) ) ;
    buf_clk cell_14433 ( .C (clk), .D (signal_19320), .Q (signal_19321) ) ;
    buf_clk cell_14439 ( .C (clk), .D (signal_19326), .Q (signal_19327) ) ;
    buf_clk cell_14445 ( .C (clk), .D (signal_19332), .Q (signal_19333) ) ;
    buf_clk cell_14451 ( .C (clk), .D (signal_19338), .Q (signal_19339) ) ;
    buf_clk cell_14457 ( .C (clk), .D (signal_19344), .Q (signal_19345) ) ;
    buf_clk cell_14463 ( .C (clk), .D (signal_19350), .Q (signal_19351) ) ;
    buf_clk cell_14469 ( .C (clk), .D (signal_19356), .Q (signal_19357) ) ;
    buf_clk cell_14475 ( .C (clk), .D (signal_19362), .Q (signal_19363) ) ;
    buf_clk cell_14481 ( .C (clk), .D (signal_19368), .Q (signal_19369) ) ;
    buf_clk cell_14487 ( .C (clk), .D (signal_19374), .Q (signal_19375) ) ;
    buf_clk cell_14493 ( .C (clk), .D (signal_19380), .Q (signal_19381) ) ;
    buf_clk cell_14499 ( .C (clk), .D (signal_19386), .Q (signal_19387) ) ;
    buf_clk cell_14505 ( .C (clk), .D (signal_19392), .Q (signal_19393) ) ;
    buf_clk cell_14511 ( .C (clk), .D (signal_19398), .Q (signal_19399) ) ;
    buf_clk cell_14517 ( .C (clk), .D (signal_19404), .Q (signal_19405) ) ;
    buf_clk cell_14523 ( .C (clk), .D (signal_19410), .Q (signal_19411) ) ;
    buf_clk cell_14529 ( .C (clk), .D (signal_19416), .Q (signal_19417) ) ;
    buf_clk cell_14535 ( .C (clk), .D (signal_19422), .Q (signal_19423) ) ;
    buf_clk cell_14541 ( .C (clk), .D (signal_19428), .Q (signal_19429) ) ;
    buf_clk cell_14547 ( .C (clk), .D (signal_19434), .Q (signal_19435) ) ;
    buf_clk cell_14553 ( .C (clk), .D (signal_19440), .Q (signal_19441) ) ;
    buf_clk cell_14559 ( .C (clk), .D (signal_19446), .Q (signal_19447) ) ;
    buf_clk cell_14565 ( .C (clk), .D (signal_19452), .Q (signal_19453) ) ;
    buf_clk cell_14571 ( .C (clk), .D (signal_19458), .Q (signal_19459) ) ;
    buf_clk cell_14577 ( .C (clk), .D (signal_19464), .Q (signal_19465) ) ;
    buf_clk cell_14583 ( .C (clk), .D (signal_19470), .Q (signal_19471) ) ;
    buf_clk cell_14589 ( .C (clk), .D (signal_19476), .Q (signal_19477) ) ;
    buf_clk cell_14595 ( .C (clk), .D (signal_19482), .Q (signal_19483) ) ;
    buf_clk cell_14601 ( .C (clk), .D (signal_19488), .Q (signal_19489) ) ;
    buf_clk cell_14607 ( .C (clk), .D (signal_19494), .Q (signal_19495) ) ;
    buf_clk cell_14613 ( .C (clk), .D (signal_19500), .Q (signal_19501) ) ;
    buf_clk cell_14619 ( .C (clk), .D (signal_19506), .Q (signal_19507) ) ;
    buf_clk cell_14625 ( .C (clk), .D (signal_19512), .Q (signal_19513) ) ;
    buf_clk cell_14631 ( .C (clk), .D (signal_19518), .Q (signal_19519) ) ;
    buf_clk cell_14637 ( .C (clk), .D (signal_19524), .Q (signal_19525) ) ;
    buf_clk cell_14643 ( .C (clk), .D (signal_19530), .Q (signal_19531) ) ;
    buf_clk cell_14649 ( .C (clk), .D (signal_19536), .Q (signal_19537) ) ;
    buf_clk cell_14655 ( .C (clk), .D (signal_19542), .Q (signal_19543) ) ;
    buf_clk cell_14661 ( .C (clk), .D (signal_19548), .Q (signal_19549) ) ;
    buf_clk cell_14667 ( .C (clk), .D (signal_19554), .Q (signal_19555) ) ;
    buf_clk cell_14673 ( .C (clk), .D (signal_19560), .Q (signal_19561) ) ;
    buf_clk cell_14679 ( .C (clk), .D (signal_19566), .Q (signal_19567) ) ;
    buf_clk cell_14685 ( .C (clk), .D (signal_19572), .Q (signal_19573) ) ;
    buf_clk cell_14691 ( .C (clk), .D (signal_19578), .Q (signal_19579) ) ;
    buf_clk cell_14697 ( .C (clk), .D (signal_19584), .Q (signal_19585) ) ;
    buf_clk cell_14703 ( .C (clk), .D (signal_19590), .Q (signal_19591) ) ;
    buf_clk cell_14709 ( .C (clk), .D (signal_19596), .Q (signal_19597) ) ;
    buf_clk cell_14715 ( .C (clk), .D (signal_19602), .Q (signal_19603) ) ;
    buf_clk cell_14721 ( .C (clk), .D (signal_19608), .Q (signal_19609) ) ;
    buf_clk cell_14727 ( .C (clk), .D (signal_19614), .Q (signal_19615) ) ;
    buf_clk cell_14733 ( .C (clk), .D (signal_19620), .Q (signal_19621) ) ;
    buf_clk cell_14739 ( .C (clk), .D (signal_19626), .Q (signal_19627) ) ;
    buf_clk cell_14745 ( .C (clk), .D (signal_19632), .Q (signal_19633) ) ;
    buf_clk cell_14751 ( .C (clk), .D (signal_19638), .Q (signal_19639) ) ;
    buf_clk cell_14757 ( .C (clk), .D (signal_19644), .Q (signal_19645) ) ;
    buf_clk cell_14763 ( .C (clk), .D (signal_19650), .Q (signal_19651) ) ;
    buf_clk cell_14769 ( .C (clk), .D (signal_19656), .Q (signal_19657) ) ;
    buf_clk cell_14775 ( .C (clk), .D (signal_19662), .Q (signal_19663) ) ;
    buf_clk cell_14781 ( .C (clk), .D (signal_19668), .Q (signal_19669) ) ;
    buf_clk cell_14787 ( .C (clk), .D (signal_19674), .Q (signal_19675) ) ;
    buf_clk cell_14793 ( .C (clk), .D (signal_19680), .Q (signal_19681) ) ;
    buf_clk cell_14799 ( .C (clk), .D (signal_19686), .Q (signal_19687) ) ;
    buf_clk cell_14805 ( .C (clk), .D (signal_19692), .Q (signal_19693) ) ;
    buf_clk cell_14811 ( .C (clk), .D (signal_19698), .Q (signal_19699) ) ;
    buf_clk cell_14817 ( .C (clk), .D (signal_19704), .Q (signal_19705) ) ;
    buf_clk cell_14823 ( .C (clk), .D (signal_19710), .Q (signal_19711) ) ;
    buf_clk cell_14829 ( .C (clk), .D (signal_19716), .Q (signal_19717) ) ;
    buf_clk cell_14835 ( .C (clk), .D (signal_19722), .Q (signal_19723) ) ;
    buf_clk cell_14841 ( .C (clk), .D (signal_19728), .Q (signal_19729) ) ;
    buf_clk cell_14847 ( .C (clk), .D (signal_19734), .Q (signal_19735) ) ;
    buf_clk cell_14853 ( .C (clk), .D (signal_19740), .Q (signal_19741) ) ;
    buf_clk cell_14859 ( .C (clk), .D (signal_19746), .Q (signal_19747) ) ;
    buf_clk cell_14865 ( .C (clk), .D (signal_19752), .Q (signal_19753) ) ;
    buf_clk cell_14871 ( .C (clk), .D (signal_19758), .Q (signal_19759) ) ;
    buf_clk cell_14877 ( .C (clk), .D (signal_19764), .Q (signal_19765) ) ;
    buf_clk cell_14883 ( .C (clk), .D (signal_19770), .Q (signal_19771) ) ;
    buf_clk cell_14889 ( .C (clk), .D (signal_19776), .Q (signal_19777) ) ;
    buf_clk cell_14895 ( .C (clk), .D (signal_19782), .Q (signal_19783) ) ;
    buf_clk cell_14901 ( .C (clk), .D (signal_19788), .Q (signal_19789) ) ;
    buf_clk cell_14907 ( .C (clk), .D (signal_19794), .Q (signal_19795) ) ;
    buf_clk cell_14913 ( .C (clk), .D (signal_19800), .Q (signal_19801) ) ;
    buf_clk cell_14919 ( .C (clk), .D (signal_19806), .Q (signal_19807) ) ;
    buf_clk cell_14925 ( .C (clk), .D (signal_19812), .Q (signal_19813) ) ;
    buf_clk cell_14931 ( .C (clk), .D (signal_19818), .Q (signal_19819) ) ;
    buf_clk cell_14937 ( .C (clk), .D (signal_19824), .Q (signal_19825) ) ;
    buf_clk cell_14943 ( .C (clk), .D (signal_19830), .Q (signal_19831) ) ;
    buf_clk cell_14949 ( .C (clk), .D (signal_19836), .Q (signal_19837) ) ;
    buf_clk cell_14955 ( .C (clk), .D (signal_19842), .Q (signal_19843) ) ;
    buf_clk cell_14961 ( .C (clk), .D (signal_19848), .Q (signal_19849) ) ;
    buf_clk cell_14967 ( .C (clk), .D (signal_19854), .Q (signal_19855) ) ;
    buf_clk cell_14973 ( .C (clk), .D (signal_19860), .Q (signal_19861) ) ;
    buf_clk cell_14979 ( .C (clk), .D (signal_19866), .Q (signal_19867) ) ;
    buf_clk cell_14985 ( .C (clk), .D (signal_19872), .Q (signal_19873) ) ;
    buf_clk cell_14991 ( .C (clk), .D (signal_19878), .Q (signal_19879) ) ;
    buf_clk cell_14997 ( .C (clk), .D (signal_19884), .Q (signal_19885) ) ;
    buf_clk cell_15003 ( .C (clk), .D (signal_19890), .Q (signal_19891) ) ;
    buf_clk cell_15009 ( .C (clk), .D (signal_19896), .Q (signal_19897) ) ;
    buf_clk cell_15015 ( .C (clk), .D (signal_19902), .Q (signal_19903) ) ;
    buf_clk cell_15021 ( .C (clk), .D (signal_19908), .Q (signal_19909) ) ;
    buf_clk cell_15027 ( .C (clk), .D (signal_19914), .Q (signal_19915) ) ;
    buf_clk cell_15033 ( .C (clk), .D (signal_19920), .Q (signal_19921) ) ;
    buf_clk cell_15039 ( .C (clk), .D (signal_19926), .Q (signal_19927) ) ;
    buf_clk cell_15045 ( .C (clk), .D (signal_19932), .Q (signal_19933) ) ;
    buf_clk cell_15051 ( .C (clk), .D (signal_19938), .Q (signal_19939) ) ;
    buf_clk cell_15057 ( .C (clk), .D (signal_19944), .Q (signal_19945) ) ;
    buf_clk cell_15063 ( .C (clk), .D (signal_19950), .Q (signal_19951) ) ;
    buf_clk cell_15069 ( .C (clk), .D (signal_19956), .Q (signal_19957) ) ;
    buf_clk cell_15075 ( .C (clk), .D (signal_19962), .Q (signal_19963) ) ;
    buf_clk cell_15081 ( .C (clk), .D (signal_19968), .Q (signal_19969) ) ;
    buf_clk cell_15087 ( .C (clk), .D (signal_19974), .Q (signal_19975) ) ;
    buf_clk cell_15093 ( .C (clk), .D (signal_19980), .Q (signal_19981) ) ;
    buf_clk cell_15099 ( .C (clk), .D (signal_19986), .Q (signal_19987) ) ;
    buf_clk cell_15105 ( .C (clk), .D (signal_19992), .Q (signal_19993) ) ;
    buf_clk cell_15111 ( .C (clk), .D (signal_19998), .Q (signal_19999) ) ;
    buf_clk cell_15117 ( .C (clk), .D (signal_20004), .Q (signal_20005) ) ;
    buf_clk cell_15123 ( .C (clk), .D (signal_20010), .Q (signal_20011) ) ;
    buf_clk cell_15129 ( .C (clk), .D (signal_20016), .Q (signal_20017) ) ;
    buf_clk cell_15135 ( .C (clk), .D (signal_20022), .Q (signal_20023) ) ;
    buf_clk cell_15141 ( .C (clk), .D (signal_20028), .Q (signal_20029) ) ;
    buf_clk cell_15147 ( .C (clk), .D (signal_20034), .Q (signal_20035) ) ;
    buf_clk cell_15153 ( .C (clk), .D (signal_20040), .Q (signal_20041) ) ;
    buf_clk cell_15159 ( .C (clk), .D (signal_20046), .Q (signal_20047) ) ;
    buf_clk cell_15165 ( .C (clk), .D (signal_20052), .Q (signal_20053) ) ;
    buf_clk cell_15171 ( .C (clk), .D (signal_20058), .Q (signal_20059) ) ;
    buf_clk cell_15177 ( .C (clk), .D (signal_20064), .Q (signal_20065) ) ;
    buf_clk cell_15183 ( .C (clk), .D (signal_20070), .Q (signal_20071) ) ;
    buf_clk cell_15189 ( .C (clk), .D (signal_20076), .Q (signal_20077) ) ;
    buf_clk cell_15195 ( .C (clk), .D (signal_20082), .Q (signal_20083) ) ;
    buf_clk cell_15201 ( .C (clk), .D (signal_20088), .Q (signal_20089) ) ;
    buf_clk cell_15207 ( .C (clk), .D (signal_20094), .Q (signal_20095) ) ;
    buf_clk cell_15213 ( .C (clk), .D (signal_20100), .Q (signal_20101) ) ;
    buf_clk cell_15219 ( .C (clk), .D (signal_20106), .Q (signal_20107) ) ;
    buf_clk cell_15225 ( .C (clk), .D (signal_20112), .Q (signal_20113) ) ;
    buf_clk cell_15231 ( .C (clk), .D (signal_20118), .Q (signal_20119) ) ;
    buf_clk cell_15237 ( .C (clk), .D (signal_20124), .Q (signal_20125) ) ;
    buf_clk cell_15243 ( .C (clk), .D (signal_20130), .Q (signal_20131) ) ;
    buf_clk cell_15249 ( .C (clk), .D (signal_20136), .Q (signal_20137) ) ;
    buf_clk cell_15255 ( .C (clk), .D (signal_20142), .Q (signal_20143) ) ;
    buf_clk cell_15261 ( .C (clk), .D (signal_20148), .Q (signal_20149) ) ;
    buf_clk cell_15267 ( .C (clk), .D (signal_20154), .Q (signal_20155) ) ;
    buf_clk cell_15273 ( .C (clk), .D (signal_20160), .Q (signal_20161) ) ;
    buf_clk cell_15279 ( .C (clk), .D (signal_20166), .Q (signal_20167) ) ;
    buf_clk cell_15285 ( .C (clk), .D (signal_20172), .Q (signal_20173) ) ;
    buf_clk cell_15291 ( .C (clk), .D (signal_20178), .Q (signal_20179) ) ;
    buf_clk cell_15297 ( .C (clk), .D (signal_20184), .Q (signal_20185) ) ;
    buf_clk cell_15303 ( .C (clk), .D (signal_20190), .Q (signal_20191) ) ;
    buf_clk cell_15309 ( .C (clk), .D (signal_20196), .Q (signal_20197) ) ;
    buf_clk cell_15315 ( .C (clk), .D (signal_20202), .Q (signal_20203) ) ;
    buf_clk cell_15321 ( .C (clk), .D (signal_20208), .Q (signal_20209) ) ;
    buf_clk cell_15327 ( .C (clk), .D (signal_20214), .Q (signal_20215) ) ;
    buf_clk cell_15333 ( .C (clk), .D (signal_20220), .Q (signal_20221) ) ;
    buf_clk cell_15339 ( .C (clk), .D (signal_20226), .Q (signal_20227) ) ;
    buf_clk cell_15345 ( .C (clk), .D (signal_20232), .Q (signal_20233) ) ;
    buf_clk cell_15351 ( .C (clk), .D (signal_20238), .Q (signal_20239) ) ;
    buf_clk cell_15357 ( .C (clk), .D (signal_20244), .Q (signal_20245) ) ;
    buf_clk cell_15363 ( .C (clk), .D (signal_20250), .Q (signal_20251) ) ;
    buf_clk cell_15369 ( .C (clk), .D (signal_20256), .Q (signal_20257) ) ;
    buf_clk cell_15375 ( .C (clk), .D (signal_20262), .Q (signal_20263) ) ;
    buf_clk cell_15381 ( .C (clk), .D (signal_20268), .Q (signal_20269) ) ;
    buf_clk cell_15387 ( .C (clk), .D (signal_20274), .Q (signal_20275) ) ;
    buf_clk cell_15393 ( .C (clk), .D (signal_20280), .Q (signal_20281) ) ;
    buf_clk cell_15399 ( .C (clk), .D (signal_20286), .Q (signal_20287) ) ;
    buf_clk cell_15405 ( .C (clk), .D (signal_20292), .Q (signal_20293) ) ;
    buf_clk cell_15411 ( .C (clk), .D (signal_20298), .Q (signal_20299) ) ;
    buf_clk cell_15417 ( .C (clk), .D (signal_20304), .Q (signal_20305) ) ;
    buf_clk cell_15423 ( .C (clk), .D (signal_20310), .Q (signal_20311) ) ;
    buf_clk cell_15429 ( .C (clk), .D (signal_20316), .Q (signal_20317) ) ;
    buf_clk cell_15435 ( .C (clk), .D (signal_20322), .Q (signal_20323) ) ;
    buf_clk cell_15441 ( .C (clk), .D (signal_20328), .Q (signal_20329) ) ;
    buf_clk cell_15447 ( .C (clk), .D (signal_20334), .Q (signal_20335) ) ;
    buf_clk cell_15453 ( .C (clk), .D (signal_20340), .Q (signal_20341) ) ;
    buf_clk cell_15459 ( .C (clk), .D (signal_20346), .Q (signal_20347) ) ;
    buf_clk cell_15465 ( .C (clk), .D (signal_20352), .Q (signal_20353) ) ;
    buf_clk cell_15471 ( .C (clk), .D (signal_20358), .Q (signal_20359) ) ;
    buf_clk cell_15477 ( .C (clk), .D (signal_20364), .Q (signal_20365) ) ;
    buf_clk cell_15483 ( .C (clk), .D (signal_20370), .Q (signal_20371) ) ;
    buf_clk cell_15489 ( .C (clk), .D (signal_20376), .Q (signal_20377) ) ;
    buf_clk cell_15495 ( .C (clk), .D (signal_20382), .Q (signal_20383) ) ;
    buf_clk cell_15501 ( .C (clk), .D (signal_20388), .Q (signal_20389) ) ;
    buf_clk cell_15507 ( .C (clk), .D (signal_20394), .Q (signal_20395) ) ;
    buf_clk cell_15513 ( .C (clk), .D (signal_20400), .Q (signal_20401) ) ;
    buf_clk cell_15519 ( .C (clk), .D (signal_20406), .Q (signal_20407) ) ;
    buf_clk cell_15525 ( .C (clk), .D (signal_20412), .Q (signal_20413) ) ;
    buf_clk cell_15531 ( .C (clk), .D (signal_20418), .Q (signal_20419) ) ;
    buf_clk cell_15537 ( .C (clk), .D (signal_20424), .Q (signal_20425) ) ;
    buf_clk cell_15543 ( .C (clk), .D (signal_20430), .Q (signal_20431) ) ;
    buf_clk cell_15549 ( .C (clk), .D (signal_20436), .Q (signal_20437) ) ;
    buf_clk cell_15555 ( .C (clk), .D (signal_20442), .Q (signal_20443) ) ;
    buf_clk cell_15561 ( .C (clk), .D (signal_20448), .Q (signal_20449) ) ;
    buf_clk cell_15567 ( .C (clk), .D (signal_20454), .Q (signal_20455) ) ;
    buf_clk cell_15573 ( .C (clk), .D (signal_20460), .Q (signal_20461) ) ;
    buf_clk cell_15579 ( .C (clk), .D (signal_20466), .Q (signal_20467) ) ;
    buf_clk cell_15585 ( .C (clk), .D (signal_20472), .Q (signal_20473) ) ;
    buf_clk cell_15591 ( .C (clk), .D (signal_20478), .Q (signal_20479) ) ;
    buf_clk cell_15597 ( .C (clk), .D (signal_20484), .Q (signal_20485) ) ;
    buf_clk cell_15603 ( .C (clk), .D (signal_20490), .Q (signal_20491) ) ;
    buf_clk cell_15609 ( .C (clk), .D (signal_20496), .Q (signal_20497) ) ;
    buf_clk cell_15615 ( .C (clk), .D (signal_20502), .Q (signal_20503) ) ;
    buf_clk cell_15621 ( .C (clk), .D (signal_20508), .Q (signal_20509) ) ;
    buf_clk cell_15627 ( .C (clk), .D (signal_20514), .Q (signal_20515) ) ;
    buf_clk cell_15633 ( .C (clk), .D (signal_20520), .Q (signal_20521) ) ;
    buf_clk cell_15639 ( .C (clk), .D (signal_20526), .Q (signal_20527) ) ;
    buf_clk cell_15645 ( .C (clk), .D (signal_20532), .Q (signal_20533) ) ;
    buf_clk cell_15651 ( .C (clk), .D (signal_20538), .Q (signal_20539) ) ;
    buf_clk cell_15657 ( .C (clk), .D (signal_20544), .Q (signal_20545) ) ;
    buf_clk cell_15663 ( .C (clk), .D (signal_20550), .Q (signal_20551) ) ;
    buf_clk cell_15669 ( .C (clk), .D (signal_20556), .Q (signal_20557) ) ;
    buf_clk cell_15675 ( .C (clk), .D (signal_20562), .Q (signal_20563) ) ;
    buf_clk cell_15681 ( .C (clk), .D (signal_20568), .Q (signal_20569) ) ;
    buf_clk cell_15687 ( .C (clk), .D (signal_20574), .Q (signal_20575) ) ;
    buf_clk cell_15693 ( .C (clk), .D (signal_20580), .Q (signal_20581) ) ;
    buf_clk cell_15699 ( .C (clk), .D (signal_20586), .Q (signal_20587) ) ;
    buf_clk cell_15705 ( .C (clk), .D (signal_20592), .Q (signal_20593) ) ;
    buf_clk cell_15711 ( .C (clk), .D (signal_20598), .Q (signal_20599) ) ;
    buf_clk cell_15717 ( .C (clk), .D (signal_20604), .Q (signal_20605) ) ;
    buf_clk cell_15723 ( .C (clk), .D (signal_20610), .Q (signal_20611) ) ;
    buf_clk cell_15729 ( .C (clk), .D (signal_20616), .Q (signal_20617) ) ;
    buf_clk cell_15735 ( .C (clk), .D (signal_20622), .Q (signal_20623) ) ;
    buf_clk cell_15741 ( .C (clk), .D (signal_20628), .Q (signal_20629) ) ;
    buf_clk cell_15747 ( .C (clk), .D (signal_20634), .Q (signal_20635) ) ;
    buf_clk cell_15753 ( .C (clk), .D (signal_20640), .Q (signal_20641) ) ;
    buf_clk cell_15759 ( .C (clk), .D (signal_20646), .Q (signal_20647) ) ;
    buf_clk cell_15765 ( .C (clk), .D (signal_20652), .Q (signal_20653) ) ;
    buf_clk cell_15771 ( .C (clk), .D (signal_20658), .Q (signal_20659) ) ;
    buf_clk cell_15777 ( .C (clk), .D (signal_20664), .Q (signal_20665) ) ;
    buf_clk cell_15783 ( .C (clk), .D (signal_20670), .Q (signal_20671) ) ;
    buf_clk cell_15789 ( .C (clk), .D (signal_20676), .Q (signal_20677) ) ;
    buf_clk cell_15795 ( .C (clk), .D (signal_20682), .Q (signal_20683) ) ;
    buf_clk cell_15801 ( .C (clk), .D (signal_20688), .Q (signal_20689) ) ;
    buf_clk cell_15807 ( .C (clk), .D (signal_20694), .Q (signal_20695) ) ;
    buf_clk cell_15813 ( .C (clk), .D (signal_20700), .Q (signal_20701) ) ;
    buf_clk cell_15819 ( .C (clk), .D (signal_20706), .Q (signal_20707) ) ;
    buf_clk cell_15825 ( .C (clk), .D (signal_20712), .Q (signal_20713) ) ;
    buf_clk cell_15831 ( .C (clk), .D (signal_20718), .Q (signal_20719) ) ;
    buf_clk cell_15837 ( .C (clk), .D (signal_20724), .Q (signal_20725) ) ;
    buf_clk cell_15843 ( .C (clk), .D (signal_20730), .Q (signal_20731) ) ;
    buf_clk cell_15849 ( .C (clk), .D (signal_20736), .Q (signal_20737) ) ;
    buf_clk cell_15855 ( .C (clk), .D (signal_20742), .Q (signal_20743) ) ;
    buf_clk cell_15861 ( .C (clk), .D (signal_20748), .Q (signal_20749) ) ;
    buf_clk cell_15867 ( .C (clk), .D (signal_20754), .Q (signal_20755) ) ;
    buf_clk cell_15873 ( .C (clk), .D (signal_20760), .Q (signal_20761) ) ;
    buf_clk cell_15879 ( .C (clk), .D (signal_20766), .Q (signal_20767) ) ;
    buf_clk cell_15885 ( .C (clk), .D (signal_20772), .Q (signal_20773) ) ;
    buf_clk cell_15891 ( .C (clk), .D (signal_20778), .Q (signal_20779) ) ;
    buf_clk cell_15897 ( .C (clk), .D (signal_20784), .Q (signal_20785) ) ;
    buf_clk cell_15903 ( .C (clk), .D (signal_20790), .Q (signal_20791) ) ;
    buf_clk cell_15909 ( .C (clk), .D (signal_20796), .Q (signal_20797) ) ;
    buf_clk cell_15915 ( .C (clk), .D (signal_20802), .Q (signal_20803) ) ;
    buf_clk cell_15921 ( .C (clk), .D (signal_20808), .Q (signal_20809) ) ;
    buf_clk cell_15927 ( .C (clk), .D (signal_20814), .Q (signal_20815) ) ;
    buf_clk cell_15933 ( .C (clk), .D (signal_20820), .Q (signal_20821) ) ;
    buf_clk cell_15939 ( .C (clk), .D (signal_20826), .Q (signal_20827) ) ;
    buf_clk cell_15945 ( .C (clk), .D (signal_20832), .Q (signal_20833) ) ;
    buf_clk cell_15951 ( .C (clk), .D (signal_20838), .Q (signal_20839) ) ;
    buf_clk cell_15957 ( .C (clk), .D (signal_20844), .Q (signal_20845) ) ;
    buf_clk cell_15963 ( .C (clk), .D (signal_20850), .Q (signal_20851) ) ;
    buf_clk cell_15969 ( .C (clk), .D (signal_20856), .Q (signal_20857) ) ;
    buf_clk cell_15975 ( .C (clk), .D (signal_20862), .Q (signal_20863) ) ;
    buf_clk cell_15981 ( .C (clk), .D (signal_20868), .Q (signal_20869) ) ;
    buf_clk cell_15987 ( .C (clk), .D (signal_20874), .Q (signal_20875) ) ;
    buf_clk cell_15993 ( .C (clk), .D (signal_20880), .Q (signal_20881) ) ;
    buf_clk cell_15999 ( .C (clk), .D (signal_20886), .Q (signal_20887) ) ;
    buf_clk cell_16005 ( .C (clk), .D (signal_20892), .Q (signal_20893) ) ;
    buf_clk cell_16011 ( .C (clk), .D (signal_20898), .Q (signal_20899) ) ;
    buf_clk cell_16017 ( .C (clk), .D (signal_20904), .Q (signal_20905) ) ;
    buf_clk cell_16023 ( .C (clk), .D (signal_20910), .Q (signal_20911) ) ;
    buf_clk cell_16029 ( .C (clk), .D (signal_20916), .Q (signal_20917) ) ;
    buf_clk cell_16035 ( .C (clk), .D (signal_20922), .Q (signal_20923) ) ;
    buf_clk cell_16041 ( .C (clk), .D (signal_20928), .Q (signal_20929) ) ;
    buf_clk cell_16047 ( .C (clk), .D (signal_20934), .Q (signal_20935) ) ;
    buf_clk cell_16053 ( .C (clk), .D (signal_20940), .Q (signal_20941) ) ;
    buf_clk cell_16059 ( .C (clk), .D (signal_20946), .Q (signal_20947) ) ;
    buf_clk cell_16065 ( .C (clk), .D (signal_20952), .Q (signal_20953) ) ;
    buf_clk cell_16071 ( .C (clk), .D (signal_20958), .Q (signal_20959) ) ;
    buf_clk cell_16077 ( .C (clk), .D (signal_20964), .Q (signal_20965) ) ;
    buf_clk cell_16083 ( .C (clk), .D (signal_20970), .Q (signal_20971) ) ;
    buf_clk cell_16089 ( .C (clk), .D (signal_20976), .Q (signal_20977) ) ;
    buf_clk cell_16095 ( .C (clk), .D (signal_20982), .Q (signal_20983) ) ;
    buf_clk cell_16101 ( .C (clk), .D (signal_20988), .Q (signal_20989) ) ;
    buf_clk cell_16107 ( .C (clk), .D (signal_20994), .Q (signal_20995) ) ;
    buf_clk cell_16113 ( .C (clk), .D (signal_21000), .Q (signal_21001) ) ;
    buf_clk cell_16119 ( .C (clk), .D (signal_21006), .Q (signal_21007) ) ;
    buf_clk cell_16125 ( .C (clk), .D (signal_21012), .Q (signal_21013) ) ;
    buf_clk cell_16131 ( .C (clk), .D (signal_21018), .Q (signal_21019) ) ;
    buf_clk cell_16137 ( .C (clk), .D (signal_21024), .Q (signal_21025) ) ;
    buf_clk cell_16143 ( .C (clk), .D (signal_21030), .Q (signal_21031) ) ;
    buf_clk cell_16149 ( .C (clk), .D (signal_21036), .Q (signal_21037) ) ;
    buf_clk cell_16155 ( .C (clk), .D (signal_21042), .Q (signal_21043) ) ;
    buf_clk cell_16161 ( .C (clk), .D (signal_21048), .Q (signal_21049) ) ;
    buf_clk cell_16167 ( .C (clk), .D (signal_21054), .Q (signal_21055) ) ;
    buf_clk cell_16173 ( .C (clk), .D (signal_21060), .Q (signal_21061) ) ;
    buf_clk cell_16179 ( .C (clk), .D (signal_21066), .Q (signal_21067) ) ;
    buf_clk cell_16185 ( .C (clk), .D (signal_21072), .Q (signal_21073) ) ;
    buf_clk cell_16191 ( .C (clk), .D (signal_21078), .Q (signal_21079) ) ;
    buf_clk cell_16197 ( .C (clk), .D (signal_21084), .Q (signal_21085) ) ;
    buf_clk cell_16203 ( .C (clk), .D (signal_21090), .Q (signal_21091) ) ;
    buf_clk cell_16209 ( .C (clk), .D (signal_21096), .Q (signal_21097) ) ;
    buf_clk cell_16215 ( .C (clk), .D (signal_21102), .Q (signal_21103) ) ;
    buf_clk cell_16221 ( .C (clk), .D (signal_21108), .Q (signal_21109) ) ;
    buf_clk cell_16227 ( .C (clk), .D (signal_21114), .Q (signal_21115) ) ;
    buf_clk cell_16233 ( .C (clk), .D (signal_21120), .Q (signal_21121) ) ;
    buf_clk cell_16239 ( .C (clk), .D (signal_21126), .Q (signal_21127) ) ;
    buf_clk cell_16245 ( .C (clk), .D (signal_21132), .Q (signal_21133) ) ;
    buf_clk cell_16251 ( .C (clk), .D (signal_21138), .Q (signal_21139) ) ;
    buf_clk cell_16257 ( .C (clk), .D (signal_21144), .Q (signal_21145) ) ;
    buf_clk cell_16263 ( .C (clk), .D (signal_21150), .Q (signal_21151) ) ;
    buf_clk cell_16269 ( .C (clk), .D (signal_21156), .Q (signal_21157) ) ;
    buf_clk cell_16275 ( .C (clk), .D (signal_21162), .Q (signal_21163) ) ;
    buf_clk cell_16281 ( .C (clk), .D (signal_21168), .Q (signal_21169) ) ;
    buf_clk cell_16287 ( .C (clk), .D (signal_21174), .Q (signal_21175) ) ;
    buf_clk cell_16293 ( .C (clk), .D (signal_21180), .Q (signal_21181) ) ;
    buf_clk cell_16299 ( .C (clk), .D (signal_21186), .Q (signal_21187) ) ;
    buf_clk cell_16305 ( .C (clk), .D (signal_21192), .Q (signal_21193) ) ;
    buf_clk cell_16311 ( .C (clk), .D (signal_21198), .Q (signal_21199) ) ;
    buf_clk cell_16317 ( .C (clk), .D (signal_21204), .Q (signal_21205) ) ;
    buf_clk cell_16323 ( .C (clk), .D (signal_21210), .Q (signal_21211) ) ;
    buf_clk cell_16329 ( .C (clk), .D (signal_21216), .Q (signal_21217) ) ;
    buf_clk cell_16335 ( .C (clk), .D (signal_21222), .Q (signal_21223) ) ;
    buf_clk cell_16341 ( .C (clk), .D (signal_21228), .Q (signal_21229) ) ;
    buf_clk cell_16347 ( .C (clk), .D (signal_21234), .Q (signal_21235) ) ;
    buf_clk cell_16353 ( .C (clk), .D (signal_21240), .Q (signal_21241) ) ;
    buf_clk cell_16359 ( .C (clk), .D (signal_21246), .Q (signal_21247) ) ;
    buf_clk cell_16365 ( .C (clk), .D (signal_21252), .Q (signal_21253) ) ;
    buf_clk cell_16371 ( .C (clk), .D (signal_21258), .Q (signal_21259) ) ;
    buf_clk cell_16377 ( .C (clk), .D (signal_21264), .Q (signal_21265) ) ;
    buf_clk cell_16383 ( .C (clk), .D (signal_21270), .Q (signal_21271) ) ;
    buf_clk cell_16389 ( .C (clk), .D (signal_21276), .Q (signal_21277) ) ;
    buf_clk cell_16395 ( .C (clk), .D (signal_21282), .Q (signal_21283) ) ;
    buf_clk cell_16401 ( .C (clk), .D (signal_21288), .Q (signal_21289) ) ;
    buf_clk cell_16407 ( .C (clk), .D (signal_21294), .Q (signal_21295) ) ;
    buf_clk cell_16413 ( .C (clk), .D (signal_21300), .Q (signal_21301) ) ;
    buf_clk cell_16419 ( .C (clk), .D (signal_21306), .Q (signal_21307) ) ;
    buf_clk cell_16425 ( .C (clk), .D (signal_21312), .Q (signal_21313) ) ;
    buf_clk cell_16431 ( .C (clk), .D (signal_21318), .Q (signal_21319) ) ;
    buf_clk cell_16437 ( .C (clk), .D (signal_21324), .Q (signal_21325) ) ;
    buf_clk cell_16443 ( .C (clk), .D (signal_21330), .Q (signal_21331) ) ;
    buf_clk cell_16449 ( .C (clk), .D (signal_21336), .Q (signal_21337) ) ;
    buf_clk cell_16455 ( .C (clk), .D (signal_21342), .Q (signal_21343) ) ;
    buf_clk cell_16461 ( .C (clk), .D (signal_21348), .Q (signal_21349) ) ;
    buf_clk cell_16467 ( .C (clk), .D (signal_21354), .Q (signal_21355) ) ;
    buf_clk cell_16473 ( .C (clk), .D (signal_21360), .Q (signal_21361) ) ;
    buf_clk cell_16479 ( .C (clk), .D (signal_21366), .Q (signal_21367) ) ;
    buf_clk cell_16485 ( .C (clk), .D (signal_21372), .Q (signal_21373) ) ;
    buf_clk cell_16491 ( .C (clk), .D (signal_21378), .Q (signal_21379) ) ;
    buf_clk cell_16497 ( .C (clk), .D (signal_21384), .Q (signal_21385) ) ;
    buf_clk cell_16503 ( .C (clk), .D (signal_21390), .Q (signal_21391) ) ;
    buf_clk cell_16509 ( .C (clk), .D (signal_21396), .Q (signal_21397) ) ;
    buf_clk cell_16515 ( .C (clk), .D (signal_21402), .Q (signal_21403) ) ;
    buf_clk cell_16521 ( .C (clk), .D (signal_21408), .Q (signal_21409) ) ;
    buf_clk cell_16527 ( .C (clk), .D (signal_21414), .Q (signal_21415) ) ;
    buf_clk cell_16533 ( .C (clk), .D (signal_21420), .Q (signal_21421) ) ;
    buf_clk cell_16539 ( .C (clk), .D (signal_21426), .Q (signal_21427) ) ;
    buf_clk cell_16545 ( .C (clk), .D (signal_21432), .Q (signal_21433) ) ;
    buf_clk cell_16551 ( .C (clk), .D (signal_21438), .Q (signal_21439) ) ;
    buf_clk cell_16557 ( .C (clk), .D (signal_21444), .Q (signal_21445) ) ;
    buf_clk cell_16563 ( .C (clk), .D (signal_21450), .Q (signal_21451) ) ;
    buf_clk cell_16569 ( .C (clk), .D (signal_21456), .Q (signal_21457) ) ;
    buf_clk cell_16575 ( .C (clk), .D (signal_21462), .Q (signal_21463) ) ;
    buf_clk cell_16581 ( .C (clk), .D (signal_21468), .Q (signal_21469) ) ;
    buf_clk cell_16587 ( .C (clk), .D (signal_21474), .Q (signal_21475) ) ;
    buf_clk cell_16593 ( .C (clk), .D (signal_21480), .Q (signal_21481) ) ;
    buf_clk cell_16599 ( .C (clk), .D (signal_21486), .Q (signal_21487) ) ;
    buf_clk cell_16605 ( .C (clk), .D (signal_21492), .Q (signal_21493) ) ;
    buf_clk cell_16611 ( .C (clk), .D (signal_21498), .Q (signal_21499) ) ;
    buf_clk cell_16617 ( .C (clk), .D (signal_21504), .Q (signal_21505) ) ;
    buf_clk cell_16623 ( .C (clk), .D (signal_21510), .Q (signal_21511) ) ;
    buf_clk cell_16629 ( .C (clk), .D (signal_21516), .Q (signal_21517) ) ;
    buf_clk cell_16635 ( .C (clk), .D (signal_21522), .Q (signal_21523) ) ;
    buf_clk cell_16641 ( .C (clk), .D (signal_21528), .Q (signal_21529) ) ;
    buf_clk cell_16647 ( .C (clk), .D (signal_21534), .Q (signal_21535) ) ;
    buf_clk cell_16653 ( .C (clk), .D (signal_21540), .Q (signal_21541) ) ;
    buf_clk cell_16659 ( .C (clk), .D (signal_21546), .Q (signal_21547) ) ;
    buf_clk cell_16665 ( .C (clk), .D (signal_21552), .Q (signal_21553) ) ;
    buf_clk cell_16671 ( .C (clk), .D (signal_21558), .Q (signal_21559) ) ;
    buf_clk cell_16677 ( .C (clk), .D (signal_21564), .Q (signal_21565) ) ;
    buf_clk cell_16683 ( .C (clk), .D (signal_21570), .Q (signal_21571) ) ;
    buf_clk cell_16689 ( .C (clk), .D (signal_21576), .Q (signal_21577) ) ;
    buf_clk cell_16695 ( .C (clk), .D (signal_21582), .Q (signal_21583) ) ;
    buf_clk cell_16701 ( .C (clk), .D (signal_21588), .Q (signal_21589) ) ;
    buf_clk cell_16707 ( .C (clk), .D (signal_21594), .Q (signal_21595) ) ;
    buf_clk cell_16713 ( .C (clk), .D (signal_21600), .Q (signal_21601) ) ;
    buf_clk cell_16719 ( .C (clk), .D (signal_21606), .Q (signal_21607) ) ;
    buf_clk cell_16725 ( .C (clk), .D (signal_21612), .Q (signal_21613) ) ;
    buf_clk cell_16731 ( .C (clk), .D (signal_21618), .Q (signal_21619) ) ;
    buf_clk cell_16737 ( .C (clk), .D (signal_21624), .Q (signal_21625) ) ;
    buf_clk cell_16743 ( .C (clk), .D (signal_21630), .Q (signal_21631) ) ;
    buf_clk cell_16749 ( .C (clk), .D (signal_21636), .Q (signal_21637) ) ;
    buf_clk cell_16755 ( .C (clk), .D (signal_21642), .Q (signal_21643) ) ;
    buf_clk cell_16761 ( .C (clk), .D (signal_21648), .Q (signal_21649) ) ;
    buf_clk cell_16767 ( .C (clk), .D (signal_21654), .Q (signal_21655) ) ;
    buf_clk cell_16773 ( .C (clk), .D (signal_21660), .Q (signal_21661) ) ;
    buf_clk cell_16779 ( .C (clk), .D (signal_21666), .Q (signal_21667) ) ;
    buf_clk cell_16785 ( .C (clk), .D (signal_21672), .Q (signal_21673) ) ;
    buf_clk cell_16791 ( .C (clk), .D (signal_21678), .Q (signal_21679) ) ;
    buf_clk cell_16797 ( .C (clk), .D (signal_21684), .Q (signal_21685) ) ;
    buf_clk cell_16803 ( .C (clk), .D (signal_21690), .Q (signal_21691) ) ;
    buf_clk cell_16809 ( .C (clk), .D (signal_21696), .Q (signal_21697) ) ;
    buf_clk cell_16815 ( .C (clk), .D (signal_21702), .Q (signal_21703) ) ;
    buf_clk cell_16821 ( .C (clk), .D (signal_21708), .Q (signal_21709) ) ;
    buf_clk cell_16827 ( .C (clk), .D (signal_21714), .Q (signal_21715) ) ;
    buf_clk cell_16833 ( .C (clk), .D (signal_21720), .Q (signal_21721) ) ;
    buf_clk cell_16839 ( .C (clk), .D (signal_21726), .Q (signal_21727) ) ;
    buf_clk cell_16845 ( .C (clk), .D (signal_21732), .Q (signal_21733) ) ;
    buf_clk cell_16851 ( .C (clk), .D (signal_21738), .Q (signal_21739) ) ;
    buf_clk cell_16857 ( .C (clk), .D (signal_21744), .Q (signal_21745) ) ;
    buf_clk cell_16863 ( .C (clk), .D (signal_21750), .Q (signal_21751) ) ;
    buf_clk cell_16869 ( .C (clk), .D (signal_21756), .Q (signal_21757) ) ;
    buf_clk cell_16875 ( .C (clk), .D (signal_21762), .Q (signal_21763) ) ;
    buf_clk cell_16881 ( .C (clk), .D (signal_21768), .Q (signal_21769) ) ;
    buf_clk cell_16887 ( .C (clk), .D (signal_21774), .Q (signal_21775) ) ;
    buf_clk cell_16893 ( .C (clk), .D (signal_21780), .Q (signal_21781) ) ;
    buf_clk cell_16899 ( .C (clk), .D (signal_21786), .Q (signal_21787) ) ;
    buf_clk cell_16905 ( .C (clk), .D (signal_21792), .Q (signal_21793) ) ;
    buf_clk cell_16911 ( .C (clk), .D (signal_21798), .Q (signal_21799) ) ;
    buf_clk cell_16917 ( .C (clk), .D (signal_21804), .Q (signal_21805) ) ;
    buf_clk cell_16923 ( .C (clk), .D (signal_21810), .Q (signal_21811) ) ;
    buf_clk cell_16929 ( .C (clk), .D (signal_21816), .Q (signal_21817) ) ;
    buf_clk cell_16935 ( .C (clk), .D (signal_21822), .Q (signal_21823) ) ;
    buf_clk cell_16941 ( .C (clk), .D (signal_21828), .Q (signal_21829) ) ;
    buf_clk cell_16947 ( .C (clk), .D (signal_21834), .Q (signal_21835) ) ;
    buf_clk cell_16953 ( .C (clk), .D (signal_21840), .Q (signal_21841) ) ;
    buf_clk cell_16959 ( .C (clk), .D (signal_21846), .Q (signal_21847) ) ;
    buf_clk cell_16965 ( .C (clk), .D (signal_21852), .Q (signal_21853) ) ;
    buf_clk cell_16971 ( .C (clk), .D (signal_21858), .Q (signal_21859) ) ;
    buf_clk cell_16977 ( .C (clk), .D (signal_21864), .Q (signal_21865) ) ;
    buf_clk cell_16983 ( .C (clk), .D (signal_21870), .Q (signal_21871) ) ;
    buf_clk cell_16989 ( .C (clk), .D (signal_21876), .Q (signal_21877) ) ;
    buf_clk cell_16995 ( .C (clk), .D (signal_21882), .Q (signal_21883) ) ;
    buf_clk cell_17001 ( .C (clk), .D (signal_21888), .Q (signal_21889) ) ;
    buf_clk cell_17007 ( .C (clk), .D (signal_21894), .Q (signal_21895) ) ;
    buf_clk cell_17013 ( .C (clk), .D (signal_21900), .Q (signal_21901) ) ;
    buf_clk cell_17019 ( .C (clk), .D (signal_21906), .Q (signal_21907) ) ;
    buf_clk cell_17025 ( .C (clk), .D (signal_21912), .Q (signal_21913) ) ;
    buf_clk cell_17031 ( .C (clk), .D (signal_21918), .Q (signal_21919) ) ;
    buf_clk cell_17037 ( .C (clk), .D (signal_21924), .Q (signal_21925) ) ;
    buf_clk cell_17043 ( .C (clk), .D (signal_21930), .Q (signal_21931) ) ;
    buf_clk cell_17049 ( .C (clk), .D (signal_21936), .Q (signal_21937) ) ;
    buf_clk cell_17055 ( .C (clk), .D (signal_21942), .Q (signal_21943) ) ;
    buf_clk cell_17061 ( .C (clk), .D (signal_21948), .Q (signal_21949) ) ;
    buf_clk cell_17067 ( .C (clk), .D (signal_21954), .Q (signal_21955) ) ;
    buf_clk cell_17073 ( .C (clk), .D (signal_21960), .Q (signal_21961) ) ;
    buf_clk cell_17079 ( .C (clk), .D (signal_21966), .Q (signal_21967) ) ;
    buf_clk cell_17085 ( .C (clk), .D (signal_21972), .Q (signal_21973) ) ;
    buf_clk cell_17091 ( .C (clk), .D (signal_21978), .Q (signal_21979) ) ;
    buf_clk cell_17097 ( .C (clk), .D (signal_21984), .Q (signal_21985) ) ;
    buf_clk cell_17103 ( .C (clk), .D (signal_21990), .Q (signal_21991) ) ;
    buf_clk cell_17109 ( .C (clk), .D (signal_21996), .Q (signal_21997) ) ;
    buf_clk cell_17115 ( .C (clk), .D (signal_22002), .Q (signal_22003) ) ;
    buf_clk cell_17121 ( .C (clk), .D (signal_22008), .Q (signal_22009) ) ;
    buf_clk cell_17127 ( .C (clk), .D (signal_22014), .Q (signal_22015) ) ;
    buf_clk cell_17133 ( .C (clk), .D (signal_22020), .Q (signal_22021) ) ;
    buf_clk cell_17139 ( .C (clk), .D (signal_22026), .Q (signal_22027) ) ;
    buf_clk cell_17145 ( .C (clk), .D (signal_22032), .Q (signal_22033) ) ;
    buf_clk cell_17151 ( .C (clk), .D (signal_22038), .Q (signal_22039) ) ;
    buf_clk cell_17157 ( .C (clk), .D (signal_22044), .Q (signal_22045) ) ;
    buf_clk cell_17163 ( .C (clk), .D (signal_22050), .Q (signal_22051) ) ;
    buf_clk cell_17169 ( .C (clk), .D (signal_22056), .Q (signal_22057) ) ;
    buf_clk cell_17175 ( .C (clk), .D (signal_22062), .Q (signal_22063) ) ;
    buf_clk cell_17181 ( .C (clk), .D (signal_22068), .Q (signal_22069) ) ;
    buf_clk cell_17187 ( .C (clk), .D (signal_22074), .Q (signal_22075) ) ;
    buf_clk cell_17193 ( .C (clk), .D (signal_22080), .Q (signal_22081) ) ;
    buf_clk cell_17199 ( .C (clk), .D (signal_22086), .Q (signal_22087) ) ;
    buf_clk cell_17205 ( .C (clk), .D (signal_22092), .Q (signal_22093) ) ;
    buf_clk cell_17211 ( .C (clk), .D (signal_22098), .Q (signal_22099) ) ;
    buf_clk cell_17217 ( .C (clk), .D (signal_22104), .Q (signal_22105) ) ;
    buf_clk cell_17223 ( .C (clk), .D (signal_22110), .Q (signal_22111) ) ;
    buf_clk cell_17229 ( .C (clk), .D (signal_22116), .Q (signal_22117) ) ;
    buf_clk cell_17235 ( .C (clk), .D (signal_22122), .Q (signal_22123) ) ;
    buf_clk cell_17241 ( .C (clk), .D (signal_22128), .Q (signal_22129) ) ;
    buf_clk cell_17247 ( .C (clk), .D (signal_22134), .Q (signal_22135) ) ;
    buf_clk cell_17253 ( .C (clk), .D (signal_22140), .Q (signal_22141) ) ;
    buf_clk cell_17259 ( .C (clk), .D (signal_22146), .Q (signal_22147) ) ;
    buf_clk cell_17265 ( .C (clk), .D (signal_22152), .Q (signal_22153) ) ;
    buf_clk cell_17271 ( .C (clk), .D (signal_22158), .Q (signal_22159) ) ;
    buf_clk cell_17277 ( .C (clk), .D (signal_22164), .Q (signal_22165) ) ;
    buf_clk cell_17283 ( .C (clk), .D (signal_22170), .Q (signal_22171) ) ;
    buf_clk cell_17289 ( .C (clk), .D (signal_22176), .Q (signal_22177) ) ;
    buf_clk cell_17295 ( .C (clk), .D (signal_22182), .Q (signal_22183) ) ;
    buf_clk cell_17301 ( .C (clk), .D (signal_22188), .Q (signal_22189) ) ;
    buf_clk cell_17307 ( .C (clk), .D (signal_22194), .Q (signal_22195) ) ;
    buf_clk cell_17313 ( .C (clk), .D (signal_22200), .Q (signal_22201) ) ;
    buf_clk cell_17319 ( .C (clk), .D (signal_22206), .Q (signal_22207) ) ;
    buf_clk cell_17325 ( .C (clk), .D (signal_22212), .Q (signal_22213) ) ;
    buf_clk cell_17331 ( .C (clk), .D (signal_22218), .Q (signal_22219) ) ;
    buf_clk cell_17337 ( .C (clk), .D (signal_22224), .Q (signal_22225) ) ;
    buf_clk cell_17343 ( .C (clk), .D (signal_22230), .Q (signal_22231) ) ;
    buf_clk cell_17349 ( .C (clk), .D (signal_22236), .Q (signal_22237) ) ;
    buf_clk cell_17355 ( .C (clk), .D (signal_22242), .Q (signal_22243) ) ;
    buf_clk cell_17361 ( .C (clk), .D (signal_22248), .Q (signal_22249) ) ;
    buf_clk cell_17367 ( .C (clk), .D (signal_22254), .Q (signal_22255) ) ;
    buf_clk cell_17373 ( .C (clk), .D (signal_22260), .Q (signal_22261) ) ;
    buf_clk cell_17379 ( .C (clk), .D (signal_22266), .Q (signal_22267) ) ;
    buf_clk cell_17385 ( .C (clk), .D (signal_22272), .Q (signal_22273) ) ;
    buf_clk cell_17391 ( .C (clk), .D (signal_22278), .Q (signal_22279) ) ;
    buf_clk cell_17397 ( .C (clk), .D (signal_22284), .Q (signal_22285) ) ;
    buf_clk cell_17403 ( .C (clk), .D (signal_22290), .Q (signal_22291) ) ;
    buf_clk cell_17409 ( .C (clk), .D (signal_22296), .Q (signal_22297) ) ;
    buf_clk cell_17415 ( .C (clk), .D (signal_22302), .Q (signal_22303) ) ;
    buf_clk cell_17421 ( .C (clk), .D (signal_22308), .Q (signal_22309) ) ;
    buf_clk cell_17427 ( .C (clk), .D (signal_22314), .Q (signal_22315) ) ;
    buf_clk cell_17433 ( .C (clk), .D (signal_22320), .Q (signal_22321) ) ;
    buf_clk cell_17439 ( .C (clk), .D (signal_22326), .Q (signal_22327) ) ;
    buf_clk cell_17445 ( .C (clk), .D (signal_22332), .Q (signal_22333) ) ;
    buf_clk cell_17451 ( .C (clk), .D (signal_22338), .Q (signal_22339) ) ;
    buf_clk cell_17457 ( .C (clk), .D (signal_22344), .Q (signal_22345) ) ;
    buf_clk cell_17463 ( .C (clk), .D (signal_22350), .Q (signal_22351) ) ;
    buf_clk cell_17469 ( .C (clk), .D (signal_22356), .Q (signal_22357) ) ;
    buf_clk cell_17475 ( .C (clk), .D (signal_22362), .Q (signal_22363) ) ;
    buf_clk cell_17481 ( .C (clk), .D (signal_22368), .Q (signal_22369) ) ;
    buf_clk cell_17487 ( .C (clk), .D (signal_22374), .Q (signal_22375) ) ;
    buf_clk cell_17493 ( .C (clk), .D (signal_22380), .Q (signal_22381) ) ;
    buf_clk cell_17499 ( .C (clk), .D (signal_22386), .Q (signal_22387) ) ;
    buf_clk cell_17505 ( .C (clk), .D (signal_22392), .Q (signal_22393) ) ;
    buf_clk cell_17511 ( .C (clk), .D (signal_22398), .Q (signal_22399) ) ;
    buf_clk cell_17517 ( .C (clk), .D (signal_22404), .Q (signal_22405) ) ;
    buf_clk cell_17523 ( .C (clk), .D (signal_22410), .Q (signal_22411) ) ;
    buf_clk cell_17529 ( .C (clk), .D (signal_22416), .Q (signal_22417) ) ;
    buf_clk cell_17535 ( .C (clk), .D (signal_22422), .Q (signal_22423) ) ;
    buf_clk cell_17541 ( .C (clk), .D (signal_22428), .Q (signal_22429) ) ;
    buf_clk cell_17547 ( .C (clk), .D (signal_22434), .Q (signal_22435) ) ;
    buf_clk cell_17553 ( .C (clk), .D (signal_22440), .Q (signal_22441) ) ;
    buf_clk cell_17559 ( .C (clk), .D (signal_22446), .Q (signal_22447) ) ;
    buf_clk cell_17565 ( .C (clk), .D (signal_22452), .Q (signal_22453) ) ;
    buf_clk cell_17571 ( .C (clk), .D (signal_22458), .Q (signal_22459) ) ;
    buf_clk cell_17577 ( .C (clk), .D (signal_22464), .Q (signal_22465) ) ;
    buf_clk cell_17583 ( .C (clk), .D (signal_22470), .Q (signal_22471) ) ;
    buf_clk cell_17589 ( .C (clk), .D (signal_22476), .Q (signal_22477) ) ;
    buf_clk cell_17597 ( .C (clk), .D (signal_22484), .Q (signal_22485) ) ;
    buf_clk cell_17605 ( .C (clk), .D (signal_22492), .Q (signal_22493) ) ;
    buf_clk cell_17613 ( .C (clk), .D (signal_22500), .Q (signal_22501) ) ;
    buf_clk cell_17621 ( .C (clk), .D (signal_22508), .Q (signal_22509) ) ;
    buf_clk cell_17629 ( .C (clk), .D (signal_22516), .Q (signal_22517) ) ;
    buf_clk cell_17637 ( .C (clk), .D (signal_22524), .Q (signal_22525) ) ;
    buf_clk cell_17645 ( .C (clk), .D (signal_22532), .Q (signal_22533) ) ;
    buf_clk cell_17653 ( .C (clk), .D (signal_22540), .Q (signal_22541) ) ;
    buf_clk cell_17661 ( .C (clk), .D (signal_22548), .Q (signal_22549) ) ;
    buf_clk cell_17669 ( .C (clk), .D (signal_22556), .Q (signal_22557) ) ;
    buf_clk cell_17677 ( .C (clk), .D (signal_22564), .Q (signal_22565) ) ;
    buf_clk cell_17685 ( .C (clk), .D (signal_22572), .Q (signal_22573) ) ;
    buf_clk cell_17693 ( .C (clk), .D (signal_22580), .Q (signal_22581) ) ;
    buf_clk cell_17701 ( .C (clk), .D (signal_22588), .Q (signal_22589) ) ;
    buf_clk cell_17709 ( .C (clk), .D (signal_22596), .Q (signal_22597) ) ;
    buf_clk cell_17717 ( .C (clk), .D (signal_22604), .Q (signal_22605) ) ;
    buf_clk cell_17725 ( .C (clk), .D (signal_22612), .Q (signal_22613) ) ;
    buf_clk cell_17733 ( .C (clk), .D (signal_22620), .Q (signal_22621) ) ;
    buf_clk cell_17741 ( .C (clk), .D (signal_22628), .Q (signal_22629) ) ;
    buf_clk cell_17749 ( .C (clk), .D (signal_22636), .Q (signal_22637) ) ;
    buf_clk cell_17757 ( .C (clk), .D (signal_22644), .Q (signal_22645) ) ;
    buf_clk cell_17765 ( .C (clk), .D (signal_22652), .Q (signal_22653) ) ;
    buf_clk cell_17773 ( .C (clk), .D (signal_22660), .Q (signal_22661) ) ;
    buf_clk cell_17781 ( .C (clk), .D (signal_22668), .Q (signal_22669) ) ;
    buf_clk cell_17789 ( .C (clk), .D (signal_22676), .Q (signal_22677) ) ;
    buf_clk cell_17797 ( .C (clk), .D (signal_22684), .Q (signal_22685) ) ;
    buf_clk cell_17805 ( .C (clk), .D (signal_22692), .Q (signal_22693) ) ;
    buf_clk cell_17813 ( .C (clk), .D (signal_22700), .Q (signal_22701) ) ;
    buf_clk cell_17821 ( .C (clk), .D (signal_22708), .Q (signal_22709) ) ;
    buf_clk cell_17829 ( .C (clk), .D (signal_22716), .Q (signal_22717) ) ;
    buf_clk cell_17837 ( .C (clk), .D (signal_22724), .Q (signal_22725) ) ;
    buf_clk cell_17845 ( .C (clk), .D (signal_22732), .Q (signal_22733) ) ;
    buf_clk cell_17853 ( .C (clk), .D (signal_22740), .Q (signal_22741) ) ;
    buf_clk cell_17861 ( .C (clk), .D (signal_22748), .Q (signal_22749) ) ;
    buf_clk cell_17869 ( .C (clk), .D (signal_22756), .Q (signal_22757) ) ;
    buf_clk cell_17877 ( .C (clk), .D (signal_22764), .Q (signal_22765) ) ;
    buf_clk cell_17885 ( .C (clk), .D (signal_22772), .Q (signal_22773) ) ;
    buf_clk cell_17893 ( .C (clk), .D (signal_22780), .Q (signal_22781) ) ;
    buf_clk cell_17901 ( .C (clk), .D (signal_22788), .Q (signal_22789) ) ;
    buf_clk cell_17909 ( .C (clk), .D (signal_22796), .Q (signal_22797) ) ;
    buf_clk cell_17917 ( .C (clk), .D (signal_22804), .Q (signal_22805) ) ;
    buf_clk cell_17925 ( .C (clk), .D (signal_22812), .Q (signal_22813) ) ;
    buf_clk cell_17933 ( .C (clk), .D (signal_22820), .Q (signal_22821) ) ;
    buf_clk cell_17941 ( .C (clk), .D (signal_22828), .Q (signal_22829) ) ;
    buf_clk cell_17949 ( .C (clk), .D (signal_22836), .Q (signal_22837) ) ;
    buf_clk cell_17957 ( .C (clk), .D (signal_22844), .Q (signal_22845) ) ;
    buf_clk cell_17965 ( .C (clk), .D (signal_22852), .Q (signal_22853) ) ;
    buf_clk cell_17973 ( .C (clk), .D (signal_22860), .Q (signal_22861) ) ;
    buf_clk cell_17981 ( .C (clk), .D (signal_22868), .Q (signal_22869) ) ;
    buf_clk cell_17989 ( .C (clk), .D (signal_22876), .Q (signal_22877) ) ;
    buf_clk cell_17997 ( .C (clk), .D (signal_22884), .Q (signal_22885) ) ;
    buf_clk cell_18005 ( .C (clk), .D (signal_22892), .Q (signal_22893) ) ;
    buf_clk cell_18013 ( .C (clk), .D (signal_22900), .Q (signal_22901) ) ;
    buf_clk cell_18021 ( .C (clk), .D (signal_22908), .Q (signal_22909) ) ;
    buf_clk cell_18029 ( .C (clk), .D (signal_22916), .Q (signal_22917) ) ;
    buf_clk cell_18037 ( .C (clk), .D (signal_22924), .Q (signal_22925) ) ;
    buf_clk cell_18045 ( .C (clk), .D (signal_22932), .Q (signal_22933) ) ;
    buf_clk cell_18053 ( .C (clk), .D (signal_22940), .Q (signal_22941) ) ;
    buf_clk cell_18061 ( .C (clk), .D (signal_22948), .Q (signal_22949) ) ;
    buf_clk cell_18069 ( .C (clk), .D (signal_22956), .Q (signal_22957) ) ;
    buf_clk cell_18077 ( .C (clk), .D (signal_22964), .Q (signal_22965) ) ;
    buf_clk cell_18085 ( .C (clk), .D (signal_22972), .Q (signal_22973) ) ;
    buf_clk cell_18093 ( .C (clk), .D (signal_22980), .Q (signal_22981) ) ;
    buf_clk cell_18101 ( .C (clk), .D (signal_22988), .Q (signal_22989) ) ;
    buf_clk cell_18109 ( .C (clk), .D (signal_22996), .Q (signal_22997) ) ;
    buf_clk cell_18117 ( .C (clk), .D (signal_23004), .Q (signal_23005) ) ;
    buf_clk cell_18125 ( .C (clk), .D (signal_23012), .Q (signal_23013) ) ;
    buf_clk cell_18133 ( .C (clk), .D (signal_23020), .Q (signal_23021) ) ;
    buf_clk cell_18141 ( .C (clk), .D (signal_23028), .Q (signal_23029) ) ;
    buf_clk cell_18149 ( .C (clk), .D (signal_23036), .Q (signal_23037) ) ;
    buf_clk cell_18157 ( .C (clk), .D (signal_23044), .Q (signal_23045) ) ;
    buf_clk cell_18165 ( .C (clk), .D (signal_23052), .Q (signal_23053) ) ;
    buf_clk cell_18173 ( .C (clk), .D (signal_23060), .Q (signal_23061) ) ;
    buf_clk cell_18181 ( .C (clk), .D (signal_23068), .Q (signal_23069) ) ;
    buf_clk cell_18189 ( .C (clk), .D (signal_23076), .Q (signal_23077) ) ;
    buf_clk cell_18197 ( .C (clk), .D (signal_23084), .Q (signal_23085) ) ;
    buf_clk cell_18205 ( .C (clk), .D (signal_23092), .Q (signal_23093) ) ;
    buf_clk cell_18213 ( .C (clk), .D (signal_23100), .Q (signal_23101) ) ;
    buf_clk cell_18221 ( .C (clk), .D (signal_23108), .Q (signal_23109) ) ;
    buf_clk cell_18229 ( .C (clk), .D (signal_23116), .Q (signal_23117) ) ;
    buf_clk cell_18237 ( .C (clk), .D (signal_23124), .Q (signal_23125) ) ;
    buf_clk cell_18245 ( .C (clk), .D (signal_23132), .Q (signal_23133) ) ;
    buf_clk cell_18253 ( .C (clk), .D (signal_23140), .Q (signal_23141) ) ;
    buf_clk cell_18261 ( .C (clk), .D (signal_23148), .Q (signal_23149) ) ;
    buf_clk cell_18269 ( .C (clk), .D (signal_23156), .Q (signal_23157) ) ;
    buf_clk cell_18277 ( .C (clk), .D (signal_23164), .Q (signal_23165) ) ;
    buf_clk cell_18285 ( .C (clk), .D (signal_23172), .Q (signal_23173) ) ;
    buf_clk cell_18293 ( .C (clk), .D (signal_23180), .Q (signal_23181) ) ;
    buf_clk cell_18301 ( .C (clk), .D (signal_23188), .Q (signal_23189) ) ;
    buf_clk cell_18309 ( .C (clk), .D (signal_23196), .Q (signal_23197) ) ;
    buf_clk cell_18317 ( .C (clk), .D (signal_23204), .Q (signal_23205) ) ;
    buf_clk cell_18325 ( .C (clk), .D (signal_23212), .Q (signal_23213) ) ;
    buf_clk cell_18333 ( .C (clk), .D (signal_23220), .Q (signal_23221) ) ;
    buf_clk cell_18341 ( .C (clk), .D (signal_23228), .Q (signal_23229) ) ;
    buf_clk cell_18349 ( .C (clk), .D (signal_23236), .Q (signal_23237) ) ;
    buf_clk cell_18357 ( .C (clk), .D (signal_23244), .Q (signal_23245) ) ;
    buf_clk cell_18365 ( .C (clk), .D (signal_23252), .Q (signal_23253) ) ;
    buf_clk cell_18373 ( .C (clk), .D (signal_23260), .Q (signal_23261) ) ;
    buf_clk cell_18381 ( .C (clk), .D (signal_23268), .Q (signal_23269) ) ;
    buf_clk cell_18389 ( .C (clk), .D (signal_23276), .Q (signal_23277) ) ;
    buf_clk cell_18397 ( .C (clk), .D (signal_23284), .Q (signal_23285) ) ;
    buf_clk cell_18409 ( .C (clk), .D (signal_23296), .Q (signal_23297) ) ;
    buf_clk cell_18417 ( .C (clk), .D (signal_23304), .Q (signal_23305) ) ;
    buf_clk cell_18425 ( .C (clk), .D (signal_23312), .Q (signal_23313) ) ;
    buf_clk cell_18433 ( .C (clk), .D (signal_23320), .Q (signal_23321) ) ;
    buf_clk cell_18441 ( .C (clk), .D (signal_23328), .Q (signal_23329) ) ;
    buf_clk cell_18449 ( .C (clk), .D (signal_23336), .Q (signal_23337) ) ;
    buf_clk cell_18457 ( .C (clk), .D (signal_23344), .Q (signal_23345) ) ;
    buf_clk cell_18465 ( .C (clk), .D (signal_23352), .Q (signal_23353) ) ;
    buf_clk cell_18473 ( .C (clk), .D (signal_23360), .Q (signal_23361) ) ;
    buf_clk cell_18481 ( .C (clk), .D (signal_23368), .Q (signal_23369) ) ;
    buf_clk cell_18489 ( .C (clk), .D (signal_23376), .Q (signal_23377) ) ;
    buf_clk cell_18497 ( .C (clk), .D (signal_23384), .Q (signal_23385) ) ;
    buf_clk cell_18505 ( .C (clk), .D (signal_23392), .Q (signal_23393) ) ;
    buf_clk cell_18513 ( .C (clk), .D (signal_23400), .Q (signal_23401) ) ;
    buf_clk cell_18521 ( .C (clk), .D (signal_23408), .Q (signal_23409) ) ;
    buf_clk cell_18529 ( .C (clk), .D (signal_23416), .Q (signal_23417) ) ;
    buf_clk cell_18537 ( .C (clk), .D (signal_23424), .Q (signal_23425) ) ;
    buf_clk cell_18545 ( .C (clk), .D (signal_23432), .Q (signal_23433) ) ;
    buf_clk cell_18553 ( .C (clk), .D (signal_23440), .Q (signal_23441) ) ;
    buf_clk cell_18561 ( .C (clk), .D (signal_23448), .Q (signal_23449) ) ;
    buf_clk cell_18569 ( .C (clk), .D (signal_23456), .Q (signal_23457) ) ;
    buf_clk cell_18577 ( .C (clk), .D (signal_23464), .Q (signal_23465) ) ;
    buf_clk cell_18585 ( .C (clk), .D (signal_23472), .Q (signal_23473) ) ;
    buf_clk cell_18593 ( .C (clk), .D (signal_23480), .Q (signal_23481) ) ;
    buf_clk cell_18601 ( .C (clk), .D (signal_23488), .Q (signal_23489) ) ;
    buf_clk cell_18609 ( .C (clk), .D (signal_23496), .Q (signal_23497) ) ;
    buf_clk cell_18617 ( .C (clk), .D (signal_23504), .Q (signal_23505) ) ;
    buf_clk cell_18625 ( .C (clk), .D (signal_23512), .Q (signal_23513) ) ;
    buf_clk cell_18633 ( .C (clk), .D (signal_23520), .Q (signal_23521) ) ;
    buf_clk cell_18641 ( .C (clk), .D (signal_23528), .Q (signal_23529) ) ;
    buf_clk cell_18653 ( .C (clk), .D (signal_23540), .Q (signal_23541) ) ;
    buf_clk cell_18661 ( .C (clk), .D (signal_23548), .Q (signal_23549) ) ;
    buf_clk cell_18669 ( .C (clk), .D (signal_23556), .Q (signal_23557) ) ;
    buf_clk cell_18677 ( .C (clk), .D (signal_23564), .Q (signal_23565) ) ;
    buf_clk cell_18685 ( .C (clk), .D (signal_23572), .Q (signal_23573) ) ;
    buf_clk cell_18693 ( .C (clk), .D (signal_23580), .Q (signal_23581) ) ;
    buf_clk cell_18701 ( .C (clk), .D (signal_23588), .Q (signal_23589) ) ;
    buf_clk cell_18709 ( .C (clk), .D (signal_23596), .Q (signal_23597) ) ;
    buf_clk cell_18717 ( .C (clk), .D (signal_23604), .Q (signal_23605) ) ;
    buf_clk cell_18725 ( .C (clk), .D (signal_23612), .Q (signal_23613) ) ;
    buf_clk cell_18733 ( .C (clk), .D (signal_23620), .Q (signal_23621) ) ;
    buf_clk cell_18741 ( .C (clk), .D (signal_23628), .Q (signal_23629) ) ;
    buf_clk cell_18753 ( .C (clk), .D (signal_23640), .Q (signal_23641) ) ;
    buf_clk cell_18761 ( .C (clk), .D (signal_23648), .Q (signal_23649) ) ;
    buf_clk cell_18769 ( .C (clk), .D (signal_23656), .Q (signal_23657) ) ;
    buf_clk cell_18777 ( .C (clk), .D (signal_23664), .Q (signal_23665) ) ;
    buf_clk cell_18785 ( .C (clk), .D (signal_23672), .Q (signal_23673) ) ;
    buf_clk cell_18793 ( .C (clk), .D (signal_23680), .Q (signal_23681) ) ;
    buf_clk cell_18801 ( .C (clk), .D (signal_23688), .Q (signal_23689) ) ;
    buf_clk cell_18809 ( .C (clk), .D (signal_23696), .Q (signal_23697) ) ;
    buf_clk cell_18817 ( .C (clk), .D (signal_23704), .Q (signal_23705) ) ;
    buf_clk cell_18825 ( .C (clk), .D (signal_23712), .Q (signal_23713) ) ;
    buf_clk cell_18833 ( .C (clk), .D (signal_23720), .Q (signal_23721) ) ;
    buf_clk cell_18841 ( .C (clk), .D (signal_23728), .Q (signal_23729) ) ;
    buf_clk cell_18849 ( .C (clk), .D (signal_23736), .Q (signal_23737) ) ;
    buf_clk cell_18857 ( .C (clk), .D (signal_23744), .Q (signal_23745) ) ;
    buf_clk cell_18865 ( .C (clk), .D (signal_23752), .Q (signal_23753) ) ;
    buf_clk cell_18873 ( .C (clk), .D (signal_23760), .Q (signal_23761) ) ;
    buf_clk cell_18881 ( .C (clk), .D (signal_23768), .Q (signal_23769) ) ;
    buf_clk cell_18889 ( .C (clk), .D (signal_23776), .Q (signal_23777) ) ;
    buf_clk cell_18897 ( .C (clk), .D (signal_23784), .Q (signal_23785) ) ;
    buf_clk cell_18905 ( .C (clk), .D (signal_23792), .Q (signal_23793) ) ;
    buf_clk cell_18913 ( .C (clk), .D (signal_23800), .Q (signal_23801) ) ;
    buf_clk cell_18921 ( .C (clk), .D (signal_23808), .Q (signal_23809) ) ;
    buf_clk cell_18929 ( .C (clk), .D (signal_23816), .Q (signal_23817) ) ;
    buf_clk cell_18937 ( .C (clk), .D (signal_23824), .Q (signal_23825) ) ;
    buf_clk cell_18945 ( .C (clk), .D (signal_23832), .Q (signal_23833) ) ;
    buf_clk cell_18953 ( .C (clk), .D (signal_23840), .Q (signal_23841) ) ;
    buf_clk cell_18961 ( .C (clk), .D (signal_23848), .Q (signal_23849) ) ;
    buf_clk cell_18969 ( .C (clk), .D (signal_23856), .Q (signal_23857) ) ;
    buf_clk cell_18977 ( .C (clk), .D (signal_23864), .Q (signal_23865) ) ;
    buf_clk cell_18985 ( .C (clk), .D (signal_23872), .Q (signal_23873) ) ;
    buf_clk cell_18993 ( .C (clk), .D (signal_23880), .Q (signal_23881) ) ;
    buf_clk cell_19001 ( .C (clk), .D (signal_23888), .Q (signal_23889) ) ;
    buf_clk cell_19009 ( .C (clk), .D (signal_23896), .Q (signal_23897) ) ;
    buf_clk cell_19017 ( .C (clk), .D (signal_23904), .Q (signal_23905) ) ;
    buf_clk cell_19025 ( .C (clk), .D (signal_23912), .Q (signal_23913) ) ;
    buf_clk cell_19033 ( .C (clk), .D (signal_23920), .Q (signal_23921) ) ;
    buf_clk cell_19041 ( .C (clk), .D (signal_23928), .Q (signal_23929) ) ;
    buf_clk cell_19049 ( .C (clk), .D (signal_23936), .Q (signal_23937) ) ;
    buf_clk cell_19057 ( .C (clk), .D (signal_23944), .Q (signal_23945) ) ;
    buf_clk cell_19065 ( .C (clk), .D (signal_23952), .Q (signal_23953) ) ;
    buf_clk cell_19073 ( .C (clk), .D (signal_23960), .Q (signal_23961) ) ;
    buf_clk cell_19081 ( .C (clk), .D (signal_23968), .Q (signal_23969) ) ;
    buf_clk cell_19089 ( .C (clk), .D (signal_23976), .Q (signal_23977) ) ;
    buf_clk cell_19097 ( .C (clk), .D (signal_23984), .Q (signal_23985) ) ;
    buf_clk cell_19105 ( .C (clk), .D (signal_23992), .Q (signal_23993) ) ;
    buf_clk cell_19113 ( .C (clk), .D (signal_24000), .Q (signal_24001) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5415 ( .a ({signal_12800, signal_12798}), .b ({signal_8926, signal_5606}), .clk (clk), .r (Fresh[240]), .c ({signal_9021, signal_5651}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5416 ( .a ({signal_12960, signal_12958}), .b ({signal_8925, signal_5605}), .clk (clk), .r (Fresh[241]), .c ({signal_9022, signal_5652}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5417 ( .a ({signal_12800, signal_12798}), .b ({signal_8921, signal_5571}), .clk (clk), .r (Fresh[242]), .c ({signal_9023, signal_5653}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5418 ( .a ({signal_8838, signal_5478}), .b ({signal_12960, signal_12958}), .clk (clk), .r (Fresh[243]), .c ({signal_9024, signal_5654}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5422 ( .a ({signal_12812, signal_12810}), .b ({signal_8930, signal_5616}), .clk (clk), .r (Fresh[244]), .c ({signal_9025, signal_5658}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5423 ( .a ({signal_13000, signal_12998}), .b ({signal_8929, signal_5615}), .clk (clk), .r (Fresh[245]), .c ({signal_9026, signal_5659}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5424 ( .a ({signal_12812, signal_12810}), .b ({signal_8922, signal_5578}), .clk (clk), .r (Fresh[246]), .c ({signal_9027, signal_5660}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5425 ( .a ({signal_8840, signal_5480}), .b ({signal_13000, signal_12998}), .clk (clk), .r (Fresh[247]), .c ({signal_9028, signal_5661}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5429 ( .a ({signal_12824, signal_12822}), .b ({signal_8934, signal_5626}), .clk (clk), .r (Fresh[248]), .c ({signal_9029, signal_5665}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5430 ( .a ({signal_13040, signal_13038}), .b ({signal_8933, signal_5625}), .clk (clk), .r (Fresh[249]), .c ({signal_9030, signal_5666}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5431 ( .a ({signal_12824, signal_12822}), .b ({signal_8923, signal_5585}), .clk (clk), .r (Fresh[250]), .c ({signal_9031, signal_5667}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5432 ( .a ({signal_8842, signal_5482}), .b ({signal_13040, signal_13038}), .clk (clk), .r (Fresh[251]), .c ({signal_9032, signal_5668}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5433 ( .a ({signal_12836, signal_12834}), .b ({signal_8907, signal_5630}), .clk (clk), .r (Fresh[252]), .c ({signal_8949, signal_5669}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5434 ( .a ({signal_13044, signal_13042}), .b ({signal_8906, signal_5629}), .clk (clk), .r (Fresh[253]), .c ({signal_8950, signal_5670}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5435 ( .a ({signal_12836, signal_12834}), .b ({signal_8875, signal_5586}), .clk (clk), .r (Fresh[254]), .c ({signal_8951, signal_5671}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5436 ( .a ({signal_8770, signal_5484}), .b ({signal_13044, signal_13042}), .clk (clk), .r (Fresh[255]), .c ({signal_8952, signal_5672}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5437 ( .a ({signal_12848, signal_12846}), .b ({signal_8911, signal_5634}), .clk (clk), .r (Fresh[256]), .c ({signal_8953, signal_5673}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5438 ( .a ({signal_13048, signal_13046}), .b ({signal_8910, signal_5633}), .clk (clk), .r (Fresh[257]), .c ({signal_8954, signal_5674}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5439 ( .a ({signal_12848, signal_12846}), .b ({signal_8876, signal_5587}), .clk (clk), .r (Fresh[258]), .c ({signal_8955, signal_5675}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5440 ( .a ({signal_8772, signal_5486}), .b ({signal_13048, signal_13046}), .clk (clk), .r (Fresh[259]), .c ({signal_8956, signal_5676}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5441 ( .a ({signal_12860, signal_12858}), .b ({signal_8915, signal_5638}), .clk (clk), .r (Fresh[260]), .c ({signal_8957, signal_5677}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5442 ( .a ({signal_13052, signal_13050}), .b ({signal_8914, signal_5637}), .clk (clk), .r (Fresh[261]), .c ({signal_8958, signal_5678}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5443 ( .a ({signal_12860, signal_12858}), .b ({signal_8877, signal_5588}), .clk (clk), .r (Fresh[262]), .c ({signal_8959, signal_5679}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5444 ( .a ({signal_8774, signal_5488}), .b ({signal_13052, signal_13050}), .clk (clk), .r (Fresh[263]), .c ({signal_8960, signal_5680}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5445 ( .a ({signal_12872, signal_12870}), .b ({signal_8919, signal_5642}), .clk (clk), .r (Fresh[264]), .c ({signal_8961, signal_5681}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5446 ( .a ({signal_13056, signal_13054}), .b ({signal_8918, signal_5641}), .clk (clk), .r (Fresh[265]), .c ({signal_8962, signal_5682}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5447 ( .a ({signal_12872, signal_12870}), .b ({signal_8878, signal_5589}), .clk (clk), .r (Fresh[266]), .c ({signal_8963, signal_5683}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5448 ( .a ({signal_8776, signal_5490}), .b ({signal_13056, signal_13054}), .clk (clk), .r (Fresh[267]), .c ({signal_8964, signal_5684}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5508 ( .a ({signal_12884, signal_12882}), .b ({signal_8967, signal_5687}), .clk (clk), .r (Fresh[268]), .c ({signal_9036, signal_5744}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5509 ( .a ({signal_13060, signal_13058}), .b ({signal_8966, signal_5686}), .clk (clk), .r (Fresh[269]), .c ({signal_9037, signal_5745}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5510 ( .a ({signal_12884, signal_12882}), .b ({signal_8936, signal_5644}), .clk (clk), .r (Fresh[270]), .c ({signal_9038, signal_5746}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5511 ( .a ({signal_8850, signal_5558}), .b ({signal_13060, signal_13058}), .clk (clk), .r (Fresh[271]), .c ({signal_9039, signal_5747}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5512 ( .a ({signal_12896, signal_12894}), .b ({signal_8971, signal_5691}), .clk (clk), .r (Fresh[272]), .c ({signal_9040, signal_5748}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5513 ( .a ({signal_13064, signal_13062}), .b ({signal_8970, signal_5690}), .clk (clk), .r (Fresh[273]), .c ({signal_9041, signal_5749}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5514 ( .a ({signal_12896, signal_12894}), .b ({signal_8937, signal_5645}), .clk (clk), .r (Fresh[274]), .c ({signal_9042, signal_5750}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5515 ( .a ({signal_8852, signal_5560}), .b ({signal_13064, signal_13062}), .clk (clk), .r (Fresh[275]), .c ({signal_9043, signal_5751}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5516 ( .a ({signal_12908, signal_12906}), .b ({signal_8975, signal_5695}), .clk (clk), .r (Fresh[276]), .c ({signal_9044, signal_5752}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5517 ( .a ({signal_13068, signal_13066}), .b ({signal_8974, signal_5694}), .clk (clk), .r (Fresh[277]), .c ({signal_9045, signal_5753}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5518 ( .a ({signal_12908, signal_12906}), .b ({signal_8938, signal_5646}), .clk (clk), .r (Fresh[278]), .c ({signal_9046, signal_5754}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5519 ( .a ({signal_8854, signal_5562}), .b ({signal_13068, signal_13066}), .clk (clk), .r (Fresh[279]), .c ({signal_9047, signal_5755}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5520 ( .a ({signal_12920, signal_12918}), .b ({signal_8979, signal_5699}), .clk (clk), .r (Fresh[280]), .c ({signal_9048, signal_5756}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5521 ( .a ({signal_13072, signal_13070}), .b ({signal_8978, signal_5698}), .clk (clk), .r (Fresh[281]), .c ({signal_9049, signal_5757}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5522 ( .a ({signal_12920, signal_12918}), .b ({signal_8939, signal_5647}), .clk (clk), .r (Fresh[282]), .c ({signal_9050, signal_5758}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5523 ( .a ({signal_8856, signal_5564}), .b ({signal_13072, signal_13070}), .clk (clk), .r (Fresh[283]), .c ({signal_9051, signal_5759}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5524 ( .a ({signal_12932, signal_12930}), .b ({signal_8983, signal_5703}), .clk (clk), .r (Fresh[284]), .c ({signal_9052, signal_5760}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5525 ( .a ({signal_13076, signal_13074}), .b ({signal_8982, signal_5702}), .clk (clk), .r (Fresh[285]), .c ({signal_9053, signal_5761}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5526 ( .a ({signal_12932, signal_12930}), .b ({signal_8940, signal_5648}), .clk (clk), .r (Fresh[286]), .c ({signal_9054, signal_5762}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5527 ( .a ({signal_8858, signal_5566}), .b ({signal_13076, signal_13074}), .clk (clk), .r (Fresh[287]), .c ({signal_9055, signal_5763}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5528 ( .a ({signal_12944, signal_12942}), .b ({signal_8987, signal_5707}), .clk (clk), .r (Fresh[288]), .c ({signal_9056, signal_5764}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5529 ( .a ({signal_13080, signal_13078}), .b ({signal_8986, signal_5706}), .clk (clk), .r (Fresh[289]), .c ({signal_9057, signal_5765}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5530 ( .a ({signal_12944, signal_12942}), .b ({signal_8941, signal_5649}), .clk (clk), .r (Fresh[290]), .c ({signal_9058, signal_5766}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5531 ( .a ({signal_8860, signal_5568}), .b ({signal_13080, signal_13078}), .clk (clk), .r (Fresh[291]), .c ({signal_9059, signal_5767}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5532 ( .a ({signal_12956, signal_12954}), .b ({signal_8991, signal_5711}), .clk (clk), .r (Fresh[292]), .c ({signal_9060, signal_5768}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5533 ( .a ({signal_13084, signal_13082}), .b ({signal_8990, signal_5710}), .clk (clk), .r (Fresh[293]), .c ({signal_9061, signal_5769}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5534 ( .a ({signal_12956, signal_12954}), .b ({signal_8942, signal_5650}), .clk (clk), .r (Fresh[294]), .c ({signal_9062, signal_5770}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5535 ( .a ({signal_8862, signal_5570}), .b ({signal_13084, signal_13082}), .clk (clk), .r (Fresh[295]), .c ({signal_9063, signal_5771}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5536 ( .a ({signal_12972, signal_12970}), .b ({signal_8995, signal_5716}), .clk (clk), .r (Fresh[296]), .c ({signal_9064, signal_5772}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5537 ( .a ({signal_13088, signal_13086}), .b ({signal_8994, signal_5715}), .clk (clk), .r (Fresh[297]), .c ({signal_9065, signal_5773}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5538 ( .a ({signal_12972, signal_12970}), .b ({signal_8943, signal_5655}), .clk (clk), .r (Fresh[298]), .c ({signal_9066, signal_5774}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5539 ( .a ({signal_8864, signal_5573}), .b ({signal_13088, signal_13086}), .clk (clk), .r (Fresh[299]), .c ({signal_9067, signal_5775}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5540 ( .a ({signal_12984, signal_12982}), .b ({signal_8999, signal_5720}), .clk (clk), .r (Fresh[300]), .c ({signal_9068, signal_5776}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5541 ( .a ({signal_13092, signal_13090}), .b ({signal_8998, signal_5719}), .clk (clk), .r (Fresh[301]), .c ({signal_9069, signal_5777}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5542 ( .a ({signal_12984, signal_12982}), .b ({signal_8944, signal_5656}), .clk (clk), .r (Fresh[302]), .c ({signal_9070, signal_5778}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5543 ( .a ({signal_8866, signal_5575}), .b ({signal_13092, signal_13090}), .clk (clk), .r (Fresh[303]), .c ({signal_9071, signal_5779}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5544 ( .a ({signal_12996, signal_12994}), .b ({signal_9003, signal_5724}), .clk (clk), .r (Fresh[304]), .c ({signal_9072, signal_5780}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5545 ( .a ({signal_13096, signal_13094}), .b ({signal_9002, signal_5723}), .clk (clk), .r (Fresh[305]), .c ({signal_9073, signal_5781}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5546 ( .a ({signal_12996, signal_12994}), .b ({signal_8945, signal_5657}), .clk (clk), .r (Fresh[306]), .c ({signal_9074, signal_5782}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5547 ( .a ({signal_8868, signal_5577}), .b ({signal_13096, signal_13094}), .clk (clk), .r (Fresh[307]), .c ({signal_9075, signal_5783}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5548 ( .a ({signal_13012, signal_13010}), .b ({signal_9007, signal_5729}), .clk (clk), .r (Fresh[308]), .c ({signal_9076, signal_5784}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5549 ( .a ({signal_13100, signal_13098}), .b ({signal_9006, signal_5728}), .clk (clk), .r (Fresh[309]), .c ({signal_9077, signal_5785}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5550 ( .a ({signal_13012, signal_13010}), .b ({signal_8946, signal_5662}), .clk (clk), .r (Fresh[310]), .c ({signal_9078, signal_5786}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5551 ( .a ({signal_8870, signal_5580}), .b ({signal_13100, signal_13098}), .clk (clk), .r (Fresh[311]), .c ({signal_9079, signal_5787}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5552 ( .a ({signal_13024, signal_13022}), .b ({signal_9011, signal_5733}), .clk (clk), .r (Fresh[312]), .c ({signal_9080, signal_5788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5553 ( .a ({signal_13104, signal_13102}), .b ({signal_9010, signal_5732}), .clk (clk), .r (Fresh[313]), .c ({signal_9081, signal_5789}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5554 ( .a ({signal_13024, signal_13022}), .b ({signal_8947, signal_5663}), .clk (clk), .r (Fresh[314]), .c ({signal_9082, signal_5790}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5555 ( .a ({signal_8872, signal_5582}), .b ({signal_13104, signal_13102}), .clk (clk), .r (Fresh[315]), .c ({signal_9083, signal_5791}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5556 ( .a ({signal_13036, signal_13034}), .b ({signal_9015, signal_5737}), .clk (clk), .r (Fresh[316]), .c ({signal_9084, signal_5792}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5557 ( .a ({signal_13108, signal_13106}), .b ({signal_9014, signal_5736}), .clk (clk), .r (Fresh[317]), .c ({signal_9085, signal_5793}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5558 ( .a ({signal_13036, signal_13034}), .b ({signal_8948, signal_5664}), .clk (clk), .r (Fresh[318]), .c ({signal_9086, signal_5794}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5559 ( .a ({signal_8874, signal_5584}), .b ({signal_13108, signal_13106}), .clk (clk), .r (Fresh[319]), .c ({signal_9087, signal_5795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5567 ( .a ({signal_13112, signal_13110}), .b ({signal_9021, signal_5651}), .c ({signal_9117, signal_5803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5568 ( .a ({signal_13116, signal_13114}), .b ({signal_9023, signal_5653}), .c ({signal_9118, signal_5804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5569 ( .a ({signal_13120, signal_13118}), .b ({signal_9022, signal_5652}), .c ({signal_9119, signal_5805}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5570 ( .a ({signal_9024, signal_5654}), .b ({signal_13124, signal_13122}), .c ({signal_9120, signal_5806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5574 ( .a ({signal_13128, signal_13126}), .b ({signal_9025, signal_5658}), .c ({signal_9121, signal_5810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5575 ( .a ({signal_13132, signal_13130}), .b ({signal_9027, signal_5660}), .c ({signal_9122, signal_5811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5576 ( .a ({signal_13136, signal_13134}), .b ({signal_9026, signal_5659}), .c ({signal_9123, signal_5812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5577 ( .a ({signal_9028, signal_5661}), .b ({signal_13140, signal_13138}), .c ({signal_9124, signal_5813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5581 ( .a ({signal_13144, signal_13142}), .b ({signal_9029, signal_5665}), .c ({signal_9125, signal_5817}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5582 ( .a ({signal_13148, signal_13146}), .b ({signal_9031, signal_5667}), .c ({signal_9126, signal_5818}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5583 ( .a ({signal_13152, signal_13150}), .b ({signal_9030, signal_5666}), .c ({signal_9127, signal_5819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5584 ( .a ({signal_9032, signal_5668}), .b ({signal_13156, signal_13154}), .c ({signal_9128, signal_5820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5585 ( .a ({signal_13160, signal_13158}), .b ({signal_8949, signal_5669}), .c ({signal_9101, signal_5821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5586 ( .a ({signal_13164, signal_13162}), .b ({signal_8951, signal_5671}), .c ({signal_9102, signal_5822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5587 ( .a ({signal_13168, signal_13166}), .b ({signal_8950, signal_5670}), .c ({signal_9103, signal_5823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5588 ( .a ({signal_8952, signal_5672}), .b ({signal_13172, signal_13170}), .c ({signal_9104, signal_5824}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5589 ( .a ({signal_13176, signal_13174}), .b ({signal_8953, signal_5673}), .c ({signal_9105, signal_5825}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5590 ( .a ({signal_13180, signal_13178}), .b ({signal_8955, signal_5675}), .c ({signal_9106, signal_5826}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5591 ( .a ({signal_13184, signal_13182}), .b ({signal_8954, signal_5674}), .c ({signal_9107, signal_5827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5592 ( .a ({signal_8956, signal_5676}), .b ({signal_13188, signal_13186}), .c ({signal_9108, signal_5828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5593 ( .a ({signal_13192, signal_13190}), .b ({signal_8957, signal_5677}), .c ({signal_9109, signal_5829}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5594 ( .a ({signal_13196, signal_13194}), .b ({signal_8959, signal_5679}), .c ({signal_9110, signal_5830}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5595 ( .a ({signal_13200, signal_13198}), .b ({signal_8958, signal_5678}), .c ({signal_9111, signal_5831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5596 ( .a ({signal_8960, signal_5680}), .b ({signal_13204, signal_13202}), .c ({signal_9112, signal_5832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5597 ( .a ({signal_13208, signal_13206}), .b ({signal_8961, signal_5681}), .c ({signal_9113, signal_5833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5598 ( .a ({signal_13212, signal_13210}), .b ({signal_8963, signal_5683}), .c ({signal_9114, signal_5834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5599 ( .a ({signal_13216, signal_13214}), .b ({signal_8962, signal_5682}), .c ({signal_9115, signal_5835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5600 ( .a ({signal_8964, signal_5684}), .b ({signal_13220, signal_13218}), .c ({signal_9116, signal_5836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5657 ( .a ({signal_13224, signal_13222}), .b ({signal_9036, signal_5744}), .c ({signal_9161, signal_5893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5658 ( .a ({signal_13228, signal_13226}), .b ({signal_9038, signal_5746}), .c ({signal_9162, signal_5894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5659 ( .a ({signal_13232, signal_13230}), .b ({signal_9037, signal_5745}), .c ({signal_9163, signal_5895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5660 ( .a ({signal_9039, signal_5747}), .b ({signal_13236, signal_13234}), .c ({signal_9164, signal_5896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5661 ( .a ({signal_13240, signal_13238}), .b ({signal_9040, signal_5748}), .c ({signal_9165, signal_5897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5662 ( .a ({signal_13244, signal_13242}), .b ({signal_9042, signal_5750}), .c ({signal_9166, signal_5898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5663 ( .a ({signal_13248, signal_13246}), .b ({signal_9041, signal_5749}), .c ({signal_9167, signal_5899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5664 ( .a ({signal_9043, signal_5751}), .b ({signal_13252, signal_13250}), .c ({signal_9168, signal_5900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5665 ( .a ({signal_13256, signal_13254}), .b ({signal_9044, signal_5752}), .c ({signal_9169, signal_5901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5666 ( .a ({signal_13260, signal_13258}), .b ({signal_9046, signal_5754}), .c ({signal_9170, signal_5902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5667 ( .a ({signal_13264, signal_13262}), .b ({signal_9045, signal_5753}), .c ({signal_9171, signal_5903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5668 ( .a ({signal_9047, signal_5755}), .b ({signal_13268, signal_13266}), .c ({signal_9172, signal_5904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5669 ( .a ({signal_13272, signal_13270}), .b ({signal_9048, signal_5756}), .c ({signal_9173, signal_5905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5670 ( .a ({signal_13276, signal_13274}), .b ({signal_9050, signal_5758}), .c ({signal_9174, signal_5906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5671 ( .a ({signal_13280, signal_13278}), .b ({signal_9049, signal_5757}), .c ({signal_9175, signal_5907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5672 ( .a ({signal_9051, signal_5759}), .b ({signal_13284, signal_13282}), .c ({signal_9176, signal_5908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5673 ( .a ({signal_13288, signal_13286}), .b ({signal_9052, signal_5760}), .c ({signal_9177, signal_5909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5674 ( .a ({signal_13292, signal_13290}), .b ({signal_9054, signal_5762}), .c ({signal_9178, signal_5910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5675 ( .a ({signal_13296, signal_13294}), .b ({signal_9053, signal_5761}), .c ({signal_9179, signal_5911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5676 ( .a ({signal_9055, signal_5763}), .b ({signal_13300, signal_13298}), .c ({signal_9180, signal_5912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5677 ( .a ({signal_13304, signal_13302}), .b ({signal_9056, signal_5764}), .c ({signal_9181, signal_5913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5678 ( .a ({signal_13308, signal_13306}), .b ({signal_9058, signal_5766}), .c ({signal_9182, signal_5914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5679 ( .a ({signal_13312, signal_13310}), .b ({signal_9057, signal_5765}), .c ({signal_9183, signal_5915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5680 ( .a ({signal_9059, signal_5767}), .b ({signal_13316, signal_13314}), .c ({signal_9184, signal_5916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5681 ( .a ({signal_13320, signal_13318}), .b ({signal_9060, signal_5768}), .c ({signal_9185, signal_5917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5682 ( .a ({signal_13324, signal_13322}), .b ({signal_9062, signal_5770}), .c ({signal_9186, signal_5918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5683 ( .a ({signal_13328, signal_13326}), .b ({signal_9061, signal_5769}), .c ({signal_9187, signal_5919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5684 ( .a ({signal_9063, signal_5771}), .b ({signal_13332, signal_13330}), .c ({signal_9188, signal_5920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5685 ( .a ({signal_9118, signal_5804}), .b ({signal_9120, signal_5806}), .c ({signal_9253, signal_5921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5686 ( .a ({signal_9117, signal_5803}), .b ({signal_9119, signal_5805}), .c ({signal_9254, signal_5922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5687 ( .a ({signal_9117, signal_5803}), .b ({signal_9118, signal_5804}), .c ({signal_9255, signal_5923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5688 ( .a ({signal_9119, signal_5805}), .b ({signal_9120, signal_5806}), .c ({signal_9256, signal_5924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5689 ( .a ({signal_13336, signal_13334}), .b ({signal_9064, signal_5772}), .c ({signal_9189, signal_5925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5690 ( .a ({signal_13340, signal_13338}), .b ({signal_9066, signal_5774}), .c ({signal_9190, signal_5926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5691 ( .a ({signal_13344, signal_13342}), .b ({signal_9065, signal_5773}), .c ({signal_9191, signal_5927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5692 ( .a ({signal_9067, signal_5775}), .b ({signal_13348, signal_13346}), .c ({signal_9192, signal_5928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5693 ( .a ({signal_13352, signal_13350}), .b ({signal_9068, signal_5776}), .c ({signal_9193, signal_5929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5694 ( .a ({signal_13356, signal_13354}), .b ({signal_9070, signal_5778}), .c ({signal_9194, signal_5930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5695 ( .a ({signal_13360, signal_13358}), .b ({signal_9069, signal_5777}), .c ({signal_9195, signal_5931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5696 ( .a ({signal_9071, signal_5779}), .b ({signal_13364, signal_13362}), .c ({signal_9196, signal_5932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5697 ( .a ({signal_13368, signal_13366}), .b ({signal_9072, signal_5780}), .c ({signal_9197, signal_5933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5698 ( .a ({signal_13372, signal_13370}), .b ({signal_9074, signal_5782}), .c ({signal_9198, signal_5934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5699 ( .a ({signal_13376, signal_13374}), .b ({signal_9073, signal_5781}), .c ({signal_9199, signal_5935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5700 ( .a ({signal_9075, signal_5783}), .b ({signal_13380, signal_13378}), .c ({signal_9200, signal_5936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5701 ( .a ({signal_9122, signal_5811}), .b ({signal_9124, signal_5813}), .c ({signal_9257, signal_5937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5702 ( .a ({signal_9121, signal_5810}), .b ({signal_9123, signal_5812}), .c ({signal_9258, signal_5938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5703 ( .a ({signal_9121, signal_5810}), .b ({signal_9122, signal_5811}), .c ({signal_9259, signal_5939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5704 ( .a ({signal_9123, signal_5812}), .b ({signal_9124, signal_5813}), .c ({signal_9260, signal_5940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5705 ( .a ({signal_13384, signal_13382}), .b ({signal_9076, signal_5784}), .c ({signal_9201, signal_5941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5706 ( .a ({signal_13388, signal_13386}), .b ({signal_9078, signal_5786}), .c ({signal_9202, signal_5942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5707 ( .a ({signal_13392, signal_13390}), .b ({signal_9077, signal_5785}), .c ({signal_9203, signal_5943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5708 ( .a ({signal_9079, signal_5787}), .b ({signal_13396, signal_13394}), .c ({signal_9204, signal_5944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5709 ( .a ({signal_13400, signal_13398}), .b ({signal_9080, signal_5788}), .c ({signal_9205, signal_5945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5710 ( .a ({signal_13404, signal_13402}), .b ({signal_9082, signal_5790}), .c ({signal_9206, signal_5946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5711 ( .a ({signal_13408, signal_13406}), .b ({signal_9081, signal_5789}), .c ({signal_9207, signal_5947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5712 ( .a ({signal_9083, signal_5791}), .b ({signal_13412, signal_13410}), .c ({signal_9208, signal_5948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5713 ( .a ({signal_13416, signal_13414}), .b ({signal_9084, signal_5792}), .c ({signal_9209, signal_5949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5714 ( .a ({signal_13420, signal_13418}), .b ({signal_9086, signal_5794}), .c ({signal_9210, signal_5950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5715 ( .a ({signal_13424, signal_13422}), .b ({signal_9085, signal_5793}), .c ({signal_9211, signal_5951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5716 ( .a ({signal_9087, signal_5795}), .b ({signal_13428, signal_13426}), .c ({signal_9212, signal_5952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5717 ( .a ({signal_9126, signal_5818}), .b ({signal_9128, signal_5820}), .c ({signal_9261, signal_5953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5718 ( .a ({signal_9125, signal_5817}), .b ({signal_9127, signal_5819}), .c ({signal_9262, signal_5954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5719 ( .a ({signal_9125, signal_5817}), .b ({signal_9126, signal_5818}), .c ({signal_9263, signal_5955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5720 ( .a ({signal_9127, signal_5819}), .b ({signal_9128, signal_5820}), .c ({signal_9264, signal_5956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5721 ( .a ({signal_9102, signal_5822}), .b ({signal_9104, signal_5824}), .c ({signal_9213, signal_5957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5722 ( .a ({signal_9101, signal_5821}), .b ({signal_9103, signal_5823}), .c ({signal_9214, signal_5958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5723 ( .a ({signal_9101, signal_5821}), .b ({signal_9102, signal_5822}), .c ({signal_9215, signal_5959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5724 ( .a ({signal_9103, signal_5823}), .b ({signal_9104, signal_5824}), .c ({signal_9216, signal_5960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5725 ( .a ({signal_9106, signal_5826}), .b ({signal_9108, signal_5828}), .c ({signal_9217, signal_5961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5726 ( .a ({signal_9105, signal_5825}), .b ({signal_9107, signal_5827}), .c ({signal_9218, signal_5962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5727 ( .a ({signal_9105, signal_5825}), .b ({signal_9106, signal_5826}), .c ({signal_9219, signal_5963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5728 ( .a ({signal_9107, signal_5827}), .b ({signal_9108, signal_5828}), .c ({signal_9220, signal_5964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5729 ( .a ({signal_9110, signal_5830}), .b ({signal_9112, signal_5832}), .c ({signal_9221, signal_5965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5730 ( .a ({signal_9109, signal_5829}), .b ({signal_9111, signal_5831}), .c ({signal_9222, signal_5966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5731 ( .a ({signal_9109, signal_5829}), .b ({signal_9110, signal_5830}), .c ({signal_9223, signal_5967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5732 ( .a ({signal_9111, signal_5831}), .b ({signal_9112, signal_5832}), .c ({signal_9224, signal_5968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5733 ( .a ({signal_9114, signal_5834}), .b ({signal_9116, signal_5836}), .c ({signal_9225, signal_5969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5734 ( .a ({signal_9113, signal_5833}), .b ({signal_9115, signal_5835}), .c ({signal_9226, signal_5970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5735 ( .a ({signal_9113, signal_5833}), .b ({signal_9114, signal_5834}), .c ({signal_9227, signal_5971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5736 ( .a ({signal_9115, signal_5835}), .b ({signal_9116, signal_5836}), .c ({signal_9228, signal_5972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5897 ( .a ({signal_9162, signal_5894}), .b ({signal_9164, signal_5896}), .c ({signal_9401, signal_6133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5898 ( .a ({signal_9161, signal_5893}), .b ({signal_9163, signal_5895}), .c ({signal_9402, signal_6134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5899 ( .a ({signal_9161, signal_5893}), .b ({signal_9162, signal_5894}), .c ({signal_9403, signal_6135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5900 ( .a ({signal_9163, signal_5895}), .b ({signal_9164, signal_5896}), .c ({signal_9404, signal_6136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5901 ( .a ({signal_9166, signal_5898}), .b ({signal_9168, signal_5900}), .c ({signal_9405, signal_6137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5902 ( .a ({signal_9165, signal_5897}), .b ({signal_9167, signal_5899}), .c ({signal_9406, signal_6138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5903 ( .a ({signal_9165, signal_5897}), .b ({signal_9166, signal_5898}), .c ({signal_9407, signal_6139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5904 ( .a ({signal_9167, signal_5899}), .b ({signal_9168, signal_5900}), .c ({signal_9408, signal_6140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5905 ( .a ({signal_9170, signal_5902}), .b ({signal_9172, signal_5904}), .c ({signal_9409, signal_6141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5906 ( .a ({signal_9169, signal_5901}), .b ({signal_9171, signal_5903}), .c ({signal_9410, signal_6142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5907 ( .a ({signal_9169, signal_5901}), .b ({signal_9170, signal_5902}), .c ({signal_9411, signal_6143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5908 ( .a ({signal_9171, signal_5903}), .b ({signal_9172, signal_5904}), .c ({signal_9412, signal_6144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5909 ( .a ({signal_9174, signal_5906}), .b ({signal_9176, signal_5908}), .c ({signal_9413, signal_6145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5910 ( .a ({signal_9173, signal_5905}), .b ({signal_9175, signal_5907}), .c ({signal_9414, signal_6146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5911 ( .a ({signal_9173, signal_5905}), .b ({signal_9174, signal_5906}), .c ({signal_9415, signal_6147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5912 ( .a ({signal_9175, signal_5907}), .b ({signal_9176, signal_5908}), .c ({signal_9416, signal_6148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5913 ( .a ({signal_9178, signal_5910}), .b ({signal_9180, signal_5912}), .c ({signal_9417, signal_6149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5914 ( .a ({signal_9177, signal_5909}), .b ({signal_9179, signal_5911}), .c ({signal_9418, signal_6150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5915 ( .a ({signal_9177, signal_5909}), .b ({signal_9178, signal_5910}), .c ({signal_9419, signal_6151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5916 ( .a ({signal_9179, signal_5911}), .b ({signal_9180, signal_5912}), .c ({signal_9420, signal_6152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5917 ( .a ({signal_9182, signal_5914}), .b ({signal_9184, signal_5916}), .c ({signal_9421, signal_6153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5918 ( .a ({signal_9181, signal_5913}), .b ({signal_9183, signal_5915}), .c ({signal_9422, signal_6154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5919 ( .a ({signal_9181, signal_5913}), .b ({signal_9182, signal_5914}), .c ({signal_9423, signal_6155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5920 ( .a ({signal_9183, signal_5915}), .b ({signal_9184, signal_5916}), .c ({signal_9424, signal_6156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5921 ( .a ({signal_9186, signal_5918}), .b ({signal_9188, signal_5920}), .c ({signal_9425, signal_6157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5922 ( .a ({signal_9185, signal_5917}), .b ({signal_9187, signal_5919}), .c ({signal_9426, signal_6158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5923 ( .a ({signal_9185, signal_5917}), .b ({signal_9186, signal_5918}), .c ({signal_9427, signal_6159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5924 ( .a ({signal_9187, signal_5919}), .b ({signal_9188, signal_5920}), .c ({signal_9428, signal_6160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5925 ( .a ({signal_9253, signal_5921}), .b ({signal_9254, signal_5922}), .c ({signal_9493, signal_6161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5929 ( .a ({signal_9190, signal_5926}), .b ({signal_9192, signal_5928}), .c ({signal_9429, signal_6165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5930 ( .a ({signal_9189, signal_5925}), .b ({signal_9191, signal_5927}), .c ({signal_9430, signal_6166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5931 ( .a ({signal_9189, signal_5925}), .b ({signal_9190, signal_5926}), .c ({signal_9431, signal_6167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5932 ( .a ({signal_9191, signal_5927}), .b ({signal_9192, signal_5928}), .c ({signal_9432, signal_6168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5933 ( .a ({signal_9194, signal_5930}), .b ({signal_9196, signal_5932}), .c ({signal_9433, signal_6169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5934 ( .a ({signal_9193, signal_5929}), .b ({signal_9195, signal_5931}), .c ({signal_9434, signal_6170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5935 ( .a ({signal_9193, signal_5929}), .b ({signal_9194, signal_5930}), .c ({signal_9435, signal_6171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5936 ( .a ({signal_9195, signal_5931}), .b ({signal_9196, signal_5932}), .c ({signal_9436, signal_6172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5937 ( .a ({signal_9198, signal_5934}), .b ({signal_9200, signal_5936}), .c ({signal_9437, signal_6173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5938 ( .a ({signal_9197, signal_5933}), .b ({signal_9199, signal_5935}), .c ({signal_9438, signal_6174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5939 ( .a ({signal_9197, signal_5933}), .b ({signal_9198, signal_5934}), .c ({signal_9439, signal_6175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5940 ( .a ({signal_9199, signal_5935}), .b ({signal_9200, signal_5936}), .c ({signal_9440, signal_6176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5941 ( .a ({signal_9257, signal_5937}), .b ({signal_9258, signal_5938}), .c ({signal_9497, signal_6177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5945 ( .a ({signal_9202, signal_5942}), .b ({signal_9204, signal_5944}), .c ({signal_9441, signal_6181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5946 ( .a ({signal_9201, signal_5941}), .b ({signal_9203, signal_5943}), .c ({signal_9442, signal_6182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5947 ( .a ({signal_9201, signal_5941}), .b ({signal_9202, signal_5942}), .c ({signal_9443, signal_6183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5948 ( .a ({signal_9203, signal_5943}), .b ({signal_9204, signal_5944}), .c ({signal_9444, signal_6184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5949 ( .a ({signal_9206, signal_5946}), .b ({signal_9208, signal_5948}), .c ({signal_9445, signal_6185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5950 ( .a ({signal_9205, signal_5945}), .b ({signal_9207, signal_5947}), .c ({signal_9446, signal_6186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5951 ( .a ({signal_9205, signal_5945}), .b ({signal_9206, signal_5946}), .c ({signal_9447, signal_6187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5952 ( .a ({signal_9207, signal_5947}), .b ({signal_9208, signal_5948}), .c ({signal_9448, signal_6188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5953 ( .a ({signal_9210, signal_5950}), .b ({signal_9212, signal_5952}), .c ({signal_9449, signal_6189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5954 ( .a ({signal_9209, signal_5949}), .b ({signal_9211, signal_5951}), .c ({signal_9450, signal_6190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5955 ( .a ({signal_9209, signal_5949}), .b ({signal_9210, signal_5950}), .c ({signal_9451, signal_6191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5956 ( .a ({signal_9211, signal_5951}), .b ({signal_9212, signal_5952}), .c ({signal_9452, signal_6192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5957 ( .a ({signal_9261, signal_5953}), .b ({signal_9262, signal_5954}), .c ({signal_9501, signal_6193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5961 ( .a ({signal_9213, signal_5957}), .b ({signal_9214, signal_5958}), .c ({signal_9453, signal_6197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5965 ( .a ({signal_9217, signal_5961}), .b ({signal_9218, signal_5962}), .c ({signal_9457, signal_6201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5969 ( .a ({signal_9221, signal_5965}), .b ({signal_9222, signal_5966}), .c ({signal_9461, signal_6205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5973 ( .a ({signal_9225, signal_5969}), .b ({signal_9226, signal_5970}), .c ({signal_9465, signal_6209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6095 ( .a ({signal_9401, signal_6133}), .b ({signal_9402, signal_6134}), .c ({signal_9617, signal_6331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6099 ( .a ({signal_9405, signal_6137}), .b ({signal_9406, signal_6138}), .c ({signal_9621, signal_6335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6103 ( .a ({signal_9409, signal_6141}), .b ({signal_9410, signal_6142}), .c ({signal_9625, signal_6339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6107 ( .a ({signal_9413, signal_6145}), .b ({signal_9414, signal_6146}), .c ({signal_9629, signal_6343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6111 ( .a ({signal_9417, signal_6149}), .b ({signal_9418, signal_6150}), .c ({signal_9633, signal_6347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6115 ( .a ({signal_9421, signal_6153}), .b ({signal_9422, signal_6154}), .c ({signal_9637, signal_6351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6119 ( .a ({signal_9425, signal_6157}), .b ({signal_9426, signal_6158}), .c ({signal_9641, signal_6355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6131 ( .a ({signal_9429, signal_6165}), .b ({signal_9430, signal_6166}), .c ({signal_9645, signal_6367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6135 ( .a ({signal_9433, signal_6169}), .b ({signal_9434, signal_6170}), .c ({signal_9649, signal_6371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6139 ( .a ({signal_9437, signal_6173}), .b ({signal_9438, signal_6174}), .c ({signal_9653, signal_6375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6151 ( .a ({signal_9441, signal_6181}), .b ({signal_9442, signal_6182}), .c ({signal_9657, signal_6387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6155 ( .a ({signal_9445, signal_6185}), .b ({signal_9446, signal_6186}), .c ({signal_9661, signal_6391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6159 ( .a ({signal_9449, signal_6189}), .b ({signal_9450, signal_6190}), .c ({signal_9665, signal_6395}) ) ;
    buf_clk cell_8222 ( .C (clk), .D (signal_13109), .Q (signal_13110) ) ;
    buf_clk cell_8224 ( .C (clk), .D (signal_13111), .Q (signal_13112) ) ;
    buf_clk cell_8226 ( .C (clk), .D (signal_13113), .Q (signal_13114) ) ;
    buf_clk cell_8228 ( .C (clk), .D (signal_13115), .Q (signal_13116) ) ;
    buf_clk cell_8230 ( .C (clk), .D (signal_13117), .Q (signal_13118) ) ;
    buf_clk cell_8232 ( .C (clk), .D (signal_13119), .Q (signal_13120) ) ;
    buf_clk cell_8234 ( .C (clk), .D (signal_13121), .Q (signal_13122) ) ;
    buf_clk cell_8236 ( .C (clk), .D (signal_13123), .Q (signal_13124) ) ;
    buf_clk cell_8238 ( .C (clk), .D (signal_13125), .Q (signal_13126) ) ;
    buf_clk cell_8240 ( .C (clk), .D (signal_13127), .Q (signal_13128) ) ;
    buf_clk cell_8242 ( .C (clk), .D (signal_13129), .Q (signal_13130) ) ;
    buf_clk cell_8244 ( .C (clk), .D (signal_13131), .Q (signal_13132) ) ;
    buf_clk cell_8246 ( .C (clk), .D (signal_13133), .Q (signal_13134) ) ;
    buf_clk cell_8248 ( .C (clk), .D (signal_13135), .Q (signal_13136) ) ;
    buf_clk cell_8250 ( .C (clk), .D (signal_13137), .Q (signal_13138) ) ;
    buf_clk cell_8252 ( .C (clk), .D (signal_13139), .Q (signal_13140) ) ;
    buf_clk cell_8254 ( .C (clk), .D (signal_13141), .Q (signal_13142) ) ;
    buf_clk cell_8256 ( .C (clk), .D (signal_13143), .Q (signal_13144) ) ;
    buf_clk cell_8258 ( .C (clk), .D (signal_13145), .Q (signal_13146) ) ;
    buf_clk cell_8260 ( .C (clk), .D (signal_13147), .Q (signal_13148) ) ;
    buf_clk cell_8262 ( .C (clk), .D (signal_13149), .Q (signal_13150) ) ;
    buf_clk cell_8264 ( .C (clk), .D (signal_13151), .Q (signal_13152) ) ;
    buf_clk cell_8266 ( .C (clk), .D (signal_13153), .Q (signal_13154) ) ;
    buf_clk cell_8268 ( .C (clk), .D (signal_13155), .Q (signal_13156) ) ;
    buf_clk cell_8270 ( .C (clk), .D (signal_13157), .Q (signal_13158) ) ;
    buf_clk cell_8272 ( .C (clk), .D (signal_13159), .Q (signal_13160) ) ;
    buf_clk cell_8274 ( .C (clk), .D (signal_13161), .Q (signal_13162) ) ;
    buf_clk cell_8276 ( .C (clk), .D (signal_13163), .Q (signal_13164) ) ;
    buf_clk cell_8278 ( .C (clk), .D (signal_13165), .Q (signal_13166) ) ;
    buf_clk cell_8280 ( .C (clk), .D (signal_13167), .Q (signal_13168) ) ;
    buf_clk cell_8282 ( .C (clk), .D (signal_13169), .Q (signal_13170) ) ;
    buf_clk cell_8284 ( .C (clk), .D (signal_13171), .Q (signal_13172) ) ;
    buf_clk cell_8286 ( .C (clk), .D (signal_13173), .Q (signal_13174) ) ;
    buf_clk cell_8288 ( .C (clk), .D (signal_13175), .Q (signal_13176) ) ;
    buf_clk cell_8290 ( .C (clk), .D (signal_13177), .Q (signal_13178) ) ;
    buf_clk cell_8292 ( .C (clk), .D (signal_13179), .Q (signal_13180) ) ;
    buf_clk cell_8294 ( .C (clk), .D (signal_13181), .Q (signal_13182) ) ;
    buf_clk cell_8296 ( .C (clk), .D (signal_13183), .Q (signal_13184) ) ;
    buf_clk cell_8298 ( .C (clk), .D (signal_13185), .Q (signal_13186) ) ;
    buf_clk cell_8300 ( .C (clk), .D (signal_13187), .Q (signal_13188) ) ;
    buf_clk cell_8302 ( .C (clk), .D (signal_13189), .Q (signal_13190) ) ;
    buf_clk cell_8304 ( .C (clk), .D (signal_13191), .Q (signal_13192) ) ;
    buf_clk cell_8306 ( .C (clk), .D (signal_13193), .Q (signal_13194) ) ;
    buf_clk cell_8308 ( .C (clk), .D (signal_13195), .Q (signal_13196) ) ;
    buf_clk cell_8310 ( .C (clk), .D (signal_13197), .Q (signal_13198) ) ;
    buf_clk cell_8312 ( .C (clk), .D (signal_13199), .Q (signal_13200) ) ;
    buf_clk cell_8314 ( .C (clk), .D (signal_13201), .Q (signal_13202) ) ;
    buf_clk cell_8316 ( .C (clk), .D (signal_13203), .Q (signal_13204) ) ;
    buf_clk cell_8318 ( .C (clk), .D (signal_13205), .Q (signal_13206) ) ;
    buf_clk cell_8320 ( .C (clk), .D (signal_13207), .Q (signal_13208) ) ;
    buf_clk cell_8322 ( .C (clk), .D (signal_13209), .Q (signal_13210) ) ;
    buf_clk cell_8324 ( .C (clk), .D (signal_13211), .Q (signal_13212) ) ;
    buf_clk cell_8326 ( .C (clk), .D (signal_13213), .Q (signal_13214) ) ;
    buf_clk cell_8328 ( .C (clk), .D (signal_13215), .Q (signal_13216) ) ;
    buf_clk cell_8330 ( .C (clk), .D (signal_13217), .Q (signal_13218) ) ;
    buf_clk cell_8332 ( .C (clk), .D (signal_13219), .Q (signal_13220) ) ;
    buf_clk cell_8334 ( .C (clk), .D (signal_13221), .Q (signal_13222) ) ;
    buf_clk cell_8336 ( .C (clk), .D (signal_13223), .Q (signal_13224) ) ;
    buf_clk cell_8338 ( .C (clk), .D (signal_13225), .Q (signal_13226) ) ;
    buf_clk cell_8340 ( .C (clk), .D (signal_13227), .Q (signal_13228) ) ;
    buf_clk cell_8342 ( .C (clk), .D (signal_13229), .Q (signal_13230) ) ;
    buf_clk cell_8344 ( .C (clk), .D (signal_13231), .Q (signal_13232) ) ;
    buf_clk cell_8346 ( .C (clk), .D (signal_13233), .Q (signal_13234) ) ;
    buf_clk cell_8348 ( .C (clk), .D (signal_13235), .Q (signal_13236) ) ;
    buf_clk cell_8350 ( .C (clk), .D (signal_13237), .Q (signal_13238) ) ;
    buf_clk cell_8352 ( .C (clk), .D (signal_13239), .Q (signal_13240) ) ;
    buf_clk cell_8354 ( .C (clk), .D (signal_13241), .Q (signal_13242) ) ;
    buf_clk cell_8356 ( .C (clk), .D (signal_13243), .Q (signal_13244) ) ;
    buf_clk cell_8358 ( .C (clk), .D (signal_13245), .Q (signal_13246) ) ;
    buf_clk cell_8360 ( .C (clk), .D (signal_13247), .Q (signal_13248) ) ;
    buf_clk cell_8362 ( .C (clk), .D (signal_13249), .Q (signal_13250) ) ;
    buf_clk cell_8364 ( .C (clk), .D (signal_13251), .Q (signal_13252) ) ;
    buf_clk cell_8366 ( .C (clk), .D (signal_13253), .Q (signal_13254) ) ;
    buf_clk cell_8368 ( .C (clk), .D (signal_13255), .Q (signal_13256) ) ;
    buf_clk cell_8370 ( .C (clk), .D (signal_13257), .Q (signal_13258) ) ;
    buf_clk cell_8372 ( .C (clk), .D (signal_13259), .Q (signal_13260) ) ;
    buf_clk cell_8374 ( .C (clk), .D (signal_13261), .Q (signal_13262) ) ;
    buf_clk cell_8376 ( .C (clk), .D (signal_13263), .Q (signal_13264) ) ;
    buf_clk cell_8378 ( .C (clk), .D (signal_13265), .Q (signal_13266) ) ;
    buf_clk cell_8380 ( .C (clk), .D (signal_13267), .Q (signal_13268) ) ;
    buf_clk cell_8382 ( .C (clk), .D (signal_13269), .Q (signal_13270) ) ;
    buf_clk cell_8384 ( .C (clk), .D (signal_13271), .Q (signal_13272) ) ;
    buf_clk cell_8386 ( .C (clk), .D (signal_13273), .Q (signal_13274) ) ;
    buf_clk cell_8388 ( .C (clk), .D (signal_13275), .Q (signal_13276) ) ;
    buf_clk cell_8390 ( .C (clk), .D (signal_13277), .Q (signal_13278) ) ;
    buf_clk cell_8392 ( .C (clk), .D (signal_13279), .Q (signal_13280) ) ;
    buf_clk cell_8394 ( .C (clk), .D (signal_13281), .Q (signal_13282) ) ;
    buf_clk cell_8396 ( .C (clk), .D (signal_13283), .Q (signal_13284) ) ;
    buf_clk cell_8398 ( .C (clk), .D (signal_13285), .Q (signal_13286) ) ;
    buf_clk cell_8400 ( .C (clk), .D (signal_13287), .Q (signal_13288) ) ;
    buf_clk cell_8402 ( .C (clk), .D (signal_13289), .Q (signal_13290) ) ;
    buf_clk cell_8404 ( .C (clk), .D (signal_13291), .Q (signal_13292) ) ;
    buf_clk cell_8406 ( .C (clk), .D (signal_13293), .Q (signal_13294) ) ;
    buf_clk cell_8408 ( .C (clk), .D (signal_13295), .Q (signal_13296) ) ;
    buf_clk cell_8410 ( .C (clk), .D (signal_13297), .Q (signal_13298) ) ;
    buf_clk cell_8412 ( .C (clk), .D (signal_13299), .Q (signal_13300) ) ;
    buf_clk cell_8414 ( .C (clk), .D (signal_13301), .Q (signal_13302) ) ;
    buf_clk cell_8416 ( .C (clk), .D (signal_13303), .Q (signal_13304) ) ;
    buf_clk cell_8418 ( .C (clk), .D (signal_13305), .Q (signal_13306) ) ;
    buf_clk cell_8420 ( .C (clk), .D (signal_13307), .Q (signal_13308) ) ;
    buf_clk cell_8422 ( .C (clk), .D (signal_13309), .Q (signal_13310) ) ;
    buf_clk cell_8424 ( .C (clk), .D (signal_13311), .Q (signal_13312) ) ;
    buf_clk cell_8426 ( .C (clk), .D (signal_13313), .Q (signal_13314) ) ;
    buf_clk cell_8428 ( .C (clk), .D (signal_13315), .Q (signal_13316) ) ;
    buf_clk cell_8430 ( .C (clk), .D (signal_13317), .Q (signal_13318) ) ;
    buf_clk cell_8432 ( .C (clk), .D (signal_13319), .Q (signal_13320) ) ;
    buf_clk cell_8434 ( .C (clk), .D (signal_13321), .Q (signal_13322) ) ;
    buf_clk cell_8436 ( .C (clk), .D (signal_13323), .Q (signal_13324) ) ;
    buf_clk cell_8438 ( .C (clk), .D (signal_13325), .Q (signal_13326) ) ;
    buf_clk cell_8440 ( .C (clk), .D (signal_13327), .Q (signal_13328) ) ;
    buf_clk cell_8442 ( .C (clk), .D (signal_13329), .Q (signal_13330) ) ;
    buf_clk cell_8444 ( .C (clk), .D (signal_13331), .Q (signal_13332) ) ;
    buf_clk cell_8446 ( .C (clk), .D (signal_13333), .Q (signal_13334) ) ;
    buf_clk cell_8448 ( .C (clk), .D (signal_13335), .Q (signal_13336) ) ;
    buf_clk cell_8450 ( .C (clk), .D (signal_13337), .Q (signal_13338) ) ;
    buf_clk cell_8452 ( .C (clk), .D (signal_13339), .Q (signal_13340) ) ;
    buf_clk cell_8454 ( .C (clk), .D (signal_13341), .Q (signal_13342) ) ;
    buf_clk cell_8456 ( .C (clk), .D (signal_13343), .Q (signal_13344) ) ;
    buf_clk cell_8458 ( .C (clk), .D (signal_13345), .Q (signal_13346) ) ;
    buf_clk cell_8460 ( .C (clk), .D (signal_13347), .Q (signal_13348) ) ;
    buf_clk cell_8462 ( .C (clk), .D (signal_13349), .Q (signal_13350) ) ;
    buf_clk cell_8464 ( .C (clk), .D (signal_13351), .Q (signal_13352) ) ;
    buf_clk cell_8466 ( .C (clk), .D (signal_13353), .Q (signal_13354) ) ;
    buf_clk cell_8468 ( .C (clk), .D (signal_13355), .Q (signal_13356) ) ;
    buf_clk cell_8470 ( .C (clk), .D (signal_13357), .Q (signal_13358) ) ;
    buf_clk cell_8472 ( .C (clk), .D (signal_13359), .Q (signal_13360) ) ;
    buf_clk cell_8474 ( .C (clk), .D (signal_13361), .Q (signal_13362) ) ;
    buf_clk cell_8476 ( .C (clk), .D (signal_13363), .Q (signal_13364) ) ;
    buf_clk cell_8478 ( .C (clk), .D (signal_13365), .Q (signal_13366) ) ;
    buf_clk cell_8480 ( .C (clk), .D (signal_13367), .Q (signal_13368) ) ;
    buf_clk cell_8482 ( .C (clk), .D (signal_13369), .Q (signal_13370) ) ;
    buf_clk cell_8484 ( .C (clk), .D (signal_13371), .Q (signal_13372) ) ;
    buf_clk cell_8486 ( .C (clk), .D (signal_13373), .Q (signal_13374) ) ;
    buf_clk cell_8488 ( .C (clk), .D (signal_13375), .Q (signal_13376) ) ;
    buf_clk cell_8490 ( .C (clk), .D (signal_13377), .Q (signal_13378) ) ;
    buf_clk cell_8492 ( .C (clk), .D (signal_13379), .Q (signal_13380) ) ;
    buf_clk cell_8494 ( .C (clk), .D (signal_13381), .Q (signal_13382) ) ;
    buf_clk cell_8496 ( .C (clk), .D (signal_13383), .Q (signal_13384) ) ;
    buf_clk cell_8498 ( .C (clk), .D (signal_13385), .Q (signal_13386) ) ;
    buf_clk cell_8500 ( .C (clk), .D (signal_13387), .Q (signal_13388) ) ;
    buf_clk cell_8502 ( .C (clk), .D (signal_13389), .Q (signal_13390) ) ;
    buf_clk cell_8504 ( .C (clk), .D (signal_13391), .Q (signal_13392) ) ;
    buf_clk cell_8506 ( .C (clk), .D (signal_13393), .Q (signal_13394) ) ;
    buf_clk cell_8508 ( .C (clk), .D (signal_13395), .Q (signal_13396) ) ;
    buf_clk cell_8510 ( .C (clk), .D (signal_13397), .Q (signal_13398) ) ;
    buf_clk cell_8512 ( .C (clk), .D (signal_13399), .Q (signal_13400) ) ;
    buf_clk cell_8514 ( .C (clk), .D (signal_13401), .Q (signal_13402) ) ;
    buf_clk cell_8516 ( .C (clk), .D (signal_13403), .Q (signal_13404) ) ;
    buf_clk cell_8518 ( .C (clk), .D (signal_13405), .Q (signal_13406) ) ;
    buf_clk cell_8520 ( .C (clk), .D (signal_13407), .Q (signal_13408) ) ;
    buf_clk cell_8522 ( .C (clk), .D (signal_13409), .Q (signal_13410) ) ;
    buf_clk cell_8524 ( .C (clk), .D (signal_13411), .Q (signal_13412) ) ;
    buf_clk cell_8526 ( .C (clk), .D (signal_13413), .Q (signal_13414) ) ;
    buf_clk cell_8528 ( .C (clk), .D (signal_13415), .Q (signal_13416) ) ;
    buf_clk cell_8530 ( .C (clk), .D (signal_13417), .Q (signal_13418) ) ;
    buf_clk cell_8532 ( .C (clk), .D (signal_13419), .Q (signal_13420) ) ;
    buf_clk cell_8534 ( .C (clk), .D (signal_13421), .Q (signal_13422) ) ;
    buf_clk cell_8536 ( .C (clk), .D (signal_13423), .Q (signal_13424) ) ;
    buf_clk cell_8538 ( .C (clk), .D (signal_13425), .Q (signal_13426) ) ;
    buf_clk cell_8540 ( .C (clk), .D (signal_13427), .Q (signal_13428) ) ;
    buf_clk cell_8546 ( .C (clk), .D (signal_13433), .Q (signal_13434) ) ;
    buf_clk cell_8554 ( .C (clk), .D (signal_13441), .Q (signal_13442) ) ;
    buf_clk cell_8562 ( .C (clk), .D (signal_13449), .Q (signal_13450) ) ;
    buf_clk cell_8570 ( .C (clk), .D (signal_13457), .Q (signal_13458) ) ;
    buf_clk cell_8578 ( .C (clk), .D (signal_13465), .Q (signal_13466) ) ;
    buf_clk cell_8586 ( .C (clk), .D (signal_13473), .Q (signal_13474) ) ;
    buf_clk cell_8594 ( .C (clk), .D (signal_13481), .Q (signal_13482) ) ;
    buf_clk cell_8602 ( .C (clk), .D (signal_13489), .Q (signal_13490) ) ;
    buf_clk cell_8610 ( .C (clk), .D (signal_13497), .Q (signal_13498) ) ;
    buf_clk cell_8618 ( .C (clk), .D (signal_13505), .Q (signal_13506) ) ;
    buf_clk cell_8626 ( .C (clk), .D (signal_13513), .Q (signal_13514) ) ;
    buf_clk cell_8634 ( .C (clk), .D (signal_13521), .Q (signal_13522) ) ;
    buf_clk cell_8642 ( .C (clk), .D (signal_13529), .Q (signal_13530) ) ;
    buf_clk cell_8650 ( .C (clk), .D (signal_13537), .Q (signal_13538) ) ;
    buf_clk cell_8658 ( .C (clk), .D (signal_13545), .Q (signal_13546) ) ;
    buf_clk cell_8666 ( .C (clk), .D (signal_13553), .Q (signal_13554) ) ;
    buf_clk cell_8674 ( .C (clk), .D (signal_13561), .Q (signal_13562) ) ;
    buf_clk cell_8682 ( .C (clk), .D (signal_13569), .Q (signal_13570) ) ;
    buf_clk cell_8690 ( .C (clk), .D (signal_13577), .Q (signal_13578) ) ;
    buf_clk cell_8698 ( .C (clk), .D (signal_13585), .Q (signal_13586) ) ;
    buf_clk cell_8706 ( .C (clk), .D (signal_13593), .Q (signal_13594) ) ;
    buf_clk cell_8714 ( .C (clk), .D (signal_13601), .Q (signal_13602) ) ;
    buf_clk cell_8722 ( .C (clk), .D (signal_13609), .Q (signal_13610) ) ;
    buf_clk cell_8730 ( .C (clk), .D (signal_13617), .Q (signal_13618) ) ;
    buf_clk cell_8738 ( .C (clk), .D (signal_13625), .Q (signal_13626) ) ;
    buf_clk cell_8746 ( .C (clk), .D (signal_13633), .Q (signal_13634) ) ;
    buf_clk cell_8754 ( .C (clk), .D (signal_13641), .Q (signal_13642) ) ;
    buf_clk cell_8762 ( .C (clk), .D (signal_13649), .Q (signal_13650) ) ;
    buf_clk cell_8770 ( .C (clk), .D (signal_13657), .Q (signal_13658) ) ;
    buf_clk cell_8778 ( .C (clk), .D (signal_13665), .Q (signal_13666) ) ;
    buf_clk cell_8786 ( .C (clk), .D (signal_13673), .Q (signal_13674) ) ;
    buf_clk cell_8794 ( .C (clk), .D (signal_13681), .Q (signal_13682) ) ;
    buf_clk cell_8802 ( .C (clk), .D (signal_13689), .Q (signal_13690) ) ;
    buf_clk cell_8810 ( .C (clk), .D (signal_13697), .Q (signal_13698) ) ;
    buf_clk cell_8818 ( .C (clk), .D (signal_13705), .Q (signal_13706) ) ;
    buf_clk cell_8826 ( .C (clk), .D (signal_13713), .Q (signal_13714) ) ;
    buf_clk cell_8834 ( .C (clk), .D (signal_13721), .Q (signal_13722) ) ;
    buf_clk cell_8842 ( .C (clk), .D (signal_13729), .Q (signal_13730) ) ;
    buf_clk cell_8850 ( .C (clk), .D (signal_13737), .Q (signal_13738) ) ;
    buf_clk cell_8858 ( .C (clk), .D (signal_13745), .Q (signal_13746) ) ;
    buf_clk cell_8866 ( .C (clk), .D (signal_13753), .Q (signal_13754) ) ;
    buf_clk cell_8874 ( .C (clk), .D (signal_13761), .Q (signal_13762) ) ;
    buf_clk cell_8882 ( .C (clk), .D (signal_13769), .Q (signal_13770) ) ;
    buf_clk cell_8890 ( .C (clk), .D (signal_13777), .Q (signal_13778) ) ;
    buf_clk cell_8898 ( .C (clk), .D (signal_13785), .Q (signal_13786) ) ;
    buf_clk cell_8906 ( .C (clk), .D (signal_13793), .Q (signal_13794) ) ;
    buf_clk cell_8914 ( .C (clk), .D (signal_13801), .Q (signal_13802) ) ;
    buf_clk cell_8922 ( .C (clk), .D (signal_13809), .Q (signal_13810) ) ;
    buf_clk cell_8930 ( .C (clk), .D (signal_13817), .Q (signal_13818) ) ;
    buf_clk cell_8938 ( .C (clk), .D (signal_13825), .Q (signal_13826) ) ;
    buf_clk cell_8946 ( .C (clk), .D (signal_13833), .Q (signal_13834) ) ;
    buf_clk cell_8954 ( .C (clk), .D (signal_13841), .Q (signal_13842) ) ;
    buf_clk cell_8962 ( .C (clk), .D (signal_13849), .Q (signal_13850) ) ;
    buf_clk cell_8970 ( .C (clk), .D (signal_13857), .Q (signal_13858) ) ;
    buf_clk cell_8978 ( .C (clk), .D (signal_13865), .Q (signal_13866) ) ;
    buf_clk cell_8986 ( .C (clk), .D (signal_13873), .Q (signal_13874) ) ;
    buf_clk cell_8994 ( .C (clk), .D (signal_13881), .Q (signal_13882) ) ;
    buf_clk cell_9002 ( .C (clk), .D (signal_13889), .Q (signal_13890) ) ;
    buf_clk cell_9010 ( .C (clk), .D (signal_13897), .Q (signal_13898) ) ;
    buf_clk cell_9018 ( .C (clk), .D (signal_13905), .Q (signal_13906) ) ;
    buf_clk cell_9026 ( .C (clk), .D (signal_13913), .Q (signal_13914) ) ;
    buf_clk cell_9034 ( .C (clk), .D (signal_13921), .Q (signal_13922) ) ;
    buf_clk cell_9042 ( .C (clk), .D (signal_13929), .Q (signal_13930) ) ;
    buf_clk cell_9050 ( .C (clk), .D (signal_13937), .Q (signal_13938) ) ;
    buf_clk cell_9058 ( .C (clk), .D (signal_13945), .Q (signal_13946) ) ;
    buf_clk cell_9066 ( .C (clk), .D (signal_13953), .Q (signal_13954) ) ;
    buf_clk cell_9074 ( .C (clk), .D (signal_13961), .Q (signal_13962) ) ;
    buf_clk cell_9082 ( .C (clk), .D (signal_13969), .Q (signal_13970) ) ;
    buf_clk cell_9090 ( .C (clk), .D (signal_13977), .Q (signal_13978) ) ;
    buf_clk cell_9098 ( .C (clk), .D (signal_13985), .Q (signal_13986) ) ;
    buf_clk cell_9106 ( .C (clk), .D (signal_13993), .Q (signal_13994) ) ;
    buf_clk cell_9114 ( .C (clk), .D (signal_14001), .Q (signal_14002) ) ;
    buf_clk cell_9122 ( .C (clk), .D (signal_14009), .Q (signal_14010) ) ;
    buf_clk cell_9130 ( .C (clk), .D (signal_14017), .Q (signal_14018) ) ;
    buf_clk cell_9138 ( .C (clk), .D (signal_14025), .Q (signal_14026) ) ;
    buf_clk cell_9146 ( .C (clk), .D (signal_14033), .Q (signal_14034) ) ;
    buf_clk cell_9154 ( .C (clk), .D (signal_14041), .Q (signal_14042) ) ;
    buf_clk cell_9162 ( .C (clk), .D (signal_14049), .Q (signal_14050) ) ;
    buf_clk cell_9170 ( .C (clk), .D (signal_14057), .Q (signal_14058) ) ;
    buf_clk cell_9178 ( .C (clk), .D (signal_14065), .Q (signal_14066) ) ;
    buf_clk cell_9186 ( .C (clk), .D (signal_14073), .Q (signal_14074) ) ;
    buf_clk cell_9194 ( .C (clk), .D (signal_14081), .Q (signal_14082) ) ;
    buf_clk cell_9202 ( .C (clk), .D (signal_14089), .Q (signal_14090) ) ;
    buf_clk cell_9210 ( .C (clk), .D (signal_14097), .Q (signal_14098) ) ;
    buf_clk cell_9218 ( .C (clk), .D (signal_14105), .Q (signal_14106) ) ;
    buf_clk cell_9226 ( .C (clk), .D (signal_14113), .Q (signal_14114) ) ;
    buf_clk cell_9234 ( .C (clk), .D (signal_14121), .Q (signal_14122) ) ;
    buf_clk cell_9242 ( .C (clk), .D (signal_14129), .Q (signal_14130) ) ;
    buf_clk cell_9250 ( .C (clk), .D (signal_14137), .Q (signal_14138) ) ;
    buf_clk cell_9258 ( .C (clk), .D (signal_14145), .Q (signal_14146) ) ;
    buf_clk cell_9266 ( .C (clk), .D (signal_14153), .Q (signal_14154) ) ;
    buf_clk cell_9274 ( .C (clk), .D (signal_14161), .Q (signal_14162) ) ;
    buf_clk cell_9282 ( .C (clk), .D (signal_14169), .Q (signal_14170) ) ;
    buf_clk cell_9290 ( .C (clk), .D (signal_14177), .Q (signal_14178) ) ;
    buf_clk cell_9298 ( .C (clk), .D (signal_14185), .Q (signal_14186) ) ;
    buf_clk cell_9306 ( .C (clk), .D (signal_14193), .Q (signal_14194) ) ;
    buf_clk cell_9314 ( .C (clk), .D (signal_14201), .Q (signal_14202) ) ;
    buf_clk cell_9322 ( .C (clk), .D (signal_14209), .Q (signal_14210) ) ;
    buf_clk cell_9330 ( .C (clk), .D (signal_14217), .Q (signal_14218) ) ;
    buf_clk cell_9338 ( .C (clk), .D (signal_14225), .Q (signal_14226) ) ;
    buf_clk cell_9346 ( .C (clk), .D (signal_14233), .Q (signal_14234) ) ;
    buf_clk cell_9354 ( .C (clk), .D (signal_14241), .Q (signal_14242) ) ;
    buf_clk cell_9362 ( .C (clk), .D (signal_14249), .Q (signal_14250) ) ;
    buf_clk cell_9370 ( .C (clk), .D (signal_14257), .Q (signal_14258) ) ;
    buf_clk cell_9378 ( .C (clk), .D (signal_14265), .Q (signal_14266) ) ;
    buf_clk cell_9386 ( .C (clk), .D (signal_14273), .Q (signal_14274) ) ;
    buf_clk cell_9394 ( .C (clk), .D (signal_14281), .Q (signal_14282) ) ;
    buf_clk cell_9402 ( .C (clk), .D (signal_14289), .Q (signal_14290) ) ;
    buf_clk cell_9410 ( .C (clk), .D (signal_14297), .Q (signal_14298) ) ;
    buf_clk cell_9418 ( .C (clk), .D (signal_14305), .Q (signal_14306) ) ;
    buf_clk cell_9426 ( .C (clk), .D (signal_14313), .Q (signal_14314) ) ;
    buf_clk cell_9434 ( .C (clk), .D (signal_14321), .Q (signal_14322) ) ;
    buf_clk cell_9442 ( .C (clk), .D (signal_14329), .Q (signal_14330) ) ;
    buf_clk cell_9450 ( .C (clk), .D (signal_14337), .Q (signal_14338) ) ;
    buf_clk cell_9458 ( .C (clk), .D (signal_14345), .Q (signal_14346) ) ;
    buf_clk cell_9466 ( .C (clk), .D (signal_14353), .Q (signal_14354) ) ;
    buf_clk cell_9474 ( .C (clk), .D (signal_14361), .Q (signal_14362) ) ;
    buf_clk cell_9482 ( .C (clk), .D (signal_14369), .Q (signal_14370) ) ;
    buf_clk cell_9490 ( .C (clk), .D (signal_14377), .Q (signal_14378) ) ;
    buf_clk cell_9498 ( .C (clk), .D (signal_14385), .Q (signal_14386) ) ;
    buf_clk cell_9506 ( .C (clk), .D (signal_14393), .Q (signal_14394) ) ;
    buf_clk cell_9514 ( .C (clk), .D (signal_14401), .Q (signal_14402) ) ;
    buf_clk cell_9522 ( .C (clk), .D (signal_14409), .Q (signal_14410) ) ;
    buf_clk cell_9530 ( .C (clk), .D (signal_14417), .Q (signal_14418) ) ;
    buf_clk cell_9538 ( .C (clk), .D (signal_14425), .Q (signal_14426) ) ;
    buf_clk cell_9546 ( .C (clk), .D (signal_14433), .Q (signal_14434) ) ;
    buf_clk cell_9554 ( .C (clk), .D (signal_14441), .Q (signal_14442) ) ;
    buf_clk cell_9562 ( .C (clk), .D (signal_14449), .Q (signal_14450) ) ;
    buf_clk cell_9570 ( .C (clk), .D (signal_14457), .Q (signal_14458) ) ;
    buf_clk cell_9578 ( .C (clk), .D (signal_14465), .Q (signal_14466) ) ;
    buf_clk cell_9586 ( .C (clk), .D (signal_14473), .Q (signal_14474) ) ;
    buf_clk cell_9594 ( .C (clk), .D (signal_14481), .Q (signal_14482) ) ;
    buf_clk cell_9602 ( .C (clk), .D (signal_14489), .Q (signal_14490) ) ;
    buf_clk cell_9610 ( .C (clk), .D (signal_14497), .Q (signal_14498) ) ;
    buf_clk cell_9618 ( .C (clk), .D (signal_14505), .Q (signal_14506) ) ;
    buf_clk cell_9626 ( .C (clk), .D (signal_14513), .Q (signal_14514) ) ;
    buf_clk cell_9634 ( .C (clk), .D (signal_14521), .Q (signal_14522) ) ;
    buf_clk cell_9642 ( .C (clk), .D (signal_14529), .Q (signal_14530) ) ;
    buf_clk cell_9650 ( .C (clk), .D (signal_14537), .Q (signal_14538) ) ;
    buf_clk cell_9658 ( .C (clk), .D (signal_14545), .Q (signal_14546) ) ;
    buf_clk cell_9666 ( .C (clk), .D (signal_14553), .Q (signal_14554) ) ;
    buf_clk cell_9674 ( .C (clk), .D (signal_14561), .Q (signal_14562) ) ;
    buf_clk cell_9682 ( .C (clk), .D (signal_14569), .Q (signal_14570) ) ;
    buf_clk cell_9690 ( .C (clk), .D (signal_14577), .Q (signal_14578) ) ;
    buf_clk cell_9698 ( .C (clk), .D (signal_14585), .Q (signal_14586) ) ;
    buf_clk cell_9706 ( .C (clk), .D (signal_14593), .Q (signal_14594) ) ;
    buf_clk cell_9714 ( .C (clk), .D (signal_14601), .Q (signal_14602) ) ;
    buf_clk cell_9722 ( .C (clk), .D (signal_14609), .Q (signal_14610) ) ;
    buf_clk cell_9730 ( .C (clk), .D (signal_14617), .Q (signal_14618) ) ;
    buf_clk cell_9738 ( .C (clk), .D (signal_14625), .Q (signal_14626) ) ;
    buf_clk cell_9746 ( .C (clk), .D (signal_14633), .Q (signal_14634) ) ;
    buf_clk cell_9754 ( .C (clk), .D (signal_14641), .Q (signal_14642) ) ;
    buf_clk cell_9762 ( .C (clk), .D (signal_14649), .Q (signal_14650) ) ;
    buf_clk cell_9770 ( .C (clk), .D (signal_14657), .Q (signal_14658) ) ;
    buf_clk cell_9778 ( .C (clk), .D (signal_14665), .Q (signal_14666) ) ;
    buf_clk cell_9786 ( .C (clk), .D (signal_14673), .Q (signal_14674) ) ;
    buf_clk cell_9794 ( .C (clk), .D (signal_14681), .Q (signal_14682) ) ;
    buf_clk cell_9802 ( .C (clk), .D (signal_14689), .Q (signal_14690) ) ;
    buf_clk cell_9810 ( .C (clk), .D (signal_14697), .Q (signal_14698) ) ;
    buf_clk cell_9818 ( .C (clk), .D (signal_14705), .Q (signal_14706) ) ;
    buf_clk cell_9826 ( .C (clk), .D (signal_14713), .Q (signal_14714) ) ;
    buf_clk cell_9834 ( .C (clk), .D (signal_14721), .Q (signal_14722) ) ;
    buf_clk cell_9842 ( .C (clk), .D (signal_14729), .Q (signal_14730) ) ;
    buf_clk cell_9850 ( .C (clk), .D (signal_14737), .Q (signal_14738) ) ;
    buf_clk cell_9858 ( .C (clk), .D (signal_14745), .Q (signal_14746) ) ;
    buf_clk cell_9866 ( .C (clk), .D (signal_14753), .Q (signal_14754) ) ;
    buf_clk cell_9874 ( .C (clk), .D (signal_14761), .Q (signal_14762) ) ;
    buf_clk cell_9882 ( .C (clk), .D (signal_14769), .Q (signal_14770) ) ;
    buf_clk cell_9890 ( .C (clk), .D (signal_14777), .Q (signal_14778) ) ;
    buf_clk cell_9898 ( .C (clk), .D (signal_14785), .Q (signal_14786) ) ;
    buf_clk cell_9906 ( .C (clk), .D (signal_14793), .Q (signal_14794) ) ;
    buf_clk cell_9914 ( .C (clk), .D (signal_14801), .Q (signal_14802) ) ;
    buf_clk cell_9922 ( .C (clk), .D (signal_14809), .Q (signal_14810) ) ;
    buf_clk cell_9930 ( .C (clk), .D (signal_14817), .Q (signal_14818) ) ;
    buf_clk cell_9938 ( .C (clk), .D (signal_14825), .Q (signal_14826) ) ;
    buf_clk cell_9946 ( .C (clk), .D (signal_14833), .Q (signal_14834) ) ;
    buf_clk cell_9954 ( .C (clk), .D (signal_14841), .Q (signal_14842) ) ;
    buf_clk cell_9962 ( .C (clk), .D (signal_14849), .Q (signal_14850) ) ;
    buf_clk cell_9970 ( .C (clk), .D (signal_14857), .Q (signal_14858) ) ;
    buf_clk cell_9978 ( .C (clk), .D (signal_14865), .Q (signal_14866) ) ;
    buf_clk cell_9986 ( .C (clk), .D (signal_14873), .Q (signal_14874) ) ;
    buf_clk cell_9994 ( .C (clk), .D (signal_14881), .Q (signal_14882) ) ;
    buf_clk cell_10002 ( .C (clk), .D (signal_14889), .Q (signal_14890) ) ;
    buf_clk cell_10010 ( .C (clk), .D (signal_14897), .Q (signal_14898) ) ;
    buf_clk cell_10018 ( .C (clk), .D (signal_14905), .Q (signal_14906) ) ;
    buf_clk cell_10026 ( .C (clk), .D (signal_14913), .Q (signal_14914) ) ;
    buf_clk cell_10034 ( .C (clk), .D (signal_14921), .Q (signal_14922) ) ;
    buf_clk cell_10042 ( .C (clk), .D (signal_14929), .Q (signal_14930) ) ;
    buf_clk cell_10050 ( .C (clk), .D (signal_14937), .Q (signal_14938) ) ;
    buf_clk cell_10058 ( .C (clk), .D (signal_14945), .Q (signal_14946) ) ;
    buf_clk cell_10066 ( .C (clk), .D (signal_14953), .Q (signal_14954) ) ;
    buf_clk cell_10074 ( .C (clk), .D (signal_14961), .Q (signal_14962) ) ;
    buf_clk cell_10082 ( .C (clk), .D (signal_14969), .Q (signal_14970) ) ;
    buf_clk cell_10090 ( .C (clk), .D (signal_14977), .Q (signal_14978) ) ;
    buf_clk cell_10098 ( .C (clk), .D (signal_14985), .Q (signal_14986) ) ;
    buf_clk cell_10106 ( .C (clk), .D (signal_14993), .Q (signal_14994) ) ;
    buf_clk cell_10114 ( .C (clk), .D (signal_15001), .Q (signal_15002) ) ;
    buf_clk cell_10122 ( .C (clk), .D (signal_15009), .Q (signal_15010) ) ;
    buf_clk cell_10130 ( .C (clk), .D (signal_15017), .Q (signal_15018) ) ;
    buf_clk cell_10138 ( .C (clk), .D (signal_15025), .Q (signal_15026) ) ;
    buf_clk cell_10146 ( .C (clk), .D (signal_15033), .Q (signal_15034) ) ;
    buf_clk cell_10154 ( .C (clk), .D (signal_15041), .Q (signal_15042) ) ;
    buf_clk cell_10162 ( .C (clk), .D (signal_15049), .Q (signal_15050) ) ;
    buf_clk cell_10170 ( .C (clk), .D (signal_15057), .Q (signal_15058) ) ;
    buf_clk cell_10178 ( .C (clk), .D (signal_15065), .Q (signal_15066) ) ;
    buf_clk cell_10186 ( .C (clk), .D (signal_15073), .Q (signal_15074) ) ;
    buf_clk cell_10194 ( .C (clk), .D (signal_15081), .Q (signal_15082) ) ;
    buf_clk cell_10202 ( .C (clk), .D (signal_15089), .Q (signal_15090) ) ;
    buf_clk cell_10210 ( .C (clk), .D (signal_15097), .Q (signal_15098) ) ;
    buf_clk cell_10218 ( .C (clk), .D (signal_15105), .Q (signal_15106) ) ;
    buf_clk cell_10226 ( .C (clk), .D (signal_15113), .Q (signal_15114) ) ;
    buf_clk cell_10234 ( .C (clk), .D (signal_15121), .Q (signal_15122) ) ;
    buf_clk cell_10242 ( .C (clk), .D (signal_15129), .Q (signal_15130) ) ;
    buf_clk cell_10250 ( .C (clk), .D (signal_15137), .Q (signal_15138) ) ;
    buf_clk cell_10258 ( .C (clk), .D (signal_15145), .Q (signal_15146) ) ;
    buf_clk cell_10266 ( .C (clk), .D (signal_15153), .Q (signal_15154) ) ;
    buf_clk cell_10274 ( .C (clk), .D (signal_15161), .Q (signal_15162) ) ;
    buf_clk cell_10282 ( .C (clk), .D (signal_15169), .Q (signal_15170) ) ;
    buf_clk cell_10290 ( .C (clk), .D (signal_15177), .Q (signal_15178) ) ;
    buf_clk cell_10298 ( .C (clk), .D (signal_15185), .Q (signal_15186) ) ;
    buf_clk cell_10306 ( .C (clk), .D (signal_15193), .Q (signal_15194) ) ;
    buf_clk cell_10314 ( .C (clk), .D (signal_15201), .Q (signal_15202) ) ;
    buf_clk cell_10322 ( .C (clk), .D (signal_15209), .Q (signal_15210) ) ;
    buf_clk cell_10330 ( .C (clk), .D (signal_15217), .Q (signal_15218) ) ;
    buf_clk cell_10338 ( .C (clk), .D (signal_15225), .Q (signal_15226) ) ;
    buf_clk cell_10346 ( .C (clk), .D (signal_15233), .Q (signal_15234) ) ;
    buf_clk cell_10354 ( .C (clk), .D (signal_15241), .Q (signal_15242) ) ;
    buf_clk cell_10362 ( .C (clk), .D (signal_15249), .Q (signal_15250) ) ;
    buf_clk cell_10370 ( .C (clk), .D (signal_15257), .Q (signal_15258) ) ;
    buf_clk cell_10378 ( .C (clk), .D (signal_15265), .Q (signal_15266) ) ;
    buf_clk cell_10386 ( .C (clk), .D (signal_15273), .Q (signal_15274) ) ;
    buf_clk cell_10394 ( .C (clk), .D (signal_15281), .Q (signal_15282) ) ;
    buf_clk cell_10402 ( .C (clk), .D (signal_15289), .Q (signal_15290) ) ;
    buf_clk cell_10410 ( .C (clk), .D (signal_15297), .Q (signal_15298) ) ;
    buf_clk cell_10418 ( .C (clk), .D (signal_15305), .Q (signal_15306) ) ;
    buf_clk cell_10426 ( .C (clk), .D (signal_15313), .Q (signal_15314) ) ;
    buf_clk cell_10434 ( .C (clk), .D (signal_15321), .Q (signal_15322) ) ;
    buf_clk cell_10442 ( .C (clk), .D (signal_15329), .Q (signal_15330) ) ;
    buf_clk cell_10450 ( .C (clk), .D (signal_15337), .Q (signal_15338) ) ;
    buf_clk cell_10458 ( .C (clk), .D (signal_15345), .Q (signal_15346) ) ;
    buf_clk cell_10466 ( .C (clk), .D (signal_15353), .Q (signal_15354) ) ;
    buf_clk cell_10474 ( .C (clk), .D (signal_15361), .Q (signal_15362) ) ;
    buf_clk cell_10482 ( .C (clk), .D (signal_15369), .Q (signal_15370) ) ;
    buf_clk cell_10490 ( .C (clk), .D (signal_15377), .Q (signal_15378) ) ;
    buf_clk cell_10498 ( .C (clk), .D (signal_15385), .Q (signal_15386) ) ;
    buf_clk cell_10506 ( .C (clk), .D (signal_15393), .Q (signal_15394) ) ;
    buf_clk cell_10514 ( .C (clk), .D (signal_15401), .Q (signal_15402) ) ;
    buf_clk cell_10522 ( .C (clk), .D (signal_15409), .Q (signal_15410) ) ;
    buf_clk cell_10530 ( .C (clk), .D (signal_15417), .Q (signal_15418) ) ;
    buf_clk cell_10538 ( .C (clk), .D (signal_15425), .Q (signal_15426) ) ;
    buf_clk cell_10546 ( .C (clk), .D (signal_15433), .Q (signal_15434) ) ;
    buf_clk cell_10554 ( .C (clk), .D (signal_15441), .Q (signal_15442) ) ;
    buf_clk cell_10562 ( .C (clk), .D (signal_15449), .Q (signal_15450) ) ;
    buf_clk cell_10570 ( .C (clk), .D (signal_15457), .Q (signal_15458) ) ;
    buf_clk cell_10578 ( .C (clk), .D (signal_15465), .Q (signal_15466) ) ;
    buf_clk cell_10586 ( .C (clk), .D (signal_15473), .Q (signal_15474) ) ;
    buf_clk cell_10594 ( .C (clk), .D (signal_15481), .Q (signal_15482) ) ;
    buf_clk cell_10602 ( .C (clk), .D (signal_15489), .Q (signal_15490) ) ;
    buf_clk cell_10610 ( .C (clk), .D (signal_15497), .Q (signal_15498) ) ;
    buf_clk cell_10618 ( .C (clk), .D (signal_15505), .Q (signal_15506) ) ;
    buf_clk cell_10626 ( .C (clk), .D (signal_15513), .Q (signal_15514) ) ;
    buf_clk cell_10634 ( .C (clk), .D (signal_15521), .Q (signal_15522) ) ;
    buf_clk cell_10642 ( .C (clk), .D (signal_15529), .Q (signal_15530) ) ;
    buf_clk cell_10650 ( .C (clk), .D (signal_15537), .Q (signal_15538) ) ;
    buf_clk cell_10658 ( .C (clk), .D (signal_15545), .Q (signal_15546) ) ;
    buf_clk cell_10666 ( .C (clk), .D (signal_15553), .Q (signal_15554) ) ;
    buf_clk cell_10674 ( .C (clk), .D (signal_15561), .Q (signal_15562) ) ;
    buf_clk cell_10682 ( .C (clk), .D (signal_15569), .Q (signal_15570) ) ;
    buf_clk cell_10690 ( .C (clk), .D (signal_15577), .Q (signal_15578) ) ;
    buf_clk cell_10698 ( .C (clk), .D (signal_15585), .Q (signal_15586) ) ;
    buf_clk cell_10706 ( .C (clk), .D (signal_15593), .Q (signal_15594) ) ;
    buf_clk cell_10714 ( .C (clk), .D (signal_15601), .Q (signal_15602) ) ;
    buf_clk cell_10722 ( .C (clk), .D (signal_15609), .Q (signal_15610) ) ;
    buf_clk cell_10730 ( .C (clk), .D (signal_15617), .Q (signal_15618) ) ;
    buf_clk cell_10738 ( .C (clk), .D (signal_15625), .Q (signal_15626) ) ;
    buf_clk cell_10746 ( .C (clk), .D (signal_15633), .Q (signal_15634) ) ;
    buf_clk cell_10754 ( .C (clk), .D (signal_15641), .Q (signal_15642) ) ;
    buf_clk cell_10762 ( .C (clk), .D (signal_15649), .Q (signal_15650) ) ;
    buf_clk cell_10770 ( .C (clk), .D (signal_15657), .Q (signal_15658) ) ;
    buf_clk cell_10778 ( .C (clk), .D (signal_15665), .Q (signal_15666) ) ;
    buf_clk cell_10786 ( .C (clk), .D (signal_15673), .Q (signal_15674) ) ;
    buf_clk cell_10794 ( .C (clk), .D (signal_15681), .Q (signal_15682) ) ;
    buf_clk cell_10802 ( .C (clk), .D (signal_15689), .Q (signal_15690) ) ;
    buf_clk cell_10810 ( .C (clk), .D (signal_15697), .Q (signal_15698) ) ;
    buf_clk cell_10818 ( .C (clk), .D (signal_15705), .Q (signal_15706) ) ;
    buf_clk cell_10826 ( .C (clk), .D (signal_15713), .Q (signal_15714) ) ;
    buf_clk cell_10834 ( .C (clk), .D (signal_15721), .Q (signal_15722) ) ;
    buf_clk cell_10842 ( .C (clk), .D (signal_15729), .Q (signal_15730) ) ;
    buf_clk cell_10850 ( .C (clk), .D (signal_15737), .Q (signal_15738) ) ;
    buf_clk cell_10858 ( .C (clk), .D (signal_15745), .Q (signal_15746) ) ;
    buf_clk cell_10866 ( .C (clk), .D (signal_15753), .Q (signal_15754) ) ;
    buf_clk cell_10874 ( .C (clk), .D (signal_15761), .Q (signal_15762) ) ;
    buf_clk cell_10882 ( .C (clk), .D (signal_15769), .Q (signal_15770) ) ;
    buf_clk cell_10890 ( .C (clk), .D (signal_15777), .Q (signal_15778) ) ;
    buf_clk cell_10898 ( .C (clk), .D (signal_15785), .Q (signal_15786) ) ;
    buf_clk cell_10906 ( .C (clk), .D (signal_15793), .Q (signal_15794) ) ;
    buf_clk cell_10914 ( .C (clk), .D (signal_15801), .Q (signal_15802) ) ;
    buf_clk cell_10922 ( .C (clk), .D (signal_15809), .Q (signal_15810) ) ;
    buf_clk cell_10930 ( .C (clk), .D (signal_15817), .Q (signal_15818) ) ;
    buf_clk cell_10938 ( .C (clk), .D (signal_15825), .Q (signal_15826) ) ;
    buf_clk cell_10946 ( .C (clk), .D (signal_15833), .Q (signal_15834) ) ;
    buf_clk cell_10954 ( .C (clk), .D (signal_15841), .Q (signal_15842) ) ;
    buf_clk cell_10962 ( .C (clk), .D (signal_15849), .Q (signal_15850) ) ;
    buf_clk cell_10970 ( .C (clk), .D (signal_15857), .Q (signal_15858) ) ;
    buf_clk cell_10978 ( .C (clk), .D (signal_15865), .Q (signal_15866) ) ;
    buf_clk cell_10986 ( .C (clk), .D (signal_15873), .Q (signal_15874) ) ;
    buf_clk cell_10994 ( .C (clk), .D (signal_15881), .Q (signal_15882) ) ;
    buf_clk cell_11002 ( .C (clk), .D (signal_15889), .Q (signal_15890) ) ;
    buf_clk cell_11010 ( .C (clk), .D (signal_15897), .Q (signal_15898) ) ;
    buf_clk cell_11018 ( .C (clk), .D (signal_15905), .Q (signal_15906) ) ;
    buf_clk cell_11026 ( .C (clk), .D (signal_15913), .Q (signal_15914) ) ;
    buf_clk cell_11034 ( .C (clk), .D (signal_15921), .Q (signal_15922) ) ;
    buf_clk cell_11042 ( .C (clk), .D (signal_15929), .Q (signal_15930) ) ;
    buf_clk cell_11050 ( .C (clk), .D (signal_15937), .Q (signal_15938) ) ;
    buf_clk cell_11058 ( .C (clk), .D (signal_15945), .Q (signal_15946) ) ;
    buf_clk cell_11066 ( .C (clk), .D (signal_15953), .Q (signal_15954) ) ;
    buf_clk cell_11074 ( .C (clk), .D (signal_15961), .Q (signal_15962) ) ;
    buf_clk cell_11082 ( .C (clk), .D (signal_15969), .Q (signal_15970) ) ;
    buf_clk cell_11090 ( .C (clk), .D (signal_15977), .Q (signal_15978) ) ;
    buf_clk cell_11098 ( .C (clk), .D (signal_15985), .Q (signal_15986) ) ;
    buf_clk cell_11106 ( .C (clk), .D (signal_15993), .Q (signal_15994) ) ;
    buf_clk cell_11114 ( .C (clk), .D (signal_16001), .Q (signal_16002) ) ;
    buf_clk cell_11122 ( .C (clk), .D (signal_16009), .Q (signal_16010) ) ;
    buf_clk cell_11130 ( .C (clk), .D (signal_16017), .Q (signal_16018) ) ;
    buf_clk cell_11138 ( .C (clk), .D (signal_16025), .Q (signal_16026) ) ;
    buf_clk cell_11146 ( .C (clk), .D (signal_16033), .Q (signal_16034) ) ;
    buf_clk cell_11154 ( .C (clk), .D (signal_16041), .Q (signal_16042) ) ;
    buf_clk cell_11162 ( .C (clk), .D (signal_16049), .Q (signal_16050) ) ;
    buf_clk cell_11170 ( .C (clk), .D (signal_16057), .Q (signal_16058) ) ;
    buf_clk cell_11178 ( .C (clk), .D (signal_16065), .Q (signal_16066) ) ;
    buf_clk cell_11186 ( .C (clk), .D (signal_16073), .Q (signal_16074) ) ;
    buf_clk cell_11194 ( .C (clk), .D (signal_16081), .Q (signal_16082) ) ;
    buf_clk cell_11202 ( .C (clk), .D (signal_16089), .Q (signal_16090) ) ;
    buf_clk cell_11210 ( .C (clk), .D (signal_16097), .Q (signal_16098) ) ;
    buf_clk cell_11218 ( .C (clk), .D (signal_16105), .Q (signal_16106) ) ;
    buf_clk cell_11226 ( .C (clk), .D (signal_16113), .Q (signal_16114) ) ;
    buf_clk cell_11234 ( .C (clk), .D (signal_16121), .Q (signal_16122) ) ;
    buf_clk cell_11242 ( .C (clk), .D (signal_16129), .Q (signal_16130) ) ;
    buf_clk cell_11250 ( .C (clk), .D (signal_16137), .Q (signal_16138) ) ;
    buf_clk cell_11258 ( .C (clk), .D (signal_16145), .Q (signal_16146) ) ;
    buf_clk cell_11266 ( .C (clk), .D (signal_16153), .Q (signal_16154) ) ;
    buf_clk cell_11274 ( .C (clk), .D (signal_16161), .Q (signal_16162) ) ;
    buf_clk cell_11282 ( .C (clk), .D (signal_16169), .Q (signal_16170) ) ;
    buf_clk cell_11290 ( .C (clk), .D (signal_16177), .Q (signal_16178) ) ;
    buf_clk cell_11298 ( .C (clk), .D (signal_16185), .Q (signal_16186) ) ;
    buf_clk cell_11306 ( .C (clk), .D (signal_16193), .Q (signal_16194) ) ;
    buf_clk cell_11314 ( .C (clk), .D (signal_16201), .Q (signal_16202) ) ;
    buf_clk cell_11322 ( .C (clk), .D (signal_16209), .Q (signal_16210) ) ;
    buf_clk cell_11330 ( .C (clk), .D (signal_16217), .Q (signal_16218) ) ;
    buf_clk cell_11338 ( .C (clk), .D (signal_16225), .Q (signal_16226) ) ;
    buf_clk cell_11346 ( .C (clk), .D (signal_16233), .Q (signal_16234) ) ;
    buf_clk cell_11354 ( .C (clk), .D (signal_16241), .Q (signal_16242) ) ;
    buf_clk cell_11362 ( .C (clk), .D (signal_16249), .Q (signal_16250) ) ;
    buf_clk cell_11370 ( .C (clk), .D (signal_16257), .Q (signal_16258) ) ;
    buf_clk cell_11378 ( .C (clk), .D (signal_16265), .Q (signal_16266) ) ;
    buf_clk cell_11386 ( .C (clk), .D (signal_16273), .Q (signal_16274) ) ;
    buf_clk cell_11394 ( .C (clk), .D (signal_16281), .Q (signal_16282) ) ;
    buf_clk cell_11402 ( .C (clk), .D (signal_16289), .Q (signal_16290) ) ;
    buf_clk cell_11410 ( .C (clk), .D (signal_16297), .Q (signal_16298) ) ;
    buf_clk cell_11418 ( .C (clk), .D (signal_16305), .Q (signal_16306) ) ;
    buf_clk cell_11426 ( .C (clk), .D (signal_16313), .Q (signal_16314) ) ;
    buf_clk cell_11434 ( .C (clk), .D (signal_16321), .Q (signal_16322) ) ;
    buf_clk cell_11442 ( .C (clk), .D (signal_16329), .Q (signal_16330) ) ;
    buf_clk cell_11450 ( .C (clk), .D (signal_16337), .Q (signal_16338) ) ;
    buf_clk cell_11458 ( .C (clk), .D (signal_16345), .Q (signal_16346) ) ;
    buf_clk cell_11466 ( .C (clk), .D (signal_16353), .Q (signal_16354) ) ;
    buf_clk cell_11474 ( .C (clk), .D (signal_16361), .Q (signal_16362) ) ;
    buf_clk cell_11482 ( .C (clk), .D (signal_16369), .Q (signal_16370) ) ;
    buf_clk cell_11490 ( .C (clk), .D (signal_16377), .Q (signal_16378) ) ;
    buf_clk cell_11498 ( .C (clk), .D (signal_16385), .Q (signal_16386) ) ;
    buf_clk cell_11506 ( .C (clk), .D (signal_16393), .Q (signal_16394) ) ;
    buf_clk cell_11514 ( .C (clk), .D (signal_16401), .Q (signal_16402) ) ;
    buf_clk cell_11522 ( .C (clk), .D (signal_16409), .Q (signal_16410) ) ;
    buf_clk cell_11530 ( .C (clk), .D (signal_16417), .Q (signal_16418) ) ;
    buf_clk cell_11538 ( .C (clk), .D (signal_16425), .Q (signal_16426) ) ;
    buf_clk cell_11546 ( .C (clk), .D (signal_16433), .Q (signal_16434) ) ;
    buf_clk cell_11554 ( .C (clk), .D (signal_16441), .Q (signal_16442) ) ;
    buf_clk cell_11562 ( .C (clk), .D (signal_16449), .Q (signal_16450) ) ;
    buf_clk cell_11570 ( .C (clk), .D (signal_16457), .Q (signal_16458) ) ;
    buf_clk cell_11578 ( .C (clk), .D (signal_16465), .Q (signal_16466) ) ;
    buf_clk cell_11586 ( .C (clk), .D (signal_16473), .Q (signal_16474) ) ;
    buf_clk cell_11594 ( .C (clk), .D (signal_16481), .Q (signal_16482) ) ;
    buf_clk cell_11602 ( .C (clk), .D (signal_16489), .Q (signal_16490) ) ;
    buf_clk cell_11610 ( .C (clk), .D (signal_16497), .Q (signal_16498) ) ;
    buf_clk cell_11618 ( .C (clk), .D (signal_16505), .Q (signal_16506) ) ;
    buf_clk cell_11626 ( .C (clk), .D (signal_16513), .Q (signal_16514) ) ;
    buf_clk cell_11634 ( .C (clk), .D (signal_16521), .Q (signal_16522) ) ;
    buf_clk cell_11642 ( .C (clk), .D (signal_16529), .Q (signal_16530) ) ;
    buf_clk cell_11650 ( .C (clk), .D (signal_16537), .Q (signal_16538) ) ;
    buf_clk cell_11658 ( .C (clk), .D (signal_16545), .Q (signal_16546) ) ;
    buf_clk cell_11666 ( .C (clk), .D (signal_16553), .Q (signal_16554) ) ;
    buf_clk cell_11674 ( .C (clk), .D (signal_16561), .Q (signal_16562) ) ;
    buf_clk cell_11682 ( .C (clk), .D (signal_16569), .Q (signal_16570) ) ;
    buf_clk cell_11690 ( .C (clk), .D (signal_16577), .Q (signal_16578) ) ;
    buf_clk cell_11698 ( .C (clk), .D (signal_16585), .Q (signal_16586) ) ;
    buf_clk cell_11706 ( .C (clk), .D (signal_16593), .Q (signal_16594) ) ;
    buf_clk cell_11714 ( .C (clk), .D (signal_16601), .Q (signal_16602) ) ;
    buf_clk cell_11722 ( .C (clk), .D (signal_16609), .Q (signal_16610) ) ;
    buf_clk cell_11730 ( .C (clk), .D (signal_16617), .Q (signal_16618) ) ;
    buf_clk cell_11738 ( .C (clk), .D (signal_16625), .Q (signal_16626) ) ;
    buf_clk cell_11746 ( .C (clk), .D (signal_16633), .Q (signal_16634) ) ;
    buf_clk cell_11754 ( .C (clk), .D (signal_16641), .Q (signal_16642) ) ;
    buf_clk cell_11762 ( .C (clk), .D (signal_16649), .Q (signal_16650) ) ;
    buf_clk cell_11770 ( .C (clk), .D (signal_16657), .Q (signal_16658) ) ;
    buf_clk cell_11778 ( .C (clk), .D (signal_16665), .Q (signal_16666) ) ;
    buf_clk cell_11786 ( .C (clk), .D (signal_16673), .Q (signal_16674) ) ;
    buf_clk cell_11794 ( .C (clk), .D (signal_16681), .Q (signal_16682) ) ;
    buf_clk cell_11802 ( .C (clk), .D (signal_16689), .Q (signal_16690) ) ;
    buf_clk cell_11810 ( .C (clk), .D (signal_16697), .Q (signal_16698) ) ;
    buf_clk cell_11818 ( .C (clk), .D (signal_16705), .Q (signal_16706) ) ;
    buf_clk cell_11826 ( .C (clk), .D (signal_16713), .Q (signal_16714) ) ;
    buf_clk cell_11834 ( .C (clk), .D (signal_16721), .Q (signal_16722) ) ;
    buf_clk cell_11842 ( .C (clk), .D (signal_16729), .Q (signal_16730) ) ;
    buf_clk cell_11850 ( .C (clk), .D (signal_16737), .Q (signal_16738) ) ;
    buf_clk cell_11858 ( .C (clk), .D (signal_16745), .Q (signal_16746) ) ;
    buf_clk cell_11866 ( .C (clk), .D (signal_16753), .Q (signal_16754) ) ;
    buf_clk cell_11874 ( .C (clk), .D (signal_16761), .Q (signal_16762) ) ;
    buf_clk cell_11882 ( .C (clk), .D (signal_16769), .Q (signal_16770) ) ;
    buf_clk cell_11890 ( .C (clk), .D (signal_16777), .Q (signal_16778) ) ;
    buf_clk cell_11898 ( .C (clk), .D (signal_16785), .Q (signal_16786) ) ;
    buf_clk cell_11906 ( .C (clk), .D (signal_16793), .Q (signal_16794) ) ;
    buf_clk cell_11914 ( .C (clk), .D (signal_16801), .Q (signal_16802) ) ;
    buf_clk cell_11922 ( .C (clk), .D (signal_16809), .Q (signal_16810) ) ;
    buf_clk cell_11930 ( .C (clk), .D (signal_16817), .Q (signal_16818) ) ;
    buf_clk cell_11938 ( .C (clk), .D (signal_16825), .Q (signal_16826) ) ;
    buf_clk cell_11946 ( .C (clk), .D (signal_16833), .Q (signal_16834) ) ;
    buf_clk cell_11954 ( .C (clk), .D (signal_16841), .Q (signal_16842) ) ;
    buf_clk cell_11962 ( .C (clk), .D (signal_16849), .Q (signal_16850) ) ;
    buf_clk cell_11970 ( .C (clk), .D (signal_16857), .Q (signal_16858) ) ;
    buf_clk cell_11978 ( .C (clk), .D (signal_16865), .Q (signal_16866) ) ;
    buf_clk cell_11986 ( .C (clk), .D (signal_16873), .Q (signal_16874) ) ;
    buf_clk cell_11994 ( .C (clk), .D (signal_16881), .Q (signal_16882) ) ;
    buf_clk cell_12002 ( .C (clk), .D (signal_16889), .Q (signal_16890) ) ;
    buf_clk cell_12010 ( .C (clk), .D (signal_16897), .Q (signal_16898) ) ;
    buf_clk cell_12018 ( .C (clk), .D (signal_16905), .Q (signal_16906) ) ;
    buf_clk cell_12026 ( .C (clk), .D (signal_16913), .Q (signal_16914) ) ;
    buf_clk cell_12034 ( .C (clk), .D (signal_16921), .Q (signal_16922) ) ;
    buf_clk cell_12042 ( .C (clk), .D (signal_16929), .Q (signal_16930) ) ;
    buf_clk cell_12050 ( .C (clk), .D (signal_16937), .Q (signal_16938) ) ;
    buf_clk cell_12058 ( .C (clk), .D (signal_16945), .Q (signal_16946) ) ;
    buf_clk cell_12066 ( .C (clk), .D (signal_16953), .Q (signal_16954) ) ;
    buf_clk cell_12074 ( .C (clk), .D (signal_16961), .Q (signal_16962) ) ;
    buf_clk cell_12082 ( .C (clk), .D (signal_16969), .Q (signal_16970) ) ;
    buf_clk cell_12090 ( .C (clk), .D (signal_16977), .Q (signal_16978) ) ;
    buf_clk cell_12098 ( .C (clk), .D (signal_16985), .Q (signal_16986) ) ;
    buf_clk cell_12106 ( .C (clk), .D (signal_16993), .Q (signal_16994) ) ;
    buf_clk cell_12114 ( .C (clk), .D (signal_17001), .Q (signal_17002) ) ;
    buf_clk cell_12122 ( .C (clk), .D (signal_17009), .Q (signal_17010) ) ;
    buf_clk cell_12130 ( .C (clk), .D (signal_17017), .Q (signal_17018) ) ;
    buf_clk cell_12138 ( .C (clk), .D (signal_17025), .Q (signal_17026) ) ;
    buf_clk cell_12146 ( .C (clk), .D (signal_17033), .Q (signal_17034) ) ;
    buf_clk cell_12154 ( .C (clk), .D (signal_17041), .Q (signal_17042) ) ;
    buf_clk cell_12162 ( .C (clk), .D (signal_17049), .Q (signal_17050) ) ;
    buf_clk cell_12170 ( .C (clk), .D (signal_17057), .Q (signal_17058) ) ;
    buf_clk cell_12178 ( .C (clk), .D (signal_17065), .Q (signal_17066) ) ;
    buf_clk cell_12186 ( .C (clk), .D (signal_17073), .Q (signal_17074) ) ;
    buf_clk cell_12194 ( .C (clk), .D (signal_17081), .Q (signal_17082) ) ;
    buf_clk cell_12202 ( .C (clk), .D (signal_17089), .Q (signal_17090) ) ;
    buf_clk cell_12210 ( .C (clk), .D (signal_17097), .Q (signal_17098) ) ;
    buf_clk cell_12218 ( .C (clk), .D (signal_17105), .Q (signal_17106) ) ;
    buf_clk cell_12226 ( .C (clk), .D (signal_17113), .Q (signal_17114) ) ;
    buf_clk cell_12234 ( .C (clk), .D (signal_17121), .Q (signal_17122) ) ;
    buf_clk cell_12242 ( .C (clk), .D (signal_17129), .Q (signal_17130) ) ;
    buf_clk cell_12250 ( .C (clk), .D (signal_17137), .Q (signal_17138) ) ;
    buf_clk cell_12258 ( .C (clk), .D (signal_17145), .Q (signal_17146) ) ;
    buf_clk cell_12266 ( .C (clk), .D (signal_17153), .Q (signal_17154) ) ;
    buf_clk cell_12274 ( .C (clk), .D (signal_17161), .Q (signal_17162) ) ;
    buf_clk cell_12282 ( .C (clk), .D (signal_17169), .Q (signal_17170) ) ;
    buf_clk cell_12290 ( .C (clk), .D (signal_17177), .Q (signal_17178) ) ;
    buf_clk cell_12298 ( .C (clk), .D (signal_17185), .Q (signal_17186) ) ;
    buf_clk cell_12306 ( .C (clk), .D (signal_17193), .Q (signal_17194) ) ;
    buf_clk cell_12314 ( .C (clk), .D (signal_17201), .Q (signal_17202) ) ;
    buf_clk cell_12322 ( .C (clk), .D (signal_17209), .Q (signal_17210) ) ;
    buf_clk cell_12330 ( .C (clk), .D (signal_17217), .Q (signal_17218) ) ;
    buf_clk cell_12338 ( .C (clk), .D (signal_17225), .Q (signal_17226) ) ;
    buf_clk cell_12346 ( .C (clk), .D (signal_17233), .Q (signal_17234) ) ;
    buf_clk cell_12354 ( .C (clk), .D (signal_17241), .Q (signal_17242) ) ;
    buf_clk cell_12362 ( .C (clk), .D (signal_17249), .Q (signal_17250) ) ;
    buf_clk cell_12370 ( .C (clk), .D (signal_17257), .Q (signal_17258) ) ;
    buf_clk cell_12378 ( .C (clk), .D (signal_17265), .Q (signal_17266) ) ;
    buf_clk cell_12386 ( .C (clk), .D (signal_17273), .Q (signal_17274) ) ;
    buf_clk cell_12394 ( .C (clk), .D (signal_17281), .Q (signal_17282) ) ;
    buf_clk cell_12402 ( .C (clk), .D (signal_17289), .Q (signal_17290) ) ;
    buf_clk cell_12410 ( .C (clk), .D (signal_17297), .Q (signal_17298) ) ;
    buf_clk cell_12418 ( .C (clk), .D (signal_17305), .Q (signal_17306) ) ;
    buf_clk cell_12426 ( .C (clk), .D (signal_17313), .Q (signal_17314) ) ;
    buf_clk cell_12434 ( .C (clk), .D (signal_17321), .Q (signal_17322) ) ;
    buf_clk cell_12442 ( .C (clk), .D (signal_17329), .Q (signal_17330) ) ;
    buf_clk cell_12450 ( .C (clk), .D (signal_17337), .Q (signal_17338) ) ;
    buf_clk cell_12458 ( .C (clk), .D (signal_17345), .Q (signal_17346) ) ;
    buf_clk cell_12466 ( .C (clk), .D (signal_17353), .Q (signal_17354) ) ;
    buf_clk cell_12474 ( .C (clk), .D (signal_17361), .Q (signal_17362) ) ;
    buf_clk cell_12482 ( .C (clk), .D (signal_17369), .Q (signal_17370) ) ;
    buf_clk cell_12490 ( .C (clk), .D (signal_17377), .Q (signal_17378) ) ;
    buf_clk cell_12498 ( .C (clk), .D (signal_17385), .Q (signal_17386) ) ;
    buf_clk cell_12506 ( .C (clk), .D (signal_17393), .Q (signal_17394) ) ;
    buf_clk cell_12514 ( .C (clk), .D (signal_17401), .Q (signal_17402) ) ;
    buf_clk cell_12522 ( .C (clk), .D (signal_17409), .Q (signal_17410) ) ;
    buf_clk cell_12530 ( .C (clk), .D (signal_17417), .Q (signal_17418) ) ;
    buf_clk cell_12538 ( .C (clk), .D (signal_17425), .Q (signal_17426) ) ;
    buf_clk cell_12546 ( .C (clk), .D (signal_17433), .Q (signal_17434) ) ;
    buf_clk cell_12554 ( .C (clk), .D (signal_17441), .Q (signal_17442) ) ;
    buf_clk cell_12562 ( .C (clk), .D (signal_17449), .Q (signal_17450) ) ;
    buf_clk cell_12570 ( .C (clk), .D (signal_17457), .Q (signal_17458) ) ;
    buf_clk cell_12578 ( .C (clk), .D (signal_17465), .Q (signal_17466) ) ;
    buf_clk cell_12586 ( .C (clk), .D (signal_17473), .Q (signal_17474) ) ;
    buf_clk cell_12594 ( .C (clk), .D (signal_17481), .Q (signal_17482) ) ;
    buf_clk cell_12602 ( .C (clk), .D (signal_17489), .Q (signal_17490) ) ;
    buf_clk cell_12610 ( .C (clk), .D (signal_17497), .Q (signal_17498) ) ;
    buf_clk cell_12618 ( .C (clk), .D (signal_17505), .Q (signal_17506) ) ;
    buf_clk cell_12626 ( .C (clk), .D (signal_17513), .Q (signal_17514) ) ;
    buf_clk cell_12634 ( .C (clk), .D (signal_17521), .Q (signal_17522) ) ;
    buf_clk cell_12642 ( .C (clk), .D (signal_17529), .Q (signal_17530) ) ;
    buf_clk cell_12650 ( .C (clk), .D (signal_17537), .Q (signal_17538) ) ;
    buf_clk cell_12658 ( .C (clk), .D (signal_17545), .Q (signal_17546) ) ;
    buf_clk cell_12666 ( .C (clk), .D (signal_17553), .Q (signal_17554) ) ;
    buf_clk cell_12674 ( .C (clk), .D (signal_17561), .Q (signal_17562) ) ;
    buf_clk cell_12682 ( .C (clk), .D (signal_17569), .Q (signal_17570) ) ;
    buf_clk cell_12690 ( .C (clk), .D (signal_17577), .Q (signal_17578) ) ;
    buf_clk cell_12698 ( .C (clk), .D (signal_17585), .Q (signal_17586) ) ;
    buf_clk cell_12706 ( .C (clk), .D (signal_17593), .Q (signal_17594) ) ;
    buf_clk cell_12714 ( .C (clk), .D (signal_17601), .Q (signal_17602) ) ;
    buf_clk cell_12722 ( .C (clk), .D (signal_17609), .Q (signal_17610) ) ;
    buf_clk cell_12730 ( .C (clk), .D (signal_17617), .Q (signal_17618) ) ;
    buf_clk cell_12738 ( .C (clk), .D (signal_17625), .Q (signal_17626) ) ;
    buf_clk cell_12746 ( .C (clk), .D (signal_17633), .Q (signal_17634) ) ;
    buf_clk cell_12754 ( .C (clk), .D (signal_17641), .Q (signal_17642) ) ;
    buf_clk cell_12762 ( .C (clk), .D (signal_17649), .Q (signal_17650) ) ;
    buf_clk cell_12770 ( .C (clk), .D (signal_17657), .Q (signal_17658) ) ;
    buf_clk cell_12778 ( .C (clk), .D (signal_17665), .Q (signal_17666) ) ;
    buf_clk cell_12786 ( .C (clk), .D (signal_17673), .Q (signal_17674) ) ;
    buf_clk cell_12794 ( .C (clk), .D (signal_17681), .Q (signal_17682) ) ;
    buf_clk cell_12802 ( .C (clk), .D (signal_17689), .Q (signal_17690) ) ;
    buf_clk cell_12810 ( .C (clk), .D (signal_17697), .Q (signal_17698) ) ;
    buf_clk cell_12818 ( .C (clk), .D (signal_17705), .Q (signal_17706) ) ;
    buf_clk cell_12826 ( .C (clk), .D (signal_17713), .Q (signal_17714) ) ;
    buf_clk cell_12834 ( .C (clk), .D (signal_17721), .Q (signal_17722) ) ;
    buf_clk cell_12842 ( .C (clk), .D (signal_17729), .Q (signal_17730) ) ;
    buf_clk cell_12850 ( .C (clk), .D (signal_17737), .Q (signal_17738) ) ;
    buf_clk cell_12858 ( .C (clk), .D (signal_17745), .Q (signal_17746) ) ;
    buf_clk cell_12866 ( .C (clk), .D (signal_17753), .Q (signal_17754) ) ;
    buf_clk cell_12874 ( .C (clk), .D (signal_17761), .Q (signal_17762) ) ;
    buf_clk cell_12882 ( .C (clk), .D (signal_17769), .Q (signal_17770) ) ;
    buf_clk cell_12890 ( .C (clk), .D (signal_17777), .Q (signal_17778) ) ;
    buf_clk cell_12898 ( .C (clk), .D (signal_17785), .Q (signal_17786) ) ;
    buf_clk cell_12906 ( .C (clk), .D (signal_17793), .Q (signal_17794) ) ;
    buf_clk cell_12914 ( .C (clk), .D (signal_17801), .Q (signal_17802) ) ;
    buf_clk cell_12922 ( .C (clk), .D (signal_17809), .Q (signal_17810) ) ;
    buf_clk cell_12930 ( .C (clk), .D (signal_17817), .Q (signal_17818) ) ;
    buf_clk cell_12938 ( .C (clk), .D (signal_17825), .Q (signal_17826) ) ;
    buf_clk cell_12946 ( .C (clk), .D (signal_17833), .Q (signal_17834) ) ;
    buf_clk cell_12954 ( .C (clk), .D (signal_17841), .Q (signal_17842) ) ;
    buf_clk cell_12962 ( .C (clk), .D (signal_17849), .Q (signal_17850) ) ;
    buf_clk cell_12970 ( .C (clk), .D (signal_17857), .Q (signal_17858) ) ;
    buf_clk cell_12978 ( .C (clk), .D (signal_17865), .Q (signal_17866) ) ;
    buf_clk cell_12986 ( .C (clk), .D (signal_17873), .Q (signal_17874) ) ;
    buf_clk cell_12994 ( .C (clk), .D (signal_17881), .Q (signal_17882) ) ;
    buf_clk cell_13002 ( .C (clk), .D (signal_17889), .Q (signal_17890) ) ;
    buf_clk cell_13010 ( .C (clk), .D (signal_17897), .Q (signal_17898) ) ;
    buf_clk cell_13018 ( .C (clk), .D (signal_17905), .Q (signal_17906) ) ;
    buf_clk cell_13026 ( .C (clk), .D (signal_17913), .Q (signal_17914) ) ;
    buf_clk cell_13034 ( .C (clk), .D (signal_17921), .Q (signal_17922) ) ;
    buf_clk cell_13042 ( .C (clk), .D (signal_17929), .Q (signal_17930) ) ;
    buf_clk cell_13050 ( .C (clk), .D (signal_17937), .Q (signal_17938) ) ;
    buf_clk cell_13058 ( .C (clk), .D (signal_17945), .Q (signal_17946) ) ;
    buf_clk cell_13066 ( .C (clk), .D (signal_17953), .Q (signal_17954) ) ;
    buf_clk cell_13074 ( .C (clk), .D (signal_17961), .Q (signal_17962) ) ;
    buf_clk cell_13082 ( .C (clk), .D (signal_17969), .Q (signal_17970) ) ;
    buf_clk cell_13090 ( .C (clk), .D (signal_17977), .Q (signal_17978) ) ;
    buf_clk cell_13098 ( .C (clk), .D (signal_17985), .Q (signal_17986) ) ;
    buf_clk cell_13106 ( .C (clk), .D (signal_17993), .Q (signal_17994) ) ;
    buf_clk cell_13114 ( .C (clk), .D (signal_18001), .Q (signal_18002) ) ;
    buf_clk cell_13122 ( .C (clk), .D (signal_18009), .Q (signal_18010) ) ;
    buf_clk cell_13130 ( .C (clk), .D (signal_18017), .Q (signal_18018) ) ;
    buf_clk cell_13138 ( .C (clk), .D (signal_18025), .Q (signal_18026) ) ;
    buf_clk cell_13146 ( .C (clk), .D (signal_18033), .Q (signal_18034) ) ;
    buf_clk cell_13154 ( .C (clk), .D (signal_18041), .Q (signal_18042) ) ;
    buf_clk cell_13162 ( .C (clk), .D (signal_18049), .Q (signal_18050) ) ;
    buf_clk cell_13170 ( .C (clk), .D (signal_18057), .Q (signal_18058) ) ;
    buf_clk cell_13178 ( .C (clk), .D (signal_18065), .Q (signal_18066) ) ;
    buf_clk cell_13186 ( .C (clk), .D (signal_18073), .Q (signal_18074) ) ;
    buf_clk cell_13194 ( .C (clk), .D (signal_18081), .Q (signal_18082) ) ;
    buf_clk cell_13202 ( .C (clk), .D (signal_18089), .Q (signal_18090) ) ;
    buf_clk cell_13210 ( .C (clk), .D (signal_18097), .Q (signal_18098) ) ;
    buf_clk cell_13218 ( .C (clk), .D (signal_18105), .Q (signal_18106) ) ;
    buf_clk cell_13226 ( .C (clk), .D (signal_18113), .Q (signal_18114) ) ;
    buf_clk cell_13234 ( .C (clk), .D (signal_18121), .Q (signal_18122) ) ;
    buf_clk cell_13242 ( .C (clk), .D (signal_18129), .Q (signal_18130) ) ;
    buf_clk cell_13250 ( .C (clk), .D (signal_18137), .Q (signal_18138) ) ;
    buf_clk cell_13258 ( .C (clk), .D (signal_18145), .Q (signal_18146) ) ;
    buf_clk cell_13266 ( .C (clk), .D (signal_18153), .Q (signal_18154) ) ;
    buf_clk cell_13274 ( .C (clk), .D (signal_18161), .Q (signal_18162) ) ;
    buf_clk cell_13282 ( .C (clk), .D (signal_18169), .Q (signal_18170) ) ;
    buf_clk cell_13288 ( .C (clk), .D (signal_18175), .Q (signal_18176) ) ;
    buf_clk cell_13294 ( .C (clk), .D (signal_18181), .Q (signal_18182) ) ;
    buf_clk cell_13300 ( .C (clk), .D (signal_18187), .Q (signal_18188) ) ;
    buf_clk cell_13306 ( .C (clk), .D (signal_18193), .Q (signal_18194) ) ;
    buf_clk cell_13312 ( .C (clk), .D (signal_18199), .Q (signal_18200) ) ;
    buf_clk cell_13318 ( .C (clk), .D (signal_18205), .Q (signal_18206) ) ;
    buf_clk cell_13324 ( .C (clk), .D (signal_18211), .Q (signal_18212) ) ;
    buf_clk cell_13330 ( .C (clk), .D (signal_18217), .Q (signal_18218) ) ;
    buf_clk cell_13336 ( .C (clk), .D (signal_18223), .Q (signal_18224) ) ;
    buf_clk cell_13342 ( .C (clk), .D (signal_18229), .Q (signal_18230) ) ;
    buf_clk cell_13348 ( .C (clk), .D (signal_18235), .Q (signal_18236) ) ;
    buf_clk cell_13354 ( .C (clk), .D (signal_18241), .Q (signal_18242) ) ;
    buf_clk cell_13360 ( .C (clk), .D (signal_18247), .Q (signal_18248) ) ;
    buf_clk cell_13366 ( .C (clk), .D (signal_18253), .Q (signal_18254) ) ;
    buf_clk cell_13372 ( .C (clk), .D (signal_18259), .Q (signal_18260) ) ;
    buf_clk cell_13378 ( .C (clk), .D (signal_18265), .Q (signal_18266) ) ;
    buf_clk cell_13384 ( .C (clk), .D (signal_18271), .Q (signal_18272) ) ;
    buf_clk cell_13390 ( .C (clk), .D (signal_18277), .Q (signal_18278) ) ;
    buf_clk cell_13396 ( .C (clk), .D (signal_18283), .Q (signal_18284) ) ;
    buf_clk cell_13402 ( .C (clk), .D (signal_18289), .Q (signal_18290) ) ;
    buf_clk cell_13408 ( .C (clk), .D (signal_18295), .Q (signal_18296) ) ;
    buf_clk cell_13414 ( .C (clk), .D (signal_18301), .Q (signal_18302) ) ;
    buf_clk cell_13420 ( .C (clk), .D (signal_18307), .Q (signal_18308) ) ;
    buf_clk cell_13426 ( .C (clk), .D (signal_18313), .Q (signal_18314) ) ;
    buf_clk cell_13432 ( .C (clk), .D (signal_18319), .Q (signal_18320) ) ;
    buf_clk cell_13438 ( .C (clk), .D (signal_18325), .Q (signal_18326) ) ;
    buf_clk cell_13444 ( .C (clk), .D (signal_18331), .Q (signal_18332) ) ;
    buf_clk cell_13450 ( .C (clk), .D (signal_18337), .Q (signal_18338) ) ;
    buf_clk cell_13456 ( .C (clk), .D (signal_18343), .Q (signal_18344) ) ;
    buf_clk cell_13462 ( .C (clk), .D (signal_18349), .Q (signal_18350) ) ;
    buf_clk cell_13468 ( .C (clk), .D (signal_18355), .Q (signal_18356) ) ;
    buf_clk cell_13474 ( .C (clk), .D (signal_18361), .Q (signal_18362) ) ;
    buf_clk cell_13480 ( .C (clk), .D (signal_18367), .Q (signal_18368) ) ;
    buf_clk cell_13486 ( .C (clk), .D (signal_18373), .Q (signal_18374) ) ;
    buf_clk cell_13492 ( .C (clk), .D (signal_18379), .Q (signal_18380) ) ;
    buf_clk cell_13498 ( .C (clk), .D (signal_18385), .Q (signal_18386) ) ;
    buf_clk cell_13504 ( .C (clk), .D (signal_18391), .Q (signal_18392) ) ;
    buf_clk cell_13510 ( .C (clk), .D (signal_18397), .Q (signal_18398) ) ;
    buf_clk cell_13516 ( .C (clk), .D (signal_18403), .Q (signal_18404) ) ;
    buf_clk cell_13522 ( .C (clk), .D (signal_18409), .Q (signal_18410) ) ;
    buf_clk cell_13528 ( .C (clk), .D (signal_18415), .Q (signal_18416) ) ;
    buf_clk cell_13534 ( .C (clk), .D (signal_18421), .Q (signal_18422) ) ;
    buf_clk cell_13540 ( .C (clk), .D (signal_18427), .Q (signal_18428) ) ;
    buf_clk cell_13546 ( .C (clk), .D (signal_18433), .Q (signal_18434) ) ;
    buf_clk cell_13552 ( .C (clk), .D (signal_18439), .Q (signal_18440) ) ;
    buf_clk cell_13558 ( .C (clk), .D (signal_18445), .Q (signal_18446) ) ;
    buf_clk cell_13564 ( .C (clk), .D (signal_18451), .Q (signal_18452) ) ;
    buf_clk cell_13570 ( .C (clk), .D (signal_18457), .Q (signal_18458) ) ;
    buf_clk cell_13576 ( .C (clk), .D (signal_18463), .Q (signal_18464) ) ;
    buf_clk cell_13582 ( .C (clk), .D (signal_18469), .Q (signal_18470) ) ;
    buf_clk cell_13588 ( .C (clk), .D (signal_18475), .Q (signal_18476) ) ;
    buf_clk cell_13594 ( .C (clk), .D (signal_18481), .Q (signal_18482) ) ;
    buf_clk cell_13600 ( .C (clk), .D (signal_18487), .Q (signal_18488) ) ;
    buf_clk cell_13606 ( .C (clk), .D (signal_18493), .Q (signal_18494) ) ;
    buf_clk cell_13612 ( .C (clk), .D (signal_18499), .Q (signal_18500) ) ;
    buf_clk cell_13618 ( .C (clk), .D (signal_18505), .Q (signal_18506) ) ;
    buf_clk cell_13624 ( .C (clk), .D (signal_18511), .Q (signal_18512) ) ;
    buf_clk cell_13630 ( .C (clk), .D (signal_18517), .Q (signal_18518) ) ;
    buf_clk cell_13636 ( .C (clk), .D (signal_18523), .Q (signal_18524) ) ;
    buf_clk cell_13642 ( .C (clk), .D (signal_18529), .Q (signal_18530) ) ;
    buf_clk cell_13648 ( .C (clk), .D (signal_18535), .Q (signal_18536) ) ;
    buf_clk cell_13654 ( .C (clk), .D (signal_18541), .Q (signal_18542) ) ;
    buf_clk cell_13660 ( .C (clk), .D (signal_18547), .Q (signal_18548) ) ;
    buf_clk cell_13666 ( .C (clk), .D (signal_18553), .Q (signal_18554) ) ;
    buf_clk cell_13672 ( .C (clk), .D (signal_18559), .Q (signal_18560) ) ;
    buf_clk cell_13678 ( .C (clk), .D (signal_18565), .Q (signal_18566) ) ;
    buf_clk cell_13684 ( .C (clk), .D (signal_18571), .Q (signal_18572) ) ;
    buf_clk cell_13690 ( .C (clk), .D (signal_18577), .Q (signal_18578) ) ;
    buf_clk cell_13696 ( .C (clk), .D (signal_18583), .Q (signal_18584) ) ;
    buf_clk cell_13702 ( .C (clk), .D (signal_18589), .Q (signal_18590) ) ;
    buf_clk cell_13708 ( .C (clk), .D (signal_18595), .Q (signal_18596) ) ;
    buf_clk cell_13714 ( .C (clk), .D (signal_18601), .Q (signal_18602) ) ;
    buf_clk cell_13720 ( .C (clk), .D (signal_18607), .Q (signal_18608) ) ;
    buf_clk cell_13726 ( .C (clk), .D (signal_18613), .Q (signal_18614) ) ;
    buf_clk cell_13732 ( .C (clk), .D (signal_18619), .Q (signal_18620) ) ;
    buf_clk cell_13738 ( .C (clk), .D (signal_18625), .Q (signal_18626) ) ;
    buf_clk cell_13744 ( .C (clk), .D (signal_18631), .Q (signal_18632) ) ;
    buf_clk cell_13750 ( .C (clk), .D (signal_18637), .Q (signal_18638) ) ;
    buf_clk cell_13756 ( .C (clk), .D (signal_18643), .Q (signal_18644) ) ;
    buf_clk cell_13762 ( .C (clk), .D (signal_18649), .Q (signal_18650) ) ;
    buf_clk cell_13768 ( .C (clk), .D (signal_18655), .Q (signal_18656) ) ;
    buf_clk cell_13774 ( .C (clk), .D (signal_18661), .Q (signal_18662) ) ;
    buf_clk cell_13780 ( .C (clk), .D (signal_18667), .Q (signal_18668) ) ;
    buf_clk cell_13786 ( .C (clk), .D (signal_18673), .Q (signal_18674) ) ;
    buf_clk cell_13792 ( .C (clk), .D (signal_18679), .Q (signal_18680) ) ;
    buf_clk cell_13798 ( .C (clk), .D (signal_18685), .Q (signal_18686) ) ;
    buf_clk cell_13804 ( .C (clk), .D (signal_18691), .Q (signal_18692) ) ;
    buf_clk cell_13810 ( .C (clk), .D (signal_18697), .Q (signal_18698) ) ;
    buf_clk cell_13816 ( .C (clk), .D (signal_18703), .Q (signal_18704) ) ;
    buf_clk cell_13822 ( .C (clk), .D (signal_18709), .Q (signal_18710) ) ;
    buf_clk cell_13828 ( .C (clk), .D (signal_18715), .Q (signal_18716) ) ;
    buf_clk cell_13834 ( .C (clk), .D (signal_18721), .Q (signal_18722) ) ;
    buf_clk cell_13840 ( .C (clk), .D (signal_18727), .Q (signal_18728) ) ;
    buf_clk cell_13846 ( .C (clk), .D (signal_18733), .Q (signal_18734) ) ;
    buf_clk cell_13852 ( .C (clk), .D (signal_18739), .Q (signal_18740) ) ;
    buf_clk cell_13858 ( .C (clk), .D (signal_18745), .Q (signal_18746) ) ;
    buf_clk cell_13864 ( .C (clk), .D (signal_18751), .Q (signal_18752) ) ;
    buf_clk cell_13870 ( .C (clk), .D (signal_18757), .Q (signal_18758) ) ;
    buf_clk cell_13876 ( .C (clk), .D (signal_18763), .Q (signal_18764) ) ;
    buf_clk cell_13882 ( .C (clk), .D (signal_18769), .Q (signal_18770) ) ;
    buf_clk cell_13888 ( .C (clk), .D (signal_18775), .Q (signal_18776) ) ;
    buf_clk cell_13894 ( .C (clk), .D (signal_18781), .Q (signal_18782) ) ;
    buf_clk cell_13900 ( .C (clk), .D (signal_18787), .Q (signal_18788) ) ;
    buf_clk cell_13906 ( .C (clk), .D (signal_18793), .Q (signal_18794) ) ;
    buf_clk cell_13912 ( .C (clk), .D (signal_18799), .Q (signal_18800) ) ;
    buf_clk cell_13918 ( .C (clk), .D (signal_18805), .Q (signal_18806) ) ;
    buf_clk cell_13924 ( .C (clk), .D (signal_18811), .Q (signal_18812) ) ;
    buf_clk cell_13930 ( .C (clk), .D (signal_18817), .Q (signal_18818) ) ;
    buf_clk cell_13936 ( .C (clk), .D (signal_18823), .Q (signal_18824) ) ;
    buf_clk cell_13942 ( .C (clk), .D (signal_18829), .Q (signal_18830) ) ;
    buf_clk cell_13948 ( .C (clk), .D (signal_18835), .Q (signal_18836) ) ;
    buf_clk cell_13954 ( .C (clk), .D (signal_18841), .Q (signal_18842) ) ;
    buf_clk cell_13960 ( .C (clk), .D (signal_18847), .Q (signal_18848) ) ;
    buf_clk cell_13966 ( .C (clk), .D (signal_18853), .Q (signal_18854) ) ;
    buf_clk cell_13972 ( .C (clk), .D (signal_18859), .Q (signal_18860) ) ;
    buf_clk cell_13978 ( .C (clk), .D (signal_18865), .Q (signal_18866) ) ;
    buf_clk cell_13984 ( .C (clk), .D (signal_18871), .Q (signal_18872) ) ;
    buf_clk cell_13990 ( .C (clk), .D (signal_18877), .Q (signal_18878) ) ;
    buf_clk cell_13996 ( .C (clk), .D (signal_18883), .Q (signal_18884) ) ;
    buf_clk cell_14002 ( .C (clk), .D (signal_18889), .Q (signal_18890) ) ;
    buf_clk cell_14008 ( .C (clk), .D (signal_18895), .Q (signal_18896) ) ;
    buf_clk cell_14014 ( .C (clk), .D (signal_18901), .Q (signal_18902) ) ;
    buf_clk cell_14020 ( .C (clk), .D (signal_18907), .Q (signal_18908) ) ;
    buf_clk cell_14026 ( .C (clk), .D (signal_18913), .Q (signal_18914) ) ;
    buf_clk cell_14032 ( .C (clk), .D (signal_18919), .Q (signal_18920) ) ;
    buf_clk cell_14038 ( .C (clk), .D (signal_18925), .Q (signal_18926) ) ;
    buf_clk cell_14044 ( .C (clk), .D (signal_18931), .Q (signal_18932) ) ;
    buf_clk cell_14050 ( .C (clk), .D (signal_18937), .Q (signal_18938) ) ;
    buf_clk cell_14056 ( .C (clk), .D (signal_18943), .Q (signal_18944) ) ;
    buf_clk cell_14062 ( .C (clk), .D (signal_18949), .Q (signal_18950) ) ;
    buf_clk cell_14068 ( .C (clk), .D (signal_18955), .Q (signal_18956) ) ;
    buf_clk cell_14074 ( .C (clk), .D (signal_18961), .Q (signal_18962) ) ;
    buf_clk cell_14080 ( .C (clk), .D (signal_18967), .Q (signal_18968) ) ;
    buf_clk cell_14086 ( .C (clk), .D (signal_18973), .Q (signal_18974) ) ;
    buf_clk cell_14092 ( .C (clk), .D (signal_18979), .Q (signal_18980) ) ;
    buf_clk cell_14098 ( .C (clk), .D (signal_18985), .Q (signal_18986) ) ;
    buf_clk cell_14104 ( .C (clk), .D (signal_18991), .Q (signal_18992) ) ;
    buf_clk cell_14110 ( .C (clk), .D (signal_18997), .Q (signal_18998) ) ;
    buf_clk cell_14116 ( .C (clk), .D (signal_19003), .Q (signal_19004) ) ;
    buf_clk cell_14122 ( .C (clk), .D (signal_19009), .Q (signal_19010) ) ;
    buf_clk cell_14128 ( .C (clk), .D (signal_19015), .Q (signal_19016) ) ;
    buf_clk cell_14134 ( .C (clk), .D (signal_19021), .Q (signal_19022) ) ;
    buf_clk cell_14140 ( .C (clk), .D (signal_19027), .Q (signal_19028) ) ;
    buf_clk cell_14146 ( .C (clk), .D (signal_19033), .Q (signal_19034) ) ;
    buf_clk cell_14152 ( .C (clk), .D (signal_19039), .Q (signal_19040) ) ;
    buf_clk cell_14158 ( .C (clk), .D (signal_19045), .Q (signal_19046) ) ;
    buf_clk cell_14164 ( .C (clk), .D (signal_19051), .Q (signal_19052) ) ;
    buf_clk cell_14170 ( .C (clk), .D (signal_19057), .Q (signal_19058) ) ;
    buf_clk cell_14176 ( .C (clk), .D (signal_19063), .Q (signal_19064) ) ;
    buf_clk cell_14182 ( .C (clk), .D (signal_19069), .Q (signal_19070) ) ;
    buf_clk cell_14188 ( .C (clk), .D (signal_19075), .Q (signal_19076) ) ;
    buf_clk cell_14194 ( .C (clk), .D (signal_19081), .Q (signal_19082) ) ;
    buf_clk cell_14200 ( .C (clk), .D (signal_19087), .Q (signal_19088) ) ;
    buf_clk cell_14206 ( .C (clk), .D (signal_19093), .Q (signal_19094) ) ;
    buf_clk cell_14212 ( .C (clk), .D (signal_19099), .Q (signal_19100) ) ;
    buf_clk cell_14218 ( .C (clk), .D (signal_19105), .Q (signal_19106) ) ;
    buf_clk cell_14224 ( .C (clk), .D (signal_19111), .Q (signal_19112) ) ;
    buf_clk cell_14230 ( .C (clk), .D (signal_19117), .Q (signal_19118) ) ;
    buf_clk cell_14236 ( .C (clk), .D (signal_19123), .Q (signal_19124) ) ;
    buf_clk cell_14242 ( .C (clk), .D (signal_19129), .Q (signal_19130) ) ;
    buf_clk cell_14248 ( .C (clk), .D (signal_19135), .Q (signal_19136) ) ;
    buf_clk cell_14254 ( .C (clk), .D (signal_19141), .Q (signal_19142) ) ;
    buf_clk cell_14260 ( .C (clk), .D (signal_19147), .Q (signal_19148) ) ;
    buf_clk cell_14266 ( .C (clk), .D (signal_19153), .Q (signal_19154) ) ;
    buf_clk cell_14272 ( .C (clk), .D (signal_19159), .Q (signal_19160) ) ;
    buf_clk cell_14278 ( .C (clk), .D (signal_19165), .Q (signal_19166) ) ;
    buf_clk cell_14284 ( .C (clk), .D (signal_19171), .Q (signal_19172) ) ;
    buf_clk cell_14290 ( .C (clk), .D (signal_19177), .Q (signal_19178) ) ;
    buf_clk cell_14296 ( .C (clk), .D (signal_19183), .Q (signal_19184) ) ;
    buf_clk cell_14302 ( .C (clk), .D (signal_19189), .Q (signal_19190) ) ;
    buf_clk cell_14308 ( .C (clk), .D (signal_19195), .Q (signal_19196) ) ;
    buf_clk cell_14314 ( .C (clk), .D (signal_19201), .Q (signal_19202) ) ;
    buf_clk cell_14320 ( .C (clk), .D (signal_19207), .Q (signal_19208) ) ;
    buf_clk cell_14326 ( .C (clk), .D (signal_19213), .Q (signal_19214) ) ;
    buf_clk cell_14332 ( .C (clk), .D (signal_19219), .Q (signal_19220) ) ;
    buf_clk cell_14338 ( .C (clk), .D (signal_19225), .Q (signal_19226) ) ;
    buf_clk cell_14344 ( .C (clk), .D (signal_19231), .Q (signal_19232) ) ;
    buf_clk cell_14350 ( .C (clk), .D (signal_19237), .Q (signal_19238) ) ;
    buf_clk cell_14356 ( .C (clk), .D (signal_19243), .Q (signal_19244) ) ;
    buf_clk cell_14362 ( .C (clk), .D (signal_19249), .Q (signal_19250) ) ;
    buf_clk cell_14368 ( .C (clk), .D (signal_19255), .Q (signal_19256) ) ;
    buf_clk cell_14374 ( .C (clk), .D (signal_19261), .Q (signal_19262) ) ;
    buf_clk cell_14380 ( .C (clk), .D (signal_19267), .Q (signal_19268) ) ;
    buf_clk cell_14386 ( .C (clk), .D (signal_19273), .Q (signal_19274) ) ;
    buf_clk cell_14392 ( .C (clk), .D (signal_19279), .Q (signal_19280) ) ;
    buf_clk cell_14398 ( .C (clk), .D (signal_19285), .Q (signal_19286) ) ;
    buf_clk cell_14404 ( .C (clk), .D (signal_19291), .Q (signal_19292) ) ;
    buf_clk cell_14410 ( .C (clk), .D (signal_19297), .Q (signal_19298) ) ;
    buf_clk cell_14416 ( .C (clk), .D (signal_19303), .Q (signal_19304) ) ;
    buf_clk cell_14422 ( .C (clk), .D (signal_19309), .Q (signal_19310) ) ;
    buf_clk cell_14428 ( .C (clk), .D (signal_19315), .Q (signal_19316) ) ;
    buf_clk cell_14434 ( .C (clk), .D (signal_19321), .Q (signal_19322) ) ;
    buf_clk cell_14440 ( .C (clk), .D (signal_19327), .Q (signal_19328) ) ;
    buf_clk cell_14446 ( .C (clk), .D (signal_19333), .Q (signal_19334) ) ;
    buf_clk cell_14452 ( .C (clk), .D (signal_19339), .Q (signal_19340) ) ;
    buf_clk cell_14458 ( .C (clk), .D (signal_19345), .Q (signal_19346) ) ;
    buf_clk cell_14464 ( .C (clk), .D (signal_19351), .Q (signal_19352) ) ;
    buf_clk cell_14470 ( .C (clk), .D (signal_19357), .Q (signal_19358) ) ;
    buf_clk cell_14476 ( .C (clk), .D (signal_19363), .Q (signal_19364) ) ;
    buf_clk cell_14482 ( .C (clk), .D (signal_19369), .Q (signal_19370) ) ;
    buf_clk cell_14488 ( .C (clk), .D (signal_19375), .Q (signal_19376) ) ;
    buf_clk cell_14494 ( .C (clk), .D (signal_19381), .Q (signal_19382) ) ;
    buf_clk cell_14500 ( .C (clk), .D (signal_19387), .Q (signal_19388) ) ;
    buf_clk cell_14506 ( .C (clk), .D (signal_19393), .Q (signal_19394) ) ;
    buf_clk cell_14512 ( .C (clk), .D (signal_19399), .Q (signal_19400) ) ;
    buf_clk cell_14518 ( .C (clk), .D (signal_19405), .Q (signal_19406) ) ;
    buf_clk cell_14524 ( .C (clk), .D (signal_19411), .Q (signal_19412) ) ;
    buf_clk cell_14530 ( .C (clk), .D (signal_19417), .Q (signal_19418) ) ;
    buf_clk cell_14536 ( .C (clk), .D (signal_19423), .Q (signal_19424) ) ;
    buf_clk cell_14542 ( .C (clk), .D (signal_19429), .Q (signal_19430) ) ;
    buf_clk cell_14548 ( .C (clk), .D (signal_19435), .Q (signal_19436) ) ;
    buf_clk cell_14554 ( .C (clk), .D (signal_19441), .Q (signal_19442) ) ;
    buf_clk cell_14560 ( .C (clk), .D (signal_19447), .Q (signal_19448) ) ;
    buf_clk cell_14566 ( .C (clk), .D (signal_19453), .Q (signal_19454) ) ;
    buf_clk cell_14572 ( .C (clk), .D (signal_19459), .Q (signal_19460) ) ;
    buf_clk cell_14578 ( .C (clk), .D (signal_19465), .Q (signal_19466) ) ;
    buf_clk cell_14584 ( .C (clk), .D (signal_19471), .Q (signal_19472) ) ;
    buf_clk cell_14590 ( .C (clk), .D (signal_19477), .Q (signal_19478) ) ;
    buf_clk cell_14596 ( .C (clk), .D (signal_19483), .Q (signal_19484) ) ;
    buf_clk cell_14602 ( .C (clk), .D (signal_19489), .Q (signal_19490) ) ;
    buf_clk cell_14608 ( .C (clk), .D (signal_19495), .Q (signal_19496) ) ;
    buf_clk cell_14614 ( .C (clk), .D (signal_19501), .Q (signal_19502) ) ;
    buf_clk cell_14620 ( .C (clk), .D (signal_19507), .Q (signal_19508) ) ;
    buf_clk cell_14626 ( .C (clk), .D (signal_19513), .Q (signal_19514) ) ;
    buf_clk cell_14632 ( .C (clk), .D (signal_19519), .Q (signal_19520) ) ;
    buf_clk cell_14638 ( .C (clk), .D (signal_19525), .Q (signal_19526) ) ;
    buf_clk cell_14644 ( .C (clk), .D (signal_19531), .Q (signal_19532) ) ;
    buf_clk cell_14650 ( .C (clk), .D (signal_19537), .Q (signal_19538) ) ;
    buf_clk cell_14656 ( .C (clk), .D (signal_19543), .Q (signal_19544) ) ;
    buf_clk cell_14662 ( .C (clk), .D (signal_19549), .Q (signal_19550) ) ;
    buf_clk cell_14668 ( .C (clk), .D (signal_19555), .Q (signal_19556) ) ;
    buf_clk cell_14674 ( .C (clk), .D (signal_19561), .Q (signal_19562) ) ;
    buf_clk cell_14680 ( .C (clk), .D (signal_19567), .Q (signal_19568) ) ;
    buf_clk cell_14686 ( .C (clk), .D (signal_19573), .Q (signal_19574) ) ;
    buf_clk cell_14692 ( .C (clk), .D (signal_19579), .Q (signal_19580) ) ;
    buf_clk cell_14698 ( .C (clk), .D (signal_19585), .Q (signal_19586) ) ;
    buf_clk cell_14704 ( .C (clk), .D (signal_19591), .Q (signal_19592) ) ;
    buf_clk cell_14710 ( .C (clk), .D (signal_19597), .Q (signal_19598) ) ;
    buf_clk cell_14716 ( .C (clk), .D (signal_19603), .Q (signal_19604) ) ;
    buf_clk cell_14722 ( .C (clk), .D (signal_19609), .Q (signal_19610) ) ;
    buf_clk cell_14728 ( .C (clk), .D (signal_19615), .Q (signal_19616) ) ;
    buf_clk cell_14734 ( .C (clk), .D (signal_19621), .Q (signal_19622) ) ;
    buf_clk cell_14740 ( .C (clk), .D (signal_19627), .Q (signal_19628) ) ;
    buf_clk cell_14746 ( .C (clk), .D (signal_19633), .Q (signal_19634) ) ;
    buf_clk cell_14752 ( .C (clk), .D (signal_19639), .Q (signal_19640) ) ;
    buf_clk cell_14758 ( .C (clk), .D (signal_19645), .Q (signal_19646) ) ;
    buf_clk cell_14764 ( .C (clk), .D (signal_19651), .Q (signal_19652) ) ;
    buf_clk cell_14770 ( .C (clk), .D (signal_19657), .Q (signal_19658) ) ;
    buf_clk cell_14776 ( .C (clk), .D (signal_19663), .Q (signal_19664) ) ;
    buf_clk cell_14782 ( .C (clk), .D (signal_19669), .Q (signal_19670) ) ;
    buf_clk cell_14788 ( .C (clk), .D (signal_19675), .Q (signal_19676) ) ;
    buf_clk cell_14794 ( .C (clk), .D (signal_19681), .Q (signal_19682) ) ;
    buf_clk cell_14800 ( .C (clk), .D (signal_19687), .Q (signal_19688) ) ;
    buf_clk cell_14806 ( .C (clk), .D (signal_19693), .Q (signal_19694) ) ;
    buf_clk cell_14812 ( .C (clk), .D (signal_19699), .Q (signal_19700) ) ;
    buf_clk cell_14818 ( .C (clk), .D (signal_19705), .Q (signal_19706) ) ;
    buf_clk cell_14824 ( .C (clk), .D (signal_19711), .Q (signal_19712) ) ;
    buf_clk cell_14830 ( .C (clk), .D (signal_19717), .Q (signal_19718) ) ;
    buf_clk cell_14836 ( .C (clk), .D (signal_19723), .Q (signal_19724) ) ;
    buf_clk cell_14842 ( .C (clk), .D (signal_19729), .Q (signal_19730) ) ;
    buf_clk cell_14848 ( .C (clk), .D (signal_19735), .Q (signal_19736) ) ;
    buf_clk cell_14854 ( .C (clk), .D (signal_19741), .Q (signal_19742) ) ;
    buf_clk cell_14860 ( .C (clk), .D (signal_19747), .Q (signal_19748) ) ;
    buf_clk cell_14866 ( .C (clk), .D (signal_19753), .Q (signal_19754) ) ;
    buf_clk cell_14872 ( .C (clk), .D (signal_19759), .Q (signal_19760) ) ;
    buf_clk cell_14878 ( .C (clk), .D (signal_19765), .Q (signal_19766) ) ;
    buf_clk cell_14884 ( .C (clk), .D (signal_19771), .Q (signal_19772) ) ;
    buf_clk cell_14890 ( .C (clk), .D (signal_19777), .Q (signal_19778) ) ;
    buf_clk cell_14896 ( .C (clk), .D (signal_19783), .Q (signal_19784) ) ;
    buf_clk cell_14902 ( .C (clk), .D (signal_19789), .Q (signal_19790) ) ;
    buf_clk cell_14908 ( .C (clk), .D (signal_19795), .Q (signal_19796) ) ;
    buf_clk cell_14914 ( .C (clk), .D (signal_19801), .Q (signal_19802) ) ;
    buf_clk cell_14920 ( .C (clk), .D (signal_19807), .Q (signal_19808) ) ;
    buf_clk cell_14926 ( .C (clk), .D (signal_19813), .Q (signal_19814) ) ;
    buf_clk cell_14932 ( .C (clk), .D (signal_19819), .Q (signal_19820) ) ;
    buf_clk cell_14938 ( .C (clk), .D (signal_19825), .Q (signal_19826) ) ;
    buf_clk cell_14944 ( .C (clk), .D (signal_19831), .Q (signal_19832) ) ;
    buf_clk cell_14950 ( .C (clk), .D (signal_19837), .Q (signal_19838) ) ;
    buf_clk cell_14956 ( .C (clk), .D (signal_19843), .Q (signal_19844) ) ;
    buf_clk cell_14962 ( .C (clk), .D (signal_19849), .Q (signal_19850) ) ;
    buf_clk cell_14968 ( .C (clk), .D (signal_19855), .Q (signal_19856) ) ;
    buf_clk cell_14974 ( .C (clk), .D (signal_19861), .Q (signal_19862) ) ;
    buf_clk cell_14980 ( .C (clk), .D (signal_19867), .Q (signal_19868) ) ;
    buf_clk cell_14986 ( .C (clk), .D (signal_19873), .Q (signal_19874) ) ;
    buf_clk cell_14992 ( .C (clk), .D (signal_19879), .Q (signal_19880) ) ;
    buf_clk cell_14998 ( .C (clk), .D (signal_19885), .Q (signal_19886) ) ;
    buf_clk cell_15004 ( .C (clk), .D (signal_19891), .Q (signal_19892) ) ;
    buf_clk cell_15010 ( .C (clk), .D (signal_19897), .Q (signal_19898) ) ;
    buf_clk cell_15016 ( .C (clk), .D (signal_19903), .Q (signal_19904) ) ;
    buf_clk cell_15022 ( .C (clk), .D (signal_19909), .Q (signal_19910) ) ;
    buf_clk cell_15028 ( .C (clk), .D (signal_19915), .Q (signal_19916) ) ;
    buf_clk cell_15034 ( .C (clk), .D (signal_19921), .Q (signal_19922) ) ;
    buf_clk cell_15040 ( .C (clk), .D (signal_19927), .Q (signal_19928) ) ;
    buf_clk cell_15046 ( .C (clk), .D (signal_19933), .Q (signal_19934) ) ;
    buf_clk cell_15052 ( .C (clk), .D (signal_19939), .Q (signal_19940) ) ;
    buf_clk cell_15058 ( .C (clk), .D (signal_19945), .Q (signal_19946) ) ;
    buf_clk cell_15064 ( .C (clk), .D (signal_19951), .Q (signal_19952) ) ;
    buf_clk cell_15070 ( .C (clk), .D (signal_19957), .Q (signal_19958) ) ;
    buf_clk cell_15076 ( .C (clk), .D (signal_19963), .Q (signal_19964) ) ;
    buf_clk cell_15082 ( .C (clk), .D (signal_19969), .Q (signal_19970) ) ;
    buf_clk cell_15088 ( .C (clk), .D (signal_19975), .Q (signal_19976) ) ;
    buf_clk cell_15094 ( .C (clk), .D (signal_19981), .Q (signal_19982) ) ;
    buf_clk cell_15100 ( .C (clk), .D (signal_19987), .Q (signal_19988) ) ;
    buf_clk cell_15106 ( .C (clk), .D (signal_19993), .Q (signal_19994) ) ;
    buf_clk cell_15112 ( .C (clk), .D (signal_19999), .Q (signal_20000) ) ;
    buf_clk cell_15118 ( .C (clk), .D (signal_20005), .Q (signal_20006) ) ;
    buf_clk cell_15124 ( .C (clk), .D (signal_20011), .Q (signal_20012) ) ;
    buf_clk cell_15130 ( .C (clk), .D (signal_20017), .Q (signal_20018) ) ;
    buf_clk cell_15136 ( .C (clk), .D (signal_20023), .Q (signal_20024) ) ;
    buf_clk cell_15142 ( .C (clk), .D (signal_20029), .Q (signal_20030) ) ;
    buf_clk cell_15148 ( .C (clk), .D (signal_20035), .Q (signal_20036) ) ;
    buf_clk cell_15154 ( .C (clk), .D (signal_20041), .Q (signal_20042) ) ;
    buf_clk cell_15160 ( .C (clk), .D (signal_20047), .Q (signal_20048) ) ;
    buf_clk cell_15166 ( .C (clk), .D (signal_20053), .Q (signal_20054) ) ;
    buf_clk cell_15172 ( .C (clk), .D (signal_20059), .Q (signal_20060) ) ;
    buf_clk cell_15178 ( .C (clk), .D (signal_20065), .Q (signal_20066) ) ;
    buf_clk cell_15184 ( .C (clk), .D (signal_20071), .Q (signal_20072) ) ;
    buf_clk cell_15190 ( .C (clk), .D (signal_20077), .Q (signal_20078) ) ;
    buf_clk cell_15196 ( .C (clk), .D (signal_20083), .Q (signal_20084) ) ;
    buf_clk cell_15202 ( .C (clk), .D (signal_20089), .Q (signal_20090) ) ;
    buf_clk cell_15208 ( .C (clk), .D (signal_20095), .Q (signal_20096) ) ;
    buf_clk cell_15214 ( .C (clk), .D (signal_20101), .Q (signal_20102) ) ;
    buf_clk cell_15220 ( .C (clk), .D (signal_20107), .Q (signal_20108) ) ;
    buf_clk cell_15226 ( .C (clk), .D (signal_20113), .Q (signal_20114) ) ;
    buf_clk cell_15232 ( .C (clk), .D (signal_20119), .Q (signal_20120) ) ;
    buf_clk cell_15238 ( .C (clk), .D (signal_20125), .Q (signal_20126) ) ;
    buf_clk cell_15244 ( .C (clk), .D (signal_20131), .Q (signal_20132) ) ;
    buf_clk cell_15250 ( .C (clk), .D (signal_20137), .Q (signal_20138) ) ;
    buf_clk cell_15256 ( .C (clk), .D (signal_20143), .Q (signal_20144) ) ;
    buf_clk cell_15262 ( .C (clk), .D (signal_20149), .Q (signal_20150) ) ;
    buf_clk cell_15268 ( .C (clk), .D (signal_20155), .Q (signal_20156) ) ;
    buf_clk cell_15274 ( .C (clk), .D (signal_20161), .Q (signal_20162) ) ;
    buf_clk cell_15280 ( .C (clk), .D (signal_20167), .Q (signal_20168) ) ;
    buf_clk cell_15286 ( .C (clk), .D (signal_20173), .Q (signal_20174) ) ;
    buf_clk cell_15292 ( .C (clk), .D (signal_20179), .Q (signal_20180) ) ;
    buf_clk cell_15298 ( .C (clk), .D (signal_20185), .Q (signal_20186) ) ;
    buf_clk cell_15304 ( .C (clk), .D (signal_20191), .Q (signal_20192) ) ;
    buf_clk cell_15310 ( .C (clk), .D (signal_20197), .Q (signal_20198) ) ;
    buf_clk cell_15316 ( .C (clk), .D (signal_20203), .Q (signal_20204) ) ;
    buf_clk cell_15322 ( .C (clk), .D (signal_20209), .Q (signal_20210) ) ;
    buf_clk cell_15328 ( .C (clk), .D (signal_20215), .Q (signal_20216) ) ;
    buf_clk cell_15334 ( .C (clk), .D (signal_20221), .Q (signal_20222) ) ;
    buf_clk cell_15340 ( .C (clk), .D (signal_20227), .Q (signal_20228) ) ;
    buf_clk cell_15346 ( .C (clk), .D (signal_20233), .Q (signal_20234) ) ;
    buf_clk cell_15352 ( .C (clk), .D (signal_20239), .Q (signal_20240) ) ;
    buf_clk cell_15358 ( .C (clk), .D (signal_20245), .Q (signal_20246) ) ;
    buf_clk cell_15364 ( .C (clk), .D (signal_20251), .Q (signal_20252) ) ;
    buf_clk cell_15370 ( .C (clk), .D (signal_20257), .Q (signal_20258) ) ;
    buf_clk cell_15376 ( .C (clk), .D (signal_20263), .Q (signal_20264) ) ;
    buf_clk cell_15382 ( .C (clk), .D (signal_20269), .Q (signal_20270) ) ;
    buf_clk cell_15388 ( .C (clk), .D (signal_20275), .Q (signal_20276) ) ;
    buf_clk cell_15394 ( .C (clk), .D (signal_20281), .Q (signal_20282) ) ;
    buf_clk cell_15400 ( .C (clk), .D (signal_20287), .Q (signal_20288) ) ;
    buf_clk cell_15406 ( .C (clk), .D (signal_20293), .Q (signal_20294) ) ;
    buf_clk cell_15412 ( .C (clk), .D (signal_20299), .Q (signal_20300) ) ;
    buf_clk cell_15418 ( .C (clk), .D (signal_20305), .Q (signal_20306) ) ;
    buf_clk cell_15424 ( .C (clk), .D (signal_20311), .Q (signal_20312) ) ;
    buf_clk cell_15430 ( .C (clk), .D (signal_20317), .Q (signal_20318) ) ;
    buf_clk cell_15436 ( .C (clk), .D (signal_20323), .Q (signal_20324) ) ;
    buf_clk cell_15442 ( .C (clk), .D (signal_20329), .Q (signal_20330) ) ;
    buf_clk cell_15448 ( .C (clk), .D (signal_20335), .Q (signal_20336) ) ;
    buf_clk cell_15454 ( .C (clk), .D (signal_20341), .Q (signal_20342) ) ;
    buf_clk cell_15460 ( .C (clk), .D (signal_20347), .Q (signal_20348) ) ;
    buf_clk cell_15466 ( .C (clk), .D (signal_20353), .Q (signal_20354) ) ;
    buf_clk cell_15472 ( .C (clk), .D (signal_20359), .Q (signal_20360) ) ;
    buf_clk cell_15478 ( .C (clk), .D (signal_20365), .Q (signal_20366) ) ;
    buf_clk cell_15484 ( .C (clk), .D (signal_20371), .Q (signal_20372) ) ;
    buf_clk cell_15490 ( .C (clk), .D (signal_20377), .Q (signal_20378) ) ;
    buf_clk cell_15496 ( .C (clk), .D (signal_20383), .Q (signal_20384) ) ;
    buf_clk cell_15502 ( .C (clk), .D (signal_20389), .Q (signal_20390) ) ;
    buf_clk cell_15508 ( .C (clk), .D (signal_20395), .Q (signal_20396) ) ;
    buf_clk cell_15514 ( .C (clk), .D (signal_20401), .Q (signal_20402) ) ;
    buf_clk cell_15520 ( .C (clk), .D (signal_20407), .Q (signal_20408) ) ;
    buf_clk cell_15526 ( .C (clk), .D (signal_20413), .Q (signal_20414) ) ;
    buf_clk cell_15532 ( .C (clk), .D (signal_20419), .Q (signal_20420) ) ;
    buf_clk cell_15538 ( .C (clk), .D (signal_20425), .Q (signal_20426) ) ;
    buf_clk cell_15544 ( .C (clk), .D (signal_20431), .Q (signal_20432) ) ;
    buf_clk cell_15550 ( .C (clk), .D (signal_20437), .Q (signal_20438) ) ;
    buf_clk cell_15556 ( .C (clk), .D (signal_20443), .Q (signal_20444) ) ;
    buf_clk cell_15562 ( .C (clk), .D (signal_20449), .Q (signal_20450) ) ;
    buf_clk cell_15568 ( .C (clk), .D (signal_20455), .Q (signal_20456) ) ;
    buf_clk cell_15574 ( .C (clk), .D (signal_20461), .Q (signal_20462) ) ;
    buf_clk cell_15580 ( .C (clk), .D (signal_20467), .Q (signal_20468) ) ;
    buf_clk cell_15586 ( .C (clk), .D (signal_20473), .Q (signal_20474) ) ;
    buf_clk cell_15592 ( .C (clk), .D (signal_20479), .Q (signal_20480) ) ;
    buf_clk cell_15598 ( .C (clk), .D (signal_20485), .Q (signal_20486) ) ;
    buf_clk cell_15604 ( .C (clk), .D (signal_20491), .Q (signal_20492) ) ;
    buf_clk cell_15610 ( .C (clk), .D (signal_20497), .Q (signal_20498) ) ;
    buf_clk cell_15616 ( .C (clk), .D (signal_20503), .Q (signal_20504) ) ;
    buf_clk cell_15622 ( .C (clk), .D (signal_20509), .Q (signal_20510) ) ;
    buf_clk cell_15628 ( .C (clk), .D (signal_20515), .Q (signal_20516) ) ;
    buf_clk cell_15634 ( .C (clk), .D (signal_20521), .Q (signal_20522) ) ;
    buf_clk cell_15640 ( .C (clk), .D (signal_20527), .Q (signal_20528) ) ;
    buf_clk cell_15646 ( .C (clk), .D (signal_20533), .Q (signal_20534) ) ;
    buf_clk cell_15652 ( .C (clk), .D (signal_20539), .Q (signal_20540) ) ;
    buf_clk cell_15658 ( .C (clk), .D (signal_20545), .Q (signal_20546) ) ;
    buf_clk cell_15664 ( .C (clk), .D (signal_20551), .Q (signal_20552) ) ;
    buf_clk cell_15670 ( .C (clk), .D (signal_20557), .Q (signal_20558) ) ;
    buf_clk cell_15676 ( .C (clk), .D (signal_20563), .Q (signal_20564) ) ;
    buf_clk cell_15682 ( .C (clk), .D (signal_20569), .Q (signal_20570) ) ;
    buf_clk cell_15688 ( .C (clk), .D (signal_20575), .Q (signal_20576) ) ;
    buf_clk cell_15694 ( .C (clk), .D (signal_20581), .Q (signal_20582) ) ;
    buf_clk cell_15700 ( .C (clk), .D (signal_20587), .Q (signal_20588) ) ;
    buf_clk cell_15706 ( .C (clk), .D (signal_20593), .Q (signal_20594) ) ;
    buf_clk cell_15712 ( .C (clk), .D (signal_20599), .Q (signal_20600) ) ;
    buf_clk cell_15718 ( .C (clk), .D (signal_20605), .Q (signal_20606) ) ;
    buf_clk cell_15724 ( .C (clk), .D (signal_20611), .Q (signal_20612) ) ;
    buf_clk cell_15730 ( .C (clk), .D (signal_20617), .Q (signal_20618) ) ;
    buf_clk cell_15736 ( .C (clk), .D (signal_20623), .Q (signal_20624) ) ;
    buf_clk cell_15742 ( .C (clk), .D (signal_20629), .Q (signal_20630) ) ;
    buf_clk cell_15748 ( .C (clk), .D (signal_20635), .Q (signal_20636) ) ;
    buf_clk cell_15754 ( .C (clk), .D (signal_20641), .Q (signal_20642) ) ;
    buf_clk cell_15760 ( .C (clk), .D (signal_20647), .Q (signal_20648) ) ;
    buf_clk cell_15766 ( .C (clk), .D (signal_20653), .Q (signal_20654) ) ;
    buf_clk cell_15772 ( .C (clk), .D (signal_20659), .Q (signal_20660) ) ;
    buf_clk cell_15778 ( .C (clk), .D (signal_20665), .Q (signal_20666) ) ;
    buf_clk cell_15784 ( .C (clk), .D (signal_20671), .Q (signal_20672) ) ;
    buf_clk cell_15790 ( .C (clk), .D (signal_20677), .Q (signal_20678) ) ;
    buf_clk cell_15796 ( .C (clk), .D (signal_20683), .Q (signal_20684) ) ;
    buf_clk cell_15802 ( .C (clk), .D (signal_20689), .Q (signal_20690) ) ;
    buf_clk cell_15808 ( .C (clk), .D (signal_20695), .Q (signal_20696) ) ;
    buf_clk cell_15814 ( .C (clk), .D (signal_20701), .Q (signal_20702) ) ;
    buf_clk cell_15820 ( .C (clk), .D (signal_20707), .Q (signal_20708) ) ;
    buf_clk cell_15826 ( .C (clk), .D (signal_20713), .Q (signal_20714) ) ;
    buf_clk cell_15832 ( .C (clk), .D (signal_20719), .Q (signal_20720) ) ;
    buf_clk cell_15838 ( .C (clk), .D (signal_20725), .Q (signal_20726) ) ;
    buf_clk cell_15844 ( .C (clk), .D (signal_20731), .Q (signal_20732) ) ;
    buf_clk cell_15850 ( .C (clk), .D (signal_20737), .Q (signal_20738) ) ;
    buf_clk cell_15856 ( .C (clk), .D (signal_20743), .Q (signal_20744) ) ;
    buf_clk cell_15862 ( .C (clk), .D (signal_20749), .Q (signal_20750) ) ;
    buf_clk cell_15868 ( .C (clk), .D (signal_20755), .Q (signal_20756) ) ;
    buf_clk cell_15874 ( .C (clk), .D (signal_20761), .Q (signal_20762) ) ;
    buf_clk cell_15880 ( .C (clk), .D (signal_20767), .Q (signal_20768) ) ;
    buf_clk cell_15886 ( .C (clk), .D (signal_20773), .Q (signal_20774) ) ;
    buf_clk cell_15892 ( .C (clk), .D (signal_20779), .Q (signal_20780) ) ;
    buf_clk cell_15898 ( .C (clk), .D (signal_20785), .Q (signal_20786) ) ;
    buf_clk cell_15904 ( .C (clk), .D (signal_20791), .Q (signal_20792) ) ;
    buf_clk cell_15910 ( .C (clk), .D (signal_20797), .Q (signal_20798) ) ;
    buf_clk cell_15916 ( .C (clk), .D (signal_20803), .Q (signal_20804) ) ;
    buf_clk cell_15922 ( .C (clk), .D (signal_20809), .Q (signal_20810) ) ;
    buf_clk cell_15928 ( .C (clk), .D (signal_20815), .Q (signal_20816) ) ;
    buf_clk cell_15934 ( .C (clk), .D (signal_20821), .Q (signal_20822) ) ;
    buf_clk cell_15940 ( .C (clk), .D (signal_20827), .Q (signal_20828) ) ;
    buf_clk cell_15946 ( .C (clk), .D (signal_20833), .Q (signal_20834) ) ;
    buf_clk cell_15952 ( .C (clk), .D (signal_20839), .Q (signal_20840) ) ;
    buf_clk cell_15958 ( .C (clk), .D (signal_20845), .Q (signal_20846) ) ;
    buf_clk cell_15964 ( .C (clk), .D (signal_20851), .Q (signal_20852) ) ;
    buf_clk cell_15970 ( .C (clk), .D (signal_20857), .Q (signal_20858) ) ;
    buf_clk cell_15976 ( .C (clk), .D (signal_20863), .Q (signal_20864) ) ;
    buf_clk cell_15982 ( .C (clk), .D (signal_20869), .Q (signal_20870) ) ;
    buf_clk cell_15988 ( .C (clk), .D (signal_20875), .Q (signal_20876) ) ;
    buf_clk cell_15994 ( .C (clk), .D (signal_20881), .Q (signal_20882) ) ;
    buf_clk cell_16000 ( .C (clk), .D (signal_20887), .Q (signal_20888) ) ;
    buf_clk cell_16006 ( .C (clk), .D (signal_20893), .Q (signal_20894) ) ;
    buf_clk cell_16012 ( .C (clk), .D (signal_20899), .Q (signal_20900) ) ;
    buf_clk cell_16018 ( .C (clk), .D (signal_20905), .Q (signal_20906) ) ;
    buf_clk cell_16024 ( .C (clk), .D (signal_20911), .Q (signal_20912) ) ;
    buf_clk cell_16030 ( .C (clk), .D (signal_20917), .Q (signal_20918) ) ;
    buf_clk cell_16036 ( .C (clk), .D (signal_20923), .Q (signal_20924) ) ;
    buf_clk cell_16042 ( .C (clk), .D (signal_20929), .Q (signal_20930) ) ;
    buf_clk cell_16048 ( .C (clk), .D (signal_20935), .Q (signal_20936) ) ;
    buf_clk cell_16054 ( .C (clk), .D (signal_20941), .Q (signal_20942) ) ;
    buf_clk cell_16060 ( .C (clk), .D (signal_20947), .Q (signal_20948) ) ;
    buf_clk cell_16066 ( .C (clk), .D (signal_20953), .Q (signal_20954) ) ;
    buf_clk cell_16072 ( .C (clk), .D (signal_20959), .Q (signal_20960) ) ;
    buf_clk cell_16078 ( .C (clk), .D (signal_20965), .Q (signal_20966) ) ;
    buf_clk cell_16084 ( .C (clk), .D (signal_20971), .Q (signal_20972) ) ;
    buf_clk cell_16090 ( .C (clk), .D (signal_20977), .Q (signal_20978) ) ;
    buf_clk cell_16096 ( .C (clk), .D (signal_20983), .Q (signal_20984) ) ;
    buf_clk cell_16102 ( .C (clk), .D (signal_20989), .Q (signal_20990) ) ;
    buf_clk cell_16108 ( .C (clk), .D (signal_20995), .Q (signal_20996) ) ;
    buf_clk cell_16114 ( .C (clk), .D (signal_21001), .Q (signal_21002) ) ;
    buf_clk cell_16120 ( .C (clk), .D (signal_21007), .Q (signal_21008) ) ;
    buf_clk cell_16126 ( .C (clk), .D (signal_21013), .Q (signal_21014) ) ;
    buf_clk cell_16132 ( .C (clk), .D (signal_21019), .Q (signal_21020) ) ;
    buf_clk cell_16138 ( .C (clk), .D (signal_21025), .Q (signal_21026) ) ;
    buf_clk cell_16144 ( .C (clk), .D (signal_21031), .Q (signal_21032) ) ;
    buf_clk cell_16150 ( .C (clk), .D (signal_21037), .Q (signal_21038) ) ;
    buf_clk cell_16156 ( .C (clk), .D (signal_21043), .Q (signal_21044) ) ;
    buf_clk cell_16162 ( .C (clk), .D (signal_21049), .Q (signal_21050) ) ;
    buf_clk cell_16168 ( .C (clk), .D (signal_21055), .Q (signal_21056) ) ;
    buf_clk cell_16174 ( .C (clk), .D (signal_21061), .Q (signal_21062) ) ;
    buf_clk cell_16180 ( .C (clk), .D (signal_21067), .Q (signal_21068) ) ;
    buf_clk cell_16186 ( .C (clk), .D (signal_21073), .Q (signal_21074) ) ;
    buf_clk cell_16192 ( .C (clk), .D (signal_21079), .Q (signal_21080) ) ;
    buf_clk cell_16198 ( .C (clk), .D (signal_21085), .Q (signal_21086) ) ;
    buf_clk cell_16204 ( .C (clk), .D (signal_21091), .Q (signal_21092) ) ;
    buf_clk cell_16210 ( .C (clk), .D (signal_21097), .Q (signal_21098) ) ;
    buf_clk cell_16216 ( .C (clk), .D (signal_21103), .Q (signal_21104) ) ;
    buf_clk cell_16222 ( .C (clk), .D (signal_21109), .Q (signal_21110) ) ;
    buf_clk cell_16228 ( .C (clk), .D (signal_21115), .Q (signal_21116) ) ;
    buf_clk cell_16234 ( .C (clk), .D (signal_21121), .Q (signal_21122) ) ;
    buf_clk cell_16240 ( .C (clk), .D (signal_21127), .Q (signal_21128) ) ;
    buf_clk cell_16246 ( .C (clk), .D (signal_21133), .Q (signal_21134) ) ;
    buf_clk cell_16252 ( .C (clk), .D (signal_21139), .Q (signal_21140) ) ;
    buf_clk cell_16258 ( .C (clk), .D (signal_21145), .Q (signal_21146) ) ;
    buf_clk cell_16264 ( .C (clk), .D (signal_21151), .Q (signal_21152) ) ;
    buf_clk cell_16270 ( .C (clk), .D (signal_21157), .Q (signal_21158) ) ;
    buf_clk cell_16276 ( .C (clk), .D (signal_21163), .Q (signal_21164) ) ;
    buf_clk cell_16282 ( .C (clk), .D (signal_21169), .Q (signal_21170) ) ;
    buf_clk cell_16288 ( .C (clk), .D (signal_21175), .Q (signal_21176) ) ;
    buf_clk cell_16294 ( .C (clk), .D (signal_21181), .Q (signal_21182) ) ;
    buf_clk cell_16300 ( .C (clk), .D (signal_21187), .Q (signal_21188) ) ;
    buf_clk cell_16306 ( .C (clk), .D (signal_21193), .Q (signal_21194) ) ;
    buf_clk cell_16312 ( .C (clk), .D (signal_21199), .Q (signal_21200) ) ;
    buf_clk cell_16318 ( .C (clk), .D (signal_21205), .Q (signal_21206) ) ;
    buf_clk cell_16324 ( .C (clk), .D (signal_21211), .Q (signal_21212) ) ;
    buf_clk cell_16330 ( .C (clk), .D (signal_21217), .Q (signal_21218) ) ;
    buf_clk cell_16336 ( .C (clk), .D (signal_21223), .Q (signal_21224) ) ;
    buf_clk cell_16342 ( .C (clk), .D (signal_21229), .Q (signal_21230) ) ;
    buf_clk cell_16348 ( .C (clk), .D (signal_21235), .Q (signal_21236) ) ;
    buf_clk cell_16354 ( .C (clk), .D (signal_21241), .Q (signal_21242) ) ;
    buf_clk cell_16360 ( .C (clk), .D (signal_21247), .Q (signal_21248) ) ;
    buf_clk cell_16366 ( .C (clk), .D (signal_21253), .Q (signal_21254) ) ;
    buf_clk cell_16372 ( .C (clk), .D (signal_21259), .Q (signal_21260) ) ;
    buf_clk cell_16378 ( .C (clk), .D (signal_21265), .Q (signal_21266) ) ;
    buf_clk cell_16384 ( .C (clk), .D (signal_21271), .Q (signal_21272) ) ;
    buf_clk cell_16390 ( .C (clk), .D (signal_21277), .Q (signal_21278) ) ;
    buf_clk cell_16396 ( .C (clk), .D (signal_21283), .Q (signal_21284) ) ;
    buf_clk cell_16402 ( .C (clk), .D (signal_21289), .Q (signal_21290) ) ;
    buf_clk cell_16408 ( .C (clk), .D (signal_21295), .Q (signal_21296) ) ;
    buf_clk cell_16414 ( .C (clk), .D (signal_21301), .Q (signal_21302) ) ;
    buf_clk cell_16420 ( .C (clk), .D (signal_21307), .Q (signal_21308) ) ;
    buf_clk cell_16426 ( .C (clk), .D (signal_21313), .Q (signal_21314) ) ;
    buf_clk cell_16432 ( .C (clk), .D (signal_21319), .Q (signal_21320) ) ;
    buf_clk cell_16438 ( .C (clk), .D (signal_21325), .Q (signal_21326) ) ;
    buf_clk cell_16444 ( .C (clk), .D (signal_21331), .Q (signal_21332) ) ;
    buf_clk cell_16450 ( .C (clk), .D (signal_21337), .Q (signal_21338) ) ;
    buf_clk cell_16456 ( .C (clk), .D (signal_21343), .Q (signal_21344) ) ;
    buf_clk cell_16462 ( .C (clk), .D (signal_21349), .Q (signal_21350) ) ;
    buf_clk cell_16468 ( .C (clk), .D (signal_21355), .Q (signal_21356) ) ;
    buf_clk cell_16474 ( .C (clk), .D (signal_21361), .Q (signal_21362) ) ;
    buf_clk cell_16480 ( .C (clk), .D (signal_21367), .Q (signal_21368) ) ;
    buf_clk cell_16486 ( .C (clk), .D (signal_21373), .Q (signal_21374) ) ;
    buf_clk cell_16492 ( .C (clk), .D (signal_21379), .Q (signal_21380) ) ;
    buf_clk cell_16498 ( .C (clk), .D (signal_21385), .Q (signal_21386) ) ;
    buf_clk cell_16504 ( .C (clk), .D (signal_21391), .Q (signal_21392) ) ;
    buf_clk cell_16510 ( .C (clk), .D (signal_21397), .Q (signal_21398) ) ;
    buf_clk cell_16516 ( .C (clk), .D (signal_21403), .Q (signal_21404) ) ;
    buf_clk cell_16522 ( .C (clk), .D (signal_21409), .Q (signal_21410) ) ;
    buf_clk cell_16528 ( .C (clk), .D (signal_21415), .Q (signal_21416) ) ;
    buf_clk cell_16534 ( .C (clk), .D (signal_21421), .Q (signal_21422) ) ;
    buf_clk cell_16540 ( .C (clk), .D (signal_21427), .Q (signal_21428) ) ;
    buf_clk cell_16546 ( .C (clk), .D (signal_21433), .Q (signal_21434) ) ;
    buf_clk cell_16552 ( .C (clk), .D (signal_21439), .Q (signal_21440) ) ;
    buf_clk cell_16558 ( .C (clk), .D (signal_21445), .Q (signal_21446) ) ;
    buf_clk cell_16564 ( .C (clk), .D (signal_21451), .Q (signal_21452) ) ;
    buf_clk cell_16570 ( .C (clk), .D (signal_21457), .Q (signal_21458) ) ;
    buf_clk cell_16576 ( .C (clk), .D (signal_21463), .Q (signal_21464) ) ;
    buf_clk cell_16582 ( .C (clk), .D (signal_21469), .Q (signal_21470) ) ;
    buf_clk cell_16588 ( .C (clk), .D (signal_21475), .Q (signal_21476) ) ;
    buf_clk cell_16594 ( .C (clk), .D (signal_21481), .Q (signal_21482) ) ;
    buf_clk cell_16600 ( .C (clk), .D (signal_21487), .Q (signal_21488) ) ;
    buf_clk cell_16606 ( .C (clk), .D (signal_21493), .Q (signal_21494) ) ;
    buf_clk cell_16612 ( .C (clk), .D (signal_21499), .Q (signal_21500) ) ;
    buf_clk cell_16618 ( .C (clk), .D (signal_21505), .Q (signal_21506) ) ;
    buf_clk cell_16624 ( .C (clk), .D (signal_21511), .Q (signal_21512) ) ;
    buf_clk cell_16630 ( .C (clk), .D (signal_21517), .Q (signal_21518) ) ;
    buf_clk cell_16636 ( .C (clk), .D (signal_21523), .Q (signal_21524) ) ;
    buf_clk cell_16642 ( .C (clk), .D (signal_21529), .Q (signal_21530) ) ;
    buf_clk cell_16648 ( .C (clk), .D (signal_21535), .Q (signal_21536) ) ;
    buf_clk cell_16654 ( .C (clk), .D (signal_21541), .Q (signal_21542) ) ;
    buf_clk cell_16660 ( .C (clk), .D (signal_21547), .Q (signal_21548) ) ;
    buf_clk cell_16666 ( .C (clk), .D (signal_21553), .Q (signal_21554) ) ;
    buf_clk cell_16672 ( .C (clk), .D (signal_21559), .Q (signal_21560) ) ;
    buf_clk cell_16678 ( .C (clk), .D (signal_21565), .Q (signal_21566) ) ;
    buf_clk cell_16684 ( .C (clk), .D (signal_21571), .Q (signal_21572) ) ;
    buf_clk cell_16690 ( .C (clk), .D (signal_21577), .Q (signal_21578) ) ;
    buf_clk cell_16696 ( .C (clk), .D (signal_21583), .Q (signal_21584) ) ;
    buf_clk cell_16702 ( .C (clk), .D (signal_21589), .Q (signal_21590) ) ;
    buf_clk cell_16708 ( .C (clk), .D (signal_21595), .Q (signal_21596) ) ;
    buf_clk cell_16714 ( .C (clk), .D (signal_21601), .Q (signal_21602) ) ;
    buf_clk cell_16720 ( .C (clk), .D (signal_21607), .Q (signal_21608) ) ;
    buf_clk cell_16726 ( .C (clk), .D (signal_21613), .Q (signal_21614) ) ;
    buf_clk cell_16732 ( .C (clk), .D (signal_21619), .Q (signal_21620) ) ;
    buf_clk cell_16738 ( .C (clk), .D (signal_21625), .Q (signal_21626) ) ;
    buf_clk cell_16744 ( .C (clk), .D (signal_21631), .Q (signal_21632) ) ;
    buf_clk cell_16750 ( .C (clk), .D (signal_21637), .Q (signal_21638) ) ;
    buf_clk cell_16756 ( .C (clk), .D (signal_21643), .Q (signal_21644) ) ;
    buf_clk cell_16762 ( .C (clk), .D (signal_21649), .Q (signal_21650) ) ;
    buf_clk cell_16768 ( .C (clk), .D (signal_21655), .Q (signal_21656) ) ;
    buf_clk cell_16774 ( .C (clk), .D (signal_21661), .Q (signal_21662) ) ;
    buf_clk cell_16780 ( .C (clk), .D (signal_21667), .Q (signal_21668) ) ;
    buf_clk cell_16786 ( .C (clk), .D (signal_21673), .Q (signal_21674) ) ;
    buf_clk cell_16792 ( .C (clk), .D (signal_21679), .Q (signal_21680) ) ;
    buf_clk cell_16798 ( .C (clk), .D (signal_21685), .Q (signal_21686) ) ;
    buf_clk cell_16804 ( .C (clk), .D (signal_21691), .Q (signal_21692) ) ;
    buf_clk cell_16810 ( .C (clk), .D (signal_21697), .Q (signal_21698) ) ;
    buf_clk cell_16816 ( .C (clk), .D (signal_21703), .Q (signal_21704) ) ;
    buf_clk cell_16822 ( .C (clk), .D (signal_21709), .Q (signal_21710) ) ;
    buf_clk cell_16828 ( .C (clk), .D (signal_21715), .Q (signal_21716) ) ;
    buf_clk cell_16834 ( .C (clk), .D (signal_21721), .Q (signal_21722) ) ;
    buf_clk cell_16840 ( .C (clk), .D (signal_21727), .Q (signal_21728) ) ;
    buf_clk cell_16846 ( .C (clk), .D (signal_21733), .Q (signal_21734) ) ;
    buf_clk cell_16852 ( .C (clk), .D (signal_21739), .Q (signal_21740) ) ;
    buf_clk cell_16858 ( .C (clk), .D (signal_21745), .Q (signal_21746) ) ;
    buf_clk cell_16864 ( .C (clk), .D (signal_21751), .Q (signal_21752) ) ;
    buf_clk cell_16870 ( .C (clk), .D (signal_21757), .Q (signal_21758) ) ;
    buf_clk cell_16876 ( .C (clk), .D (signal_21763), .Q (signal_21764) ) ;
    buf_clk cell_16882 ( .C (clk), .D (signal_21769), .Q (signal_21770) ) ;
    buf_clk cell_16888 ( .C (clk), .D (signal_21775), .Q (signal_21776) ) ;
    buf_clk cell_16894 ( .C (clk), .D (signal_21781), .Q (signal_21782) ) ;
    buf_clk cell_16900 ( .C (clk), .D (signal_21787), .Q (signal_21788) ) ;
    buf_clk cell_16906 ( .C (clk), .D (signal_21793), .Q (signal_21794) ) ;
    buf_clk cell_16912 ( .C (clk), .D (signal_21799), .Q (signal_21800) ) ;
    buf_clk cell_16918 ( .C (clk), .D (signal_21805), .Q (signal_21806) ) ;
    buf_clk cell_16924 ( .C (clk), .D (signal_21811), .Q (signal_21812) ) ;
    buf_clk cell_16930 ( .C (clk), .D (signal_21817), .Q (signal_21818) ) ;
    buf_clk cell_16936 ( .C (clk), .D (signal_21823), .Q (signal_21824) ) ;
    buf_clk cell_16942 ( .C (clk), .D (signal_21829), .Q (signal_21830) ) ;
    buf_clk cell_16948 ( .C (clk), .D (signal_21835), .Q (signal_21836) ) ;
    buf_clk cell_16954 ( .C (clk), .D (signal_21841), .Q (signal_21842) ) ;
    buf_clk cell_16960 ( .C (clk), .D (signal_21847), .Q (signal_21848) ) ;
    buf_clk cell_16966 ( .C (clk), .D (signal_21853), .Q (signal_21854) ) ;
    buf_clk cell_16972 ( .C (clk), .D (signal_21859), .Q (signal_21860) ) ;
    buf_clk cell_16978 ( .C (clk), .D (signal_21865), .Q (signal_21866) ) ;
    buf_clk cell_16984 ( .C (clk), .D (signal_21871), .Q (signal_21872) ) ;
    buf_clk cell_16990 ( .C (clk), .D (signal_21877), .Q (signal_21878) ) ;
    buf_clk cell_16996 ( .C (clk), .D (signal_21883), .Q (signal_21884) ) ;
    buf_clk cell_17002 ( .C (clk), .D (signal_21889), .Q (signal_21890) ) ;
    buf_clk cell_17008 ( .C (clk), .D (signal_21895), .Q (signal_21896) ) ;
    buf_clk cell_17014 ( .C (clk), .D (signal_21901), .Q (signal_21902) ) ;
    buf_clk cell_17020 ( .C (clk), .D (signal_21907), .Q (signal_21908) ) ;
    buf_clk cell_17026 ( .C (clk), .D (signal_21913), .Q (signal_21914) ) ;
    buf_clk cell_17032 ( .C (clk), .D (signal_21919), .Q (signal_21920) ) ;
    buf_clk cell_17038 ( .C (clk), .D (signal_21925), .Q (signal_21926) ) ;
    buf_clk cell_17044 ( .C (clk), .D (signal_21931), .Q (signal_21932) ) ;
    buf_clk cell_17050 ( .C (clk), .D (signal_21937), .Q (signal_21938) ) ;
    buf_clk cell_17056 ( .C (clk), .D (signal_21943), .Q (signal_21944) ) ;
    buf_clk cell_17062 ( .C (clk), .D (signal_21949), .Q (signal_21950) ) ;
    buf_clk cell_17068 ( .C (clk), .D (signal_21955), .Q (signal_21956) ) ;
    buf_clk cell_17074 ( .C (clk), .D (signal_21961), .Q (signal_21962) ) ;
    buf_clk cell_17080 ( .C (clk), .D (signal_21967), .Q (signal_21968) ) ;
    buf_clk cell_17086 ( .C (clk), .D (signal_21973), .Q (signal_21974) ) ;
    buf_clk cell_17092 ( .C (clk), .D (signal_21979), .Q (signal_21980) ) ;
    buf_clk cell_17098 ( .C (clk), .D (signal_21985), .Q (signal_21986) ) ;
    buf_clk cell_17104 ( .C (clk), .D (signal_21991), .Q (signal_21992) ) ;
    buf_clk cell_17110 ( .C (clk), .D (signal_21997), .Q (signal_21998) ) ;
    buf_clk cell_17116 ( .C (clk), .D (signal_22003), .Q (signal_22004) ) ;
    buf_clk cell_17122 ( .C (clk), .D (signal_22009), .Q (signal_22010) ) ;
    buf_clk cell_17128 ( .C (clk), .D (signal_22015), .Q (signal_22016) ) ;
    buf_clk cell_17134 ( .C (clk), .D (signal_22021), .Q (signal_22022) ) ;
    buf_clk cell_17140 ( .C (clk), .D (signal_22027), .Q (signal_22028) ) ;
    buf_clk cell_17146 ( .C (clk), .D (signal_22033), .Q (signal_22034) ) ;
    buf_clk cell_17152 ( .C (clk), .D (signal_22039), .Q (signal_22040) ) ;
    buf_clk cell_17158 ( .C (clk), .D (signal_22045), .Q (signal_22046) ) ;
    buf_clk cell_17164 ( .C (clk), .D (signal_22051), .Q (signal_22052) ) ;
    buf_clk cell_17170 ( .C (clk), .D (signal_22057), .Q (signal_22058) ) ;
    buf_clk cell_17176 ( .C (clk), .D (signal_22063), .Q (signal_22064) ) ;
    buf_clk cell_17182 ( .C (clk), .D (signal_22069), .Q (signal_22070) ) ;
    buf_clk cell_17188 ( .C (clk), .D (signal_22075), .Q (signal_22076) ) ;
    buf_clk cell_17194 ( .C (clk), .D (signal_22081), .Q (signal_22082) ) ;
    buf_clk cell_17200 ( .C (clk), .D (signal_22087), .Q (signal_22088) ) ;
    buf_clk cell_17206 ( .C (clk), .D (signal_22093), .Q (signal_22094) ) ;
    buf_clk cell_17212 ( .C (clk), .D (signal_22099), .Q (signal_22100) ) ;
    buf_clk cell_17218 ( .C (clk), .D (signal_22105), .Q (signal_22106) ) ;
    buf_clk cell_17224 ( .C (clk), .D (signal_22111), .Q (signal_22112) ) ;
    buf_clk cell_17230 ( .C (clk), .D (signal_22117), .Q (signal_22118) ) ;
    buf_clk cell_17236 ( .C (clk), .D (signal_22123), .Q (signal_22124) ) ;
    buf_clk cell_17242 ( .C (clk), .D (signal_22129), .Q (signal_22130) ) ;
    buf_clk cell_17248 ( .C (clk), .D (signal_22135), .Q (signal_22136) ) ;
    buf_clk cell_17254 ( .C (clk), .D (signal_22141), .Q (signal_22142) ) ;
    buf_clk cell_17260 ( .C (clk), .D (signal_22147), .Q (signal_22148) ) ;
    buf_clk cell_17266 ( .C (clk), .D (signal_22153), .Q (signal_22154) ) ;
    buf_clk cell_17272 ( .C (clk), .D (signal_22159), .Q (signal_22160) ) ;
    buf_clk cell_17278 ( .C (clk), .D (signal_22165), .Q (signal_22166) ) ;
    buf_clk cell_17284 ( .C (clk), .D (signal_22171), .Q (signal_22172) ) ;
    buf_clk cell_17290 ( .C (clk), .D (signal_22177), .Q (signal_22178) ) ;
    buf_clk cell_17296 ( .C (clk), .D (signal_22183), .Q (signal_22184) ) ;
    buf_clk cell_17302 ( .C (clk), .D (signal_22189), .Q (signal_22190) ) ;
    buf_clk cell_17308 ( .C (clk), .D (signal_22195), .Q (signal_22196) ) ;
    buf_clk cell_17314 ( .C (clk), .D (signal_22201), .Q (signal_22202) ) ;
    buf_clk cell_17320 ( .C (clk), .D (signal_22207), .Q (signal_22208) ) ;
    buf_clk cell_17326 ( .C (clk), .D (signal_22213), .Q (signal_22214) ) ;
    buf_clk cell_17332 ( .C (clk), .D (signal_22219), .Q (signal_22220) ) ;
    buf_clk cell_17338 ( .C (clk), .D (signal_22225), .Q (signal_22226) ) ;
    buf_clk cell_17344 ( .C (clk), .D (signal_22231), .Q (signal_22232) ) ;
    buf_clk cell_17350 ( .C (clk), .D (signal_22237), .Q (signal_22238) ) ;
    buf_clk cell_17356 ( .C (clk), .D (signal_22243), .Q (signal_22244) ) ;
    buf_clk cell_17362 ( .C (clk), .D (signal_22249), .Q (signal_22250) ) ;
    buf_clk cell_17368 ( .C (clk), .D (signal_22255), .Q (signal_22256) ) ;
    buf_clk cell_17374 ( .C (clk), .D (signal_22261), .Q (signal_22262) ) ;
    buf_clk cell_17380 ( .C (clk), .D (signal_22267), .Q (signal_22268) ) ;
    buf_clk cell_17386 ( .C (clk), .D (signal_22273), .Q (signal_22274) ) ;
    buf_clk cell_17392 ( .C (clk), .D (signal_22279), .Q (signal_22280) ) ;
    buf_clk cell_17398 ( .C (clk), .D (signal_22285), .Q (signal_22286) ) ;
    buf_clk cell_17404 ( .C (clk), .D (signal_22291), .Q (signal_22292) ) ;
    buf_clk cell_17410 ( .C (clk), .D (signal_22297), .Q (signal_22298) ) ;
    buf_clk cell_17416 ( .C (clk), .D (signal_22303), .Q (signal_22304) ) ;
    buf_clk cell_17422 ( .C (clk), .D (signal_22309), .Q (signal_22310) ) ;
    buf_clk cell_17428 ( .C (clk), .D (signal_22315), .Q (signal_22316) ) ;
    buf_clk cell_17434 ( .C (clk), .D (signal_22321), .Q (signal_22322) ) ;
    buf_clk cell_17440 ( .C (clk), .D (signal_22327), .Q (signal_22328) ) ;
    buf_clk cell_17446 ( .C (clk), .D (signal_22333), .Q (signal_22334) ) ;
    buf_clk cell_17452 ( .C (clk), .D (signal_22339), .Q (signal_22340) ) ;
    buf_clk cell_17458 ( .C (clk), .D (signal_22345), .Q (signal_22346) ) ;
    buf_clk cell_17464 ( .C (clk), .D (signal_22351), .Q (signal_22352) ) ;
    buf_clk cell_17470 ( .C (clk), .D (signal_22357), .Q (signal_22358) ) ;
    buf_clk cell_17476 ( .C (clk), .D (signal_22363), .Q (signal_22364) ) ;
    buf_clk cell_17482 ( .C (clk), .D (signal_22369), .Q (signal_22370) ) ;
    buf_clk cell_17488 ( .C (clk), .D (signal_22375), .Q (signal_22376) ) ;
    buf_clk cell_17494 ( .C (clk), .D (signal_22381), .Q (signal_22382) ) ;
    buf_clk cell_17500 ( .C (clk), .D (signal_22387), .Q (signal_22388) ) ;
    buf_clk cell_17506 ( .C (clk), .D (signal_22393), .Q (signal_22394) ) ;
    buf_clk cell_17512 ( .C (clk), .D (signal_22399), .Q (signal_22400) ) ;
    buf_clk cell_17518 ( .C (clk), .D (signal_22405), .Q (signal_22406) ) ;
    buf_clk cell_17524 ( .C (clk), .D (signal_22411), .Q (signal_22412) ) ;
    buf_clk cell_17530 ( .C (clk), .D (signal_22417), .Q (signal_22418) ) ;
    buf_clk cell_17536 ( .C (clk), .D (signal_22423), .Q (signal_22424) ) ;
    buf_clk cell_17542 ( .C (clk), .D (signal_22429), .Q (signal_22430) ) ;
    buf_clk cell_17548 ( .C (clk), .D (signal_22435), .Q (signal_22436) ) ;
    buf_clk cell_17554 ( .C (clk), .D (signal_22441), .Q (signal_22442) ) ;
    buf_clk cell_17560 ( .C (clk), .D (signal_22447), .Q (signal_22448) ) ;
    buf_clk cell_17566 ( .C (clk), .D (signal_22453), .Q (signal_22454) ) ;
    buf_clk cell_17572 ( .C (clk), .D (signal_22459), .Q (signal_22460) ) ;
    buf_clk cell_17578 ( .C (clk), .D (signal_22465), .Q (signal_22466) ) ;
    buf_clk cell_17584 ( .C (clk), .D (signal_22471), .Q (signal_22472) ) ;
    buf_clk cell_17590 ( .C (clk), .D (signal_22477), .Q (signal_22478) ) ;
    buf_clk cell_17598 ( .C (clk), .D (signal_22485), .Q (signal_22486) ) ;
    buf_clk cell_17606 ( .C (clk), .D (signal_22493), .Q (signal_22494) ) ;
    buf_clk cell_17614 ( .C (clk), .D (signal_22501), .Q (signal_22502) ) ;
    buf_clk cell_17622 ( .C (clk), .D (signal_22509), .Q (signal_22510) ) ;
    buf_clk cell_17630 ( .C (clk), .D (signal_22517), .Q (signal_22518) ) ;
    buf_clk cell_17638 ( .C (clk), .D (signal_22525), .Q (signal_22526) ) ;
    buf_clk cell_17646 ( .C (clk), .D (signal_22533), .Q (signal_22534) ) ;
    buf_clk cell_17654 ( .C (clk), .D (signal_22541), .Q (signal_22542) ) ;
    buf_clk cell_17662 ( .C (clk), .D (signal_22549), .Q (signal_22550) ) ;
    buf_clk cell_17670 ( .C (clk), .D (signal_22557), .Q (signal_22558) ) ;
    buf_clk cell_17678 ( .C (clk), .D (signal_22565), .Q (signal_22566) ) ;
    buf_clk cell_17686 ( .C (clk), .D (signal_22573), .Q (signal_22574) ) ;
    buf_clk cell_17694 ( .C (clk), .D (signal_22581), .Q (signal_22582) ) ;
    buf_clk cell_17702 ( .C (clk), .D (signal_22589), .Q (signal_22590) ) ;
    buf_clk cell_17710 ( .C (clk), .D (signal_22597), .Q (signal_22598) ) ;
    buf_clk cell_17718 ( .C (clk), .D (signal_22605), .Q (signal_22606) ) ;
    buf_clk cell_17726 ( .C (clk), .D (signal_22613), .Q (signal_22614) ) ;
    buf_clk cell_17734 ( .C (clk), .D (signal_22621), .Q (signal_22622) ) ;
    buf_clk cell_17742 ( .C (clk), .D (signal_22629), .Q (signal_22630) ) ;
    buf_clk cell_17750 ( .C (clk), .D (signal_22637), .Q (signal_22638) ) ;
    buf_clk cell_17758 ( .C (clk), .D (signal_22645), .Q (signal_22646) ) ;
    buf_clk cell_17766 ( .C (clk), .D (signal_22653), .Q (signal_22654) ) ;
    buf_clk cell_17774 ( .C (clk), .D (signal_22661), .Q (signal_22662) ) ;
    buf_clk cell_17782 ( .C (clk), .D (signal_22669), .Q (signal_22670) ) ;
    buf_clk cell_17790 ( .C (clk), .D (signal_22677), .Q (signal_22678) ) ;
    buf_clk cell_17798 ( .C (clk), .D (signal_22685), .Q (signal_22686) ) ;
    buf_clk cell_17806 ( .C (clk), .D (signal_22693), .Q (signal_22694) ) ;
    buf_clk cell_17814 ( .C (clk), .D (signal_22701), .Q (signal_22702) ) ;
    buf_clk cell_17822 ( .C (clk), .D (signal_22709), .Q (signal_22710) ) ;
    buf_clk cell_17830 ( .C (clk), .D (signal_22717), .Q (signal_22718) ) ;
    buf_clk cell_17838 ( .C (clk), .D (signal_22725), .Q (signal_22726) ) ;
    buf_clk cell_17846 ( .C (clk), .D (signal_22733), .Q (signal_22734) ) ;
    buf_clk cell_17854 ( .C (clk), .D (signal_22741), .Q (signal_22742) ) ;
    buf_clk cell_17862 ( .C (clk), .D (signal_22749), .Q (signal_22750) ) ;
    buf_clk cell_17870 ( .C (clk), .D (signal_22757), .Q (signal_22758) ) ;
    buf_clk cell_17878 ( .C (clk), .D (signal_22765), .Q (signal_22766) ) ;
    buf_clk cell_17886 ( .C (clk), .D (signal_22773), .Q (signal_22774) ) ;
    buf_clk cell_17894 ( .C (clk), .D (signal_22781), .Q (signal_22782) ) ;
    buf_clk cell_17902 ( .C (clk), .D (signal_22789), .Q (signal_22790) ) ;
    buf_clk cell_17910 ( .C (clk), .D (signal_22797), .Q (signal_22798) ) ;
    buf_clk cell_17918 ( .C (clk), .D (signal_22805), .Q (signal_22806) ) ;
    buf_clk cell_17926 ( .C (clk), .D (signal_22813), .Q (signal_22814) ) ;
    buf_clk cell_17934 ( .C (clk), .D (signal_22821), .Q (signal_22822) ) ;
    buf_clk cell_17942 ( .C (clk), .D (signal_22829), .Q (signal_22830) ) ;
    buf_clk cell_17950 ( .C (clk), .D (signal_22837), .Q (signal_22838) ) ;
    buf_clk cell_17958 ( .C (clk), .D (signal_22845), .Q (signal_22846) ) ;
    buf_clk cell_17966 ( .C (clk), .D (signal_22853), .Q (signal_22854) ) ;
    buf_clk cell_17974 ( .C (clk), .D (signal_22861), .Q (signal_22862) ) ;
    buf_clk cell_17982 ( .C (clk), .D (signal_22869), .Q (signal_22870) ) ;
    buf_clk cell_17990 ( .C (clk), .D (signal_22877), .Q (signal_22878) ) ;
    buf_clk cell_17998 ( .C (clk), .D (signal_22885), .Q (signal_22886) ) ;
    buf_clk cell_18006 ( .C (clk), .D (signal_22893), .Q (signal_22894) ) ;
    buf_clk cell_18014 ( .C (clk), .D (signal_22901), .Q (signal_22902) ) ;
    buf_clk cell_18022 ( .C (clk), .D (signal_22909), .Q (signal_22910) ) ;
    buf_clk cell_18030 ( .C (clk), .D (signal_22917), .Q (signal_22918) ) ;
    buf_clk cell_18038 ( .C (clk), .D (signal_22925), .Q (signal_22926) ) ;
    buf_clk cell_18046 ( .C (clk), .D (signal_22933), .Q (signal_22934) ) ;
    buf_clk cell_18054 ( .C (clk), .D (signal_22941), .Q (signal_22942) ) ;
    buf_clk cell_18062 ( .C (clk), .D (signal_22949), .Q (signal_22950) ) ;
    buf_clk cell_18070 ( .C (clk), .D (signal_22957), .Q (signal_22958) ) ;
    buf_clk cell_18078 ( .C (clk), .D (signal_22965), .Q (signal_22966) ) ;
    buf_clk cell_18086 ( .C (clk), .D (signal_22973), .Q (signal_22974) ) ;
    buf_clk cell_18094 ( .C (clk), .D (signal_22981), .Q (signal_22982) ) ;
    buf_clk cell_18102 ( .C (clk), .D (signal_22989), .Q (signal_22990) ) ;
    buf_clk cell_18110 ( .C (clk), .D (signal_22997), .Q (signal_22998) ) ;
    buf_clk cell_18118 ( .C (clk), .D (signal_23005), .Q (signal_23006) ) ;
    buf_clk cell_18126 ( .C (clk), .D (signal_23013), .Q (signal_23014) ) ;
    buf_clk cell_18134 ( .C (clk), .D (signal_23021), .Q (signal_23022) ) ;
    buf_clk cell_18142 ( .C (clk), .D (signal_23029), .Q (signal_23030) ) ;
    buf_clk cell_18150 ( .C (clk), .D (signal_23037), .Q (signal_23038) ) ;
    buf_clk cell_18158 ( .C (clk), .D (signal_23045), .Q (signal_23046) ) ;
    buf_clk cell_18166 ( .C (clk), .D (signal_23053), .Q (signal_23054) ) ;
    buf_clk cell_18174 ( .C (clk), .D (signal_23061), .Q (signal_23062) ) ;
    buf_clk cell_18182 ( .C (clk), .D (signal_23069), .Q (signal_23070) ) ;
    buf_clk cell_18190 ( .C (clk), .D (signal_23077), .Q (signal_23078) ) ;
    buf_clk cell_18198 ( .C (clk), .D (signal_23085), .Q (signal_23086) ) ;
    buf_clk cell_18206 ( .C (clk), .D (signal_23093), .Q (signal_23094) ) ;
    buf_clk cell_18214 ( .C (clk), .D (signal_23101), .Q (signal_23102) ) ;
    buf_clk cell_18222 ( .C (clk), .D (signal_23109), .Q (signal_23110) ) ;
    buf_clk cell_18230 ( .C (clk), .D (signal_23117), .Q (signal_23118) ) ;
    buf_clk cell_18238 ( .C (clk), .D (signal_23125), .Q (signal_23126) ) ;
    buf_clk cell_18246 ( .C (clk), .D (signal_23133), .Q (signal_23134) ) ;
    buf_clk cell_18254 ( .C (clk), .D (signal_23141), .Q (signal_23142) ) ;
    buf_clk cell_18262 ( .C (clk), .D (signal_23149), .Q (signal_23150) ) ;
    buf_clk cell_18270 ( .C (clk), .D (signal_23157), .Q (signal_23158) ) ;
    buf_clk cell_18278 ( .C (clk), .D (signal_23165), .Q (signal_23166) ) ;
    buf_clk cell_18286 ( .C (clk), .D (signal_23173), .Q (signal_23174) ) ;
    buf_clk cell_18294 ( .C (clk), .D (signal_23181), .Q (signal_23182) ) ;
    buf_clk cell_18302 ( .C (clk), .D (signal_23189), .Q (signal_23190) ) ;
    buf_clk cell_18310 ( .C (clk), .D (signal_23197), .Q (signal_23198) ) ;
    buf_clk cell_18318 ( .C (clk), .D (signal_23205), .Q (signal_23206) ) ;
    buf_clk cell_18326 ( .C (clk), .D (signal_23213), .Q (signal_23214) ) ;
    buf_clk cell_18334 ( .C (clk), .D (signal_23221), .Q (signal_23222) ) ;
    buf_clk cell_18342 ( .C (clk), .D (signal_23229), .Q (signal_23230) ) ;
    buf_clk cell_18350 ( .C (clk), .D (signal_23237), .Q (signal_23238) ) ;
    buf_clk cell_18358 ( .C (clk), .D (signal_23245), .Q (signal_23246) ) ;
    buf_clk cell_18366 ( .C (clk), .D (signal_23253), .Q (signal_23254) ) ;
    buf_clk cell_18374 ( .C (clk), .D (signal_23261), .Q (signal_23262) ) ;
    buf_clk cell_18382 ( .C (clk), .D (signal_23269), .Q (signal_23270) ) ;
    buf_clk cell_18390 ( .C (clk), .D (signal_23277), .Q (signal_23278) ) ;
    buf_clk cell_18398 ( .C (clk), .D (signal_23285), .Q (signal_23286) ) ;
    buf_clk cell_18410 ( .C (clk), .D (signal_23297), .Q (signal_23298) ) ;
    buf_clk cell_18418 ( .C (clk), .D (signal_23305), .Q (signal_23306) ) ;
    buf_clk cell_18426 ( .C (clk), .D (signal_23313), .Q (signal_23314) ) ;
    buf_clk cell_18434 ( .C (clk), .D (signal_23321), .Q (signal_23322) ) ;
    buf_clk cell_18442 ( .C (clk), .D (signal_23329), .Q (signal_23330) ) ;
    buf_clk cell_18450 ( .C (clk), .D (signal_23337), .Q (signal_23338) ) ;
    buf_clk cell_18458 ( .C (clk), .D (signal_23345), .Q (signal_23346) ) ;
    buf_clk cell_18466 ( .C (clk), .D (signal_23353), .Q (signal_23354) ) ;
    buf_clk cell_18474 ( .C (clk), .D (signal_23361), .Q (signal_23362) ) ;
    buf_clk cell_18482 ( .C (clk), .D (signal_23369), .Q (signal_23370) ) ;
    buf_clk cell_18490 ( .C (clk), .D (signal_23377), .Q (signal_23378) ) ;
    buf_clk cell_18498 ( .C (clk), .D (signal_23385), .Q (signal_23386) ) ;
    buf_clk cell_18506 ( .C (clk), .D (signal_23393), .Q (signal_23394) ) ;
    buf_clk cell_18514 ( .C (clk), .D (signal_23401), .Q (signal_23402) ) ;
    buf_clk cell_18522 ( .C (clk), .D (signal_23409), .Q (signal_23410) ) ;
    buf_clk cell_18530 ( .C (clk), .D (signal_23417), .Q (signal_23418) ) ;
    buf_clk cell_18538 ( .C (clk), .D (signal_23425), .Q (signal_23426) ) ;
    buf_clk cell_18546 ( .C (clk), .D (signal_23433), .Q (signal_23434) ) ;
    buf_clk cell_18554 ( .C (clk), .D (signal_23441), .Q (signal_23442) ) ;
    buf_clk cell_18562 ( .C (clk), .D (signal_23449), .Q (signal_23450) ) ;
    buf_clk cell_18570 ( .C (clk), .D (signal_23457), .Q (signal_23458) ) ;
    buf_clk cell_18578 ( .C (clk), .D (signal_23465), .Q (signal_23466) ) ;
    buf_clk cell_18586 ( .C (clk), .D (signal_23473), .Q (signal_23474) ) ;
    buf_clk cell_18594 ( .C (clk), .D (signal_23481), .Q (signal_23482) ) ;
    buf_clk cell_18602 ( .C (clk), .D (signal_23489), .Q (signal_23490) ) ;
    buf_clk cell_18610 ( .C (clk), .D (signal_23497), .Q (signal_23498) ) ;
    buf_clk cell_18618 ( .C (clk), .D (signal_23505), .Q (signal_23506) ) ;
    buf_clk cell_18626 ( .C (clk), .D (signal_23513), .Q (signal_23514) ) ;
    buf_clk cell_18634 ( .C (clk), .D (signal_23521), .Q (signal_23522) ) ;
    buf_clk cell_18642 ( .C (clk), .D (signal_23529), .Q (signal_23530) ) ;
    buf_clk cell_18654 ( .C (clk), .D (signal_23541), .Q (signal_23542) ) ;
    buf_clk cell_18662 ( .C (clk), .D (signal_23549), .Q (signal_23550) ) ;
    buf_clk cell_18670 ( .C (clk), .D (signal_23557), .Q (signal_23558) ) ;
    buf_clk cell_18678 ( .C (clk), .D (signal_23565), .Q (signal_23566) ) ;
    buf_clk cell_18686 ( .C (clk), .D (signal_23573), .Q (signal_23574) ) ;
    buf_clk cell_18694 ( .C (clk), .D (signal_23581), .Q (signal_23582) ) ;
    buf_clk cell_18702 ( .C (clk), .D (signal_23589), .Q (signal_23590) ) ;
    buf_clk cell_18710 ( .C (clk), .D (signal_23597), .Q (signal_23598) ) ;
    buf_clk cell_18718 ( .C (clk), .D (signal_23605), .Q (signal_23606) ) ;
    buf_clk cell_18726 ( .C (clk), .D (signal_23613), .Q (signal_23614) ) ;
    buf_clk cell_18734 ( .C (clk), .D (signal_23621), .Q (signal_23622) ) ;
    buf_clk cell_18742 ( .C (clk), .D (signal_23629), .Q (signal_23630) ) ;
    buf_clk cell_18754 ( .C (clk), .D (signal_23641), .Q (signal_23642) ) ;
    buf_clk cell_18762 ( .C (clk), .D (signal_23649), .Q (signal_23650) ) ;
    buf_clk cell_18770 ( .C (clk), .D (signal_23657), .Q (signal_23658) ) ;
    buf_clk cell_18778 ( .C (clk), .D (signal_23665), .Q (signal_23666) ) ;
    buf_clk cell_18786 ( .C (clk), .D (signal_23673), .Q (signal_23674) ) ;
    buf_clk cell_18794 ( .C (clk), .D (signal_23681), .Q (signal_23682) ) ;
    buf_clk cell_18802 ( .C (clk), .D (signal_23689), .Q (signal_23690) ) ;
    buf_clk cell_18810 ( .C (clk), .D (signal_23697), .Q (signal_23698) ) ;
    buf_clk cell_18818 ( .C (clk), .D (signal_23705), .Q (signal_23706) ) ;
    buf_clk cell_18826 ( .C (clk), .D (signal_23713), .Q (signal_23714) ) ;
    buf_clk cell_18834 ( .C (clk), .D (signal_23721), .Q (signal_23722) ) ;
    buf_clk cell_18842 ( .C (clk), .D (signal_23729), .Q (signal_23730) ) ;
    buf_clk cell_18850 ( .C (clk), .D (signal_23737), .Q (signal_23738) ) ;
    buf_clk cell_18858 ( .C (clk), .D (signal_23745), .Q (signal_23746) ) ;
    buf_clk cell_18866 ( .C (clk), .D (signal_23753), .Q (signal_23754) ) ;
    buf_clk cell_18874 ( .C (clk), .D (signal_23761), .Q (signal_23762) ) ;
    buf_clk cell_18882 ( .C (clk), .D (signal_23769), .Q (signal_23770) ) ;
    buf_clk cell_18890 ( .C (clk), .D (signal_23777), .Q (signal_23778) ) ;
    buf_clk cell_18898 ( .C (clk), .D (signal_23785), .Q (signal_23786) ) ;
    buf_clk cell_18906 ( .C (clk), .D (signal_23793), .Q (signal_23794) ) ;
    buf_clk cell_18914 ( .C (clk), .D (signal_23801), .Q (signal_23802) ) ;
    buf_clk cell_18922 ( .C (clk), .D (signal_23809), .Q (signal_23810) ) ;
    buf_clk cell_18930 ( .C (clk), .D (signal_23817), .Q (signal_23818) ) ;
    buf_clk cell_18938 ( .C (clk), .D (signal_23825), .Q (signal_23826) ) ;
    buf_clk cell_18946 ( .C (clk), .D (signal_23833), .Q (signal_23834) ) ;
    buf_clk cell_18954 ( .C (clk), .D (signal_23841), .Q (signal_23842) ) ;
    buf_clk cell_18962 ( .C (clk), .D (signal_23849), .Q (signal_23850) ) ;
    buf_clk cell_18970 ( .C (clk), .D (signal_23857), .Q (signal_23858) ) ;
    buf_clk cell_18978 ( .C (clk), .D (signal_23865), .Q (signal_23866) ) ;
    buf_clk cell_18986 ( .C (clk), .D (signal_23873), .Q (signal_23874) ) ;
    buf_clk cell_18994 ( .C (clk), .D (signal_23881), .Q (signal_23882) ) ;
    buf_clk cell_19002 ( .C (clk), .D (signal_23889), .Q (signal_23890) ) ;
    buf_clk cell_19010 ( .C (clk), .D (signal_23897), .Q (signal_23898) ) ;
    buf_clk cell_19018 ( .C (clk), .D (signal_23905), .Q (signal_23906) ) ;
    buf_clk cell_19026 ( .C (clk), .D (signal_23913), .Q (signal_23914) ) ;
    buf_clk cell_19034 ( .C (clk), .D (signal_23921), .Q (signal_23922) ) ;
    buf_clk cell_19042 ( .C (clk), .D (signal_23929), .Q (signal_23930) ) ;
    buf_clk cell_19050 ( .C (clk), .D (signal_23937), .Q (signal_23938) ) ;
    buf_clk cell_19058 ( .C (clk), .D (signal_23945), .Q (signal_23946) ) ;
    buf_clk cell_19066 ( .C (clk), .D (signal_23953), .Q (signal_23954) ) ;
    buf_clk cell_19074 ( .C (clk), .D (signal_23961), .Q (signal_23962) ) ;
    buf_clk cell_19082 ( .C (clk), .D (signal_23969), .Q (signal_23970) ) ;
    buf_clk cell_19090 ( .C (clk), .D (signal_23977), .Q (signal_23978) ) ;
    buf_clk cell_19098 ( .C (clk), .D (signal_23985), .Q (signal_23986) ) ;
    buf_clk cell_19106 ( .C (clk), .D (signal_23993), .Q (signal_23994) ) ;
    buf_clk cell_19114 ( .C (clk), .D (signal_24001), .Q (signal_24002) ) ;

    /* cells in depth 7 */
    buf_clk cell_8547 ( .C (clk), .D (signal_13434), .Q (signal_13435) ) ;
    buf_clk cell_8555 ( .C (clk), .D (signal_13442), .Q (signal_13443) ) ;
    buf_clk cell_8563 ( .C (clk), .D (signal_13450), .Q (signal_13451) ) ;
    buf_clk cell_8571 ( .C (clk), .D (signal_13458), .Q (signal_13459) ) ;
    buf_clk cell_8579 ( .C (clk), .D (signal_13466), .Q (signal_13467) ) ;
    buf_clk cell_8587 ( .C (clk), .D (signal_13474), .Q (signal_13475) ) ;
    buf_clk cell_8595 ( .C (clk), .D (signal_13482), .Q (signal_13483) ) ;
    buf_clk cell_8603 ( .C (clk), .D (signal_13490), .Q (signal_13491) ) ;
    buf_clk cell_8611 ( .C (clk), .D (signal_13498), .Q (signal_13499) ) ;
    buf_clk cell_8619 ( .C (clk), .D (signal_13506), .Q (signal_13507) ) ;
    buf_clk cell_8627 ( .C (clk), .D (signal_13514), .Q (signal_13515) ) ;
    buf_clk cell_8635 ( .C (clk), .D (signal_13522), .Q (signal_13523) ) ;
    buf_clk cell_8643 ( .C (clk), .D (signal_13530), .Q (signal_13531) ) ;
    buf_clk cell_8651 ( .C (clk), .D (signal_13538), .Q (signal_13539) ) ;
    buf_clk cell_8659 ( .C (clk), .D (signal_13546), .Q (signal_13547) ) ;
    buf_clk cell_8667 ( .C (clk), .D (signal_13554), .Q (signal_13555) ) ;
    buf_clk cell_8675 ( .C (clk), .D (signal_13562), .Q (signal_13563) ) ;
    buf_clk cell_8683 ( .C (clk), .D (signal_13570), .Q (signal_13571) ) ;
    buf_clk cell_8691 ( .C (clk), .D (signal_13578), .Q (signal_13579) ) ;
    buf_clk cell_8699 ( .C (clk), .D (signal_13586), .Q (signal_13587) ) ;
    buf_clk cell_8707 ( .C (clk), .D (signal_13594), .Q (signal_13595) ) ;
    buf_clk cell_8715 ( .C (clk), .D (signal_13602), .Q (signal_13603) ) ;
    buf_clk cell_8723 ( .C (clk), .D (signal_13610), .Q (signal_13611) ) ;
    buf_clk cell_8731 ( .C (clk), .D (signal_13618), .Q (signal_13619) ) ;
    buf_clk cell_8739 ( .C (clk), .D (signal_13626), .Q (signal_13627) ) ;
    buf_clk cell_8747 ( .C (clk), .D (signal_13634), .Q (signal_13635) ) ;
    buf_clk cell_8755 ( .C (clk), .D (signal_13642), .Q (signal_13643) ) ;
    buf_clk cell_8763 ( .C (clk), .D (signal_13650), .Q (signal_13651) ) ;
    buf_clk cell_8771 ( .C (clk), .D (signal_13658), .Q (signal_13659) ) ;
    buf_clk cell_8779 ( .C (clk), .D (signal_13666), .Q (signal_13667) ) ;
    buf_clk cell_8787 ( .C (clk), .D (signal_13674), .Q (signal_13675) ) ;
    buf_clk cell_8795 ( .C (clk), .D (signal_13682), .Q (signal_13683) ) ;
    buf_clk cell_8803 ( .C (clk), .D (signal_13690), .Q (signal_13691) ) ;
    buf_clk cell_8811 ( .C (clk), .D (signal_13698), .Q (signal_13699) ) ;
    buf_clk cell_8819 ( .C (clk), .D (signal_13706), .Q (signal_13707) ) ;
    buf_clk cell_8827 ( .C (clk), .D (signal_13714), .Q (signal_13715) ) ;
    buf_clk cell_8835 ( .C (clk), .D (signal_13722), .Q (signal_13723) ) ;
    buf_clk cell_8843 ( .C (clk), .D (signal_13730), .Q (signal_13731) ) ;
    buf_clk cell_8851 ( .C (clk), .D (signal_13738), .Q (signal_13739) ) ;
    buf_clk cell_8859 ( .C (clk), .D (signal_13746), .Q (signal_13747) ) ;
    buf_clk cell_8867 ( .C (clk), .D (signal_13754), .Q (signal_13755) ) ;
    buf_clk cell_8875 ( .C (clk), .D (signal_13762), .Q (signal_13763) ) ;
    buf_clk cell_8883 ( .C (clk), .D (signal_13770), .Q (signal_13771) ) ;
    buf_clk cell_8891 ( .C (clk), .D (signal_13778), .Q (signal_13779) ) ;
    buf_clk cell_8899 ( .C (clk), .D (signal_13786), .Q (signal_13787) ) ;
    buf_clk cell_8907 ( .C (clk), .D (signal_13794), .Q (signal_13795) ) ;
    buf_clk cell_8915 ( .C (clk), .D (signal_13802), .Q (signal_13803) ) ;
    buf_clk cell_8923 ( .C (clk), .D (signal_13810), .Q (signal_13811) ) ;
    buf_clk cell_8931 ( .C (clk), .D (signal_13818), .Q (signal_13819) ) ;
    buf_clk cell_8939 ( .C (clk), .D (signal_13826), .Q (signal_13827) ) ;
    buf_clk cell_8947 ( .C (clk), .D (signal_13834), .Q (signal_13835) ) ;
    buf_clk cell_8955 ( .C (clk), .D (signal_13842), .Q (signal_13843) ) ;
    buf_clk cell_8963 ( .C (clk), .D (signal_13850), .Q (signal_13851) ) ;
    buf_clk cell_8971 ( .C (clk), .D (signal_13858), .Q (signal_13859) ) ;
    buf_clk cell_8979 ( .C (clk), .D (signal_13866), .Q (signal_13867) ) ;
    buf_clk cell_8987 ( .C (clk), .D (signal_13874), .Q (signal_13875) ) ;
    buf_clk cell_8995 ( .C (clk), .D (signal_13882), .Q (signal_13883) ) ;
    buf_clk cell_9003 ( .C (clk), .D (signal_13890), .Q (signal_13891) ) ;
    buf_clk cell_9011 ( .C (clk), .D (signal_13898), .Q (signal_13899) ) ;
    buf_clk cell_9019 ( .C (clk), .D (signal_13906), .Q (signal_13907) ) ;
    buf_clk cell_9027 ( .C (clk), .D (signal_13914), .Q (signal_13915) ) ;
    buf_clk cell_9035 ( .C (clk), .D (signal_13922), .Q (signal_13923) ) ;
    buf_clk cell_9043 ( .C (clk), .D (signal_13930), .Q (signal_13931) ) ;
    buf_clk cell_9051 ( .C (clk), .D (signal_13938), .Q (signal_13939) ) ;
    buf_clk cell_9059 ( .C (clk), .D (signal_13946), .Q (signal_13947) ) ;
    buf_clk cell_9067 ( .C (clk), .D (signal_13954), .Q (signal_13955) ) ;
    buf_clk cell_9075 ( .C (clk), .D (signal_13962), .Q (signal_13963) ) ;
    buf_clk cell_9083 ( .C (clk), .D (signal_13970), .Q (signal_13971) ) ;
    buf_clk cell_9091 ( .C (clk), .D (signal_13978), .Q (signal_13979) ) ;
    buf_clk cell_9099 ( .C (clk), .D (signal_13986), .Q (signal_13987) ) ;
    buf_clk cell_9107 ( .C (clk), .D (signal_13994), .Q (signal_13995) ) ;
    buf_clk cell_9115 ( .C (clk), .D (signal_14002), .Q (signal_14003) ) ;
    buf_clk cell_9123 ( .C (clk), .D (signal_14010), .Q (signal_14011) ) ;
    buf_clk cell_9131 ( .C (clk), .D (signal_14018), .Q (signal_14019) ) ;
    buf_clk cell_9139 ( .C (clk), .D (signal_14026), .Q (signal_14027) ) ;
    buf_clk cell_9147 ( .C (clk), .D (signal_14034), .Q (signal_14035) ) ;
    buf_clk cell_9155 ( .C (clk), .D (signal_14042), .Q (signal_14043) ) ;
    buf_clk cell_9163 ( .C (clk), .D (signal_14050), .Q (signal_14051) ) ;
    buf_clk cell_9171 ( .C (clk), .D (signal_14058), .Q (signal_14059) ) ;
    buf_clk cell_9179 ( .C (clk), .D (signal_14066), .Q (signal_14067) ) ;
    buf_clk cell_9187 ( .C (clk), .D (signal_14074), .Q (signal_14075) ) ;
    buf_clk cell_9195 ( .C (clk), .D (signal_14082), .Q (signal_14083) ) ;
    buf_clk cell_9203 ( .C (clk), .D (signal_14090), .Q (signal_14091) ) ;
    buf_clk cell_9211 ( .C (clk), .D (signal_14098), .Q (signal_14099) ) ;
    buf_clk cell_9219 ( .C (clk), .D (signal_14106), .Q (signal_14107) ) ;
    buf_clk cell_9227 ( .C (clk), .D (signal_14114), .Q (signal_14115) ) ;
    buf_clk cell_9235 ( .C (clk), .D (signal_14122), .Q (signal_14123) ) ;
    buf_clk cell_9243 ( .C (clk), .D (signal_14130), .Q (signal_14131) ) ;
    buf_clk cell_9251 ( .C (clk), .D (signal_14138), .Q (signal_14139) ) ;
    buf_clk cell_9259 ( .C (clk), .D (signal_14146), .Q (signal_14147) ) ;
    buf_clk cell_9267 ( .C (clk), .D (signal_14154), .Q (signal_14155) ) ;
    buf_clk cell_9275 ( .C (clk), .D (signal_14162), .Q (signal_14163) ) ;
    buf_clk cell_9283 ( .C (clk), .D (signal_14170), .Q (signal_14171) ) ;
    buf_clk cell_9291 ( .C (clk), .D (signal_14178), .Q (signal_14179) ) ;
    buf_clk cell_9299 ( .C (clk), .D (signal_14186), .Q (signal_14187) ) ;
    buf_clk cell_9307 ( .C (clk), .D (signal_14194), .Q (signal_14195) ) ;
    buf_clk cell_9315 ( .C (clk), .D (signal_14202), .Q (signal_14203) ) ;
    buf_clk cell_9323 ( .C (clk), .D (signal_14210), .Q (signal_14211) ) ;
    buf_clk cell_9331 ( .C (clk), .D (signal_14218), .Q (signal_14219) ) ;
    buf_clk cell_9339 ( .C (clk), .D (signal_14226), .Q (signal_14227) ) ;
    buf_clk cell_9347 ( .C (clk), .D (signal_14234), .Q (signal_14235) ) ;
    buf_clk cell_9355 ( .C (clk), .D (signal_14242), .Q (signal_14243) ) ;
    buf_clk cell_9363 ( .C (clk), .D (signal_14250), .Q (signal_14251) ) ;
    buf_clk cell_9371 ( .C (clk), .D (signal_14258), .Q (signal_14259) ) ;
    buf_clk cell_9379 ( .C (clk), .D (signal_14266), .Q (signal_14267) ) ;
    buf_clk cell_9387 ( .C (clk), .D (signal_14274), .Q (signal_14275) ) ;
    buf_clk cell_9395 ( .C (clk), .D (signal_14282), .Q (signal_14283) ) ;
    buf_clk cell_9403 ( .C (clk), .D (signal_14290), .Q (signal_14291) ) ;
    buf_clk cell_9411 ( .C (clk), .D (signal_14298), .Q (signal_14299) ) ;
    buf_clk cell_9419 ( .C (clk), .D (signal_14306), .Q (signal_14307) ) ;
    buf_clk cell_9427 ( .C (clk), .D (signal_14314), .Q (signal_14315) ) ;
    buf_clk cell_9435 ( .C (clk), .D (signal_14322), .Q (signal_14323) ) ;
    buf_clk cell_9443 ( .C (clk), .D (signal_14330), .Q (signal_14331) ) ;
    buf_clk cell_9451 ( .C (clk), .D (signal_14338), .Q (signal_14339) ) ;
    buf_clk cell_9459 ( .C (clk), .D (signal_14346), .Q (signal_14347) ) ;
    buf_clk cell_9467 ( .C (clk), .D (signal_14354), .Q (signal_14355) ) ;
    buf_clk cell_9475 ( .C (clk), .D (signal_14362), .Q (signal_14363) ) ;
    buf_clk cell_9483 ( .C (clk), .D (signal_14370), .Q (signal_14371) ) ;
    buf_clk cell_9491 ( .C (clk), .D (signal_14378), .Q (signal_14379) ) ;
    buf_clk cell_9499 ( .C (clk), .D (signal_14386), .Q (signal_14387) ) ;
    buf_clk cell_9507 ( .C (clk), .D (signal_14394), .Q (signal_14395) ) ;
    buf_clk cell_9515 ( .C (clk), .D (signal_14402), .Q (signal_14403) ) ;
    buf_clk cell_9523 ( .C (clk), .D (signal_14410), .Q (signal_14411) ) ;
    buf_clk cell_9531 ( .C (clk), .D (signal_14418), .Q (signal_14419) ) ;
    buf_clk cell_9539 ( .C (clk), .D (signal_14426), .Q (signal_14427) ) ;
    buf_clk cell_9547 ( .C (clk), .D (signal_14434), .Q (signal_14435) ) ;
    buf_clk cell_9555 ( .C (clk), .D (signal_14442), .Q (signal_14443) ) ;
    buf_clk cell_9563 ( .C (clk), .D (signal_14450), .Q (signal_14451) ) ;
    buf_clk cell_9571 ( .C (clk), .D (signal_14458), .Q (signal_14459) ) ;
    buf_clk cell_9579 ( .C (clk), .D (signal_14466), .Q (signal_14467) ) ;
    buf_clk cell_9587 ( .C (clk), .D (signal_14474), .Q (signal_14475) ) ;
    buf_clk cell_9595 ( .C (clk), .D (signal_14482), .Q (signal_14483) ) ;
    buf_clk cell_9603 ( .C (clk), .D (signal_14490), .Q (signal_14491) ) ;
    buf_clk cell_9611 ( .C (clk), .D (signal_14498), .Q (signal_14499) ) ;
    buf_clk cell_9619 ( .C (clk), .D (signal_14506), .Q (signal_14507) ) ;
    buf_clk cell_9627 ( .C (clk), .D (signal_14514), .Q (signal_14515) ) ;
    buf_clk cell_9635 ( .C (clk), .D (signal_14522), .Q (signal_14523) ) ;
    buf_clk cell_9643 ( .C (clk), .D (signal_14530), .Q (signal_14531) ) ;
    buf_clk cell_9651 ( .C (clk), .D (signal_14538), .Q (signal_14539) ) ;
    buf_clk cell_9659 ( .C (clk), .D (signal_14546), .Q (signal_14547) ) ;
    buf_clk cell_9667 ( .C (clk), .D (signal_14554), .Q (signal_14555) ) ;
    buf_clk cell_9675 ( .C (clk), .D (signal_14562), .Q (signal_14563) ) ;
    buf_clk cell_9683 ( .C (clk), .D (signal_14570), .Q (signal_14571) ) ;
    buf_clk cell_9691 ( .C (clk), .D (signal_14578), .Q (signal_14579) ) ;
    buf_clk cell_9699 ( .C (clk), .D (signal_14586), .Q (signal_14587) ) ;
    buf_clk cell_9707 ( .C (clk), .D (signal_14594), .Q (signal_14595) ) ;
    buf_clk cell_9715 ( .C (clk), .D (signal_14602), .Q (signal_14603) ) ;
    buf_clk cell_9723 ( .C (clk), .D (signal_14610), .Q (signal_14611) ) ;
    buf_clk cell_9731 ( .C (clk), .D (signal_14618), .Q (signal_14619) ) ;
    buf_clk cell_9739 ( .C (clk), .D (signal_14626), .Q (signal_14627) ) ;
    buf_clk cell_9747 ( .C (clk), .D (signal_14634), .Q (signal_14635) ) ;
    buf_clk cell_9755 ( .C (clk), .D (signal_14642), .Q (signal_14643) ) ;
    buf_clk cell_9763 ( .C (clk), .D (signal_14650), .Q (signal_14651) ) ;
    buf_clk cell_9771 ( .C (clk), .D (signal_14658), .Q (signal_14659) ) ;
    buf_clk cell_9779 ( .C (clk), .D (signal_14666), .Q (signal_14667) ) ;
    buf_clk cell_9787 ( .C (clk), .D (signal_14674), .Q (signal_14675) ) ;
    buf_clk cell_9795 ( .C (clk), .D (signal_14682), .Q (signal_14683) ) ;
    buf_clk cell_9803 ( .C (clk), .D (signal_14690), .Q (signal_14691) ) ;
    buf_clk cell_9811 ( .C (clk), .D (signal_14698), .Q (signal_14699) ) ;
    buf_clk cell_9819 ( .C (clk), .D (signal_14706), .Q (signal_14707) ) ;
    buf_clk cell_9827 ( .C (clk), .D (signal_14714), .Q (signal_14715) ) ;
    buf_clk cell_9835 ( .C (clk), .D (signal_14722), .Q (signal_14723) ) ;
    buf_clk cell_9843 ( .C (clk), .D (signal_14730), .Q (signal_14731) ) ;
    buf_clk cell_9851 ( .C (clk), .D (signal_14738), .Q (signal_14739) ) ;
    buf_clk cell_9859 ( .C (clk), .D (signal_14746), .Q (signal_14747) ) ;
    buf_clk cell_9867 ( .C (clk), .D (signal_14754), .Q (signal_14755) ) ;
    buf_clk cell_9875 ( .C (clk), .D (signal_14762), .Q (signal_14763) ) ;
    buf_clk cell_9883 ( .C (clk), .D (signal_14770), .Q (signal_14771) ) ;
    buf_clk cell_9891 ( .C (clk), .D (signal_14778), .Q (signal_14779) ) ;
    buf_clk cell_9899 ( .C (clk), .D (signal_14786), .Q (signal_14787) ) ;
    buf_clk cell_9907 ( .C (clk), .D (signal_14794), .Q (signal_14795) ) ;
    buf_clk cell_9915 ( .C (clk), .D (signal_14802), .Q (signal_14803) ) ;
    buf_clk cell_9923 ( .C (clk), .D (signal_14810), .Q (signal_14811) ) ;
    buf_clk cell_9931 ( .C (clk), .D (signal_14818), .Q (signal_14819) ) ;
    buf_clk cell_9939 ( .C (clk), .D (signal_14826), .Q (signal_14827) ) ;
    buf_clk cell_9947 ( .C (clk), .D (signal_14834), .Q (signal_14835) ) ;
    buf_clk cell_9955 ( .C (clk), .D (signal_14842), .Q (signal_14843) ) ;
    buf_clk cell_9963 ( .C (clk), .D (signal_14850), .Q (signal_14851) ) ;
    buf_clk cell_9971 ( .C (clk), .D (signal_14858), .Q (signal_14859) ) ;
    buf_clk cell_9979 ( .C (clk), .D (signal_14866), .Q (signal_14867) ) ;
    buf_clk cell_9987 ( .C (clk), .D (signal_14874), .Q (signal_14875) ) ;
    buf_clk cell_9995 ( .C (clk), .D (signal_14882), .Q (signal_14883) ) ;
    buf_clk cell_10003 ( .C (clk), .D (signal_14890), .Q (signal_14891) ) ;
    buf_clk cell_10011 ( .C (clk), .D (signal_14898), .Q (signal_14899) ) ;
    buf_clk cell_10019 ( .C (clk), .D (signal_14906), .Q (signal_14907) ) ;
    buf_clk cell_10027 ( .C (clk), .D (signal_14914), .Q (signal_14915) ) ;
    buf_clk cell_10035 ( .C (clk), .D (signal_14922), .Q (signal_14923) ) ;
    buf_clk cell_10043 ( .C (clk), .D (signal_14930), .Q (signal_14931) ) ;
    buf_clk cell_10051 ( .C (clk), .D (signal_14938), .Q (signal_14939) ) ;
    buf_clk cell_10059 ( .C (clk), .D (signal_14946), .Q (signal_14947) ) ;
    buf_clk cell_10067 ( .C (clk), .D (signal_14954), .Q (signal_14955) ) ;
    buf_clk cell_10075 ( .C (clk), .D (signal_14962), .Q (signal_14963) ) ;
    buf_clk cell_10083 ( .C (clk), .D (signal_14970), .Q (signal_14971) ) ;
    buf_clk cell_10091 ( .C (clk), .D (signal_14978), .Q (signal_14979) ) ;
    buf_clk cell_10099 ( .C (clk), .D (signal_14986), .Q (signal_14987) ) ;
    buf_clk cell_10107 ( .C (clk), .D (signal_14994), .Q (signal_14995) ) ;
    buf_clk cell_10115 ( .C (clk), .D (signal_15002), .Q (signal_15003) ) ;
    buf_clk cell_10123 ( .C (clk), .D (signal_15010), .Q (signal_15011) ) ;
    buf_clk cell_10131 ( .C (clk), .D (signal_15018), .Q (signal_15019) ) ;
    buf_clk cell_10139 ( .C (clk), .D (signal_15026), .Q (signal_15027) ) ;
    buf_clk cell_10147 ( .C (clk), .D (signal_15034), .Q (signal_15035) ) ;
    buf_clk cell_10155 ( .C (clk), .D (signal_15042), .Q (signal_15043) ) ;
    buf_clk cell_10163 ( .C (clk), .D (signal_15050), .Q (signal_15051) ) ;
    buf_clk cell_10171 ( .C (clk), .D (signal_15058), .Q (signal_15059) ) ;
    buf_clk cell_10179 ( .C (clk), .D (signal_15066), .Q (signal_15067) ) ;
    buf_clk cell_10187 ( .C (clk), .D (signal_15074), .Q (signal_15075) ) ;
    buf_clk cell_10195 ( .C (clk), .D (signal_15082), .Q (signal_15083) ) ;
    buf_clk cell_10203 ( .C (clk), .D (signal_15090), .Q (signal_15091) ) ;
    buf_clk cell_10211 ( .C (clk), .D (signal_15098), .Q (signal_15099) ) ;
    buf_clk cell_10219 ( .C (clk), .D (signal_15106), .Q (signal_15107) ) ;
    buf_clk cell_10227 ( .C (clk), .D (signal_15114), .Q (signal_15115) ) ;
    buf_clk cell_10235 ( .C (clk), .D (signal_15122), .Q (signal_15123) ) ;
    buf_clk cell_10243 ( .C (clk), .D (signal_15130), .Q (signal_15131) ) ;
    buf_clk cell_10251 ( .C (clk), .D (signal_15138), .Q (signal_15139) ) ;
    buf_clk cell_10259 ( .C (clk), .D (signal_15146), .Q (signal_15147) ) ;
    buf_clk cell_10267 ( .C (clk), .D (signal_15154), .Q (signal_15155) ) ;
    buf_clk cell_10275 ( .C (clk), .D (signal_15162), .Q (signal_15163) ) ;
    buf_clk cell_10283 ( .C (clk), .D (signal_15170), .Q (signal_15171) ) ;
    buf_clk cell_10291 ( .C (clk), .D (signal_15178), .Q (signal_15179) ) ;
    buf_clk cell_10299 ( .C (clk), .D (signal_15186), .Q (signal_15187) ) ;
    buf_clk cell_10307 ( .C (clk), .D (signal_15194), .Q (signal_15195) ) ;
    buf_clk cell_10315 ( .C (clk), .D (signal_15202), .Q (signal_15203) ) ;
    buf_clk cell_10323 ( .C (clk), .D (signal_15210), .Q (signal_15211) ) ;
    buf_clk cell_10331 ( .C (clk), .D (signal_15218), .Q (signal_15219) ) ;
    buf_clk cell_10339 ( .C (clk), .D (signal_15226), .Q (signal_15227) ) ;
    buf_clk cell_10347 ( .C (clk), .D (signal_15234), .Q (signal_15235) ) ;
    buf_clk cell_10355 ( .C (clk), .D (signal_15242), .Q (signal_15243) ) ;
    buf_clk cell_10363 ( .C (clk), .D (signal_15250), .Q (signal_15251) ) ;
    buf_clk cell_10371 ( .C (clk), .D (signal_15258), .Q (signal_15259) ) ;
    buf_clk cell_10379 ( .C (clk), .D (signal_15266), .Q (signal_15267) ) ;
    buf_clk cell_10387 ( .C (clk), .D (signal_15274), .Q (signal_15275) ) ;
    buf_clk cell_10395 ( .C (clk), .D (signal_15282), .Q (signal_15283) ) ;
    buf_clk cell_10403 ( .C (clk), .D (signal_15290), .Q (signal_15291) ) ;
    buf_clk cell_10411 ( .C (clk), .D (signal_15298), .Q (signal_15299) ) ;
    buf_clk cell_10419 ( .C (clk), .D (signal_15306), .Q (signal_15307) ) ;
    buf_clk cell_10427 ( .C (clk), .D (signal_15314), .Q (signal_15315) ) ;
    buf_clk cell_10435 ( .C (clk), .D (signal_15322), .Q (signal_15323) ) ;
    buf_clk cell_10443 ( .C (clk), .D (signal_15330), .Q (signal_15331) ) ;
    buf_clk cell_10451 ( .C (clk), .D (signal_15338), .Q (signal_15339) ) ;
    buf_clk cell_10459 ( .C (clk), .D (signal_15346), .Q (signal_15347) ) ;
    buf_clk cell_10467 ( .C (clk), .D (signal_15354), .Q (signal_15355) ) ;
    buf_clk cell_10475 ( .C (clk), .D (signal_15362), .Q (signal_15363) ) ;
    buf_clk cell_10483 ( .C (clk), .D (signal_15370), .Q (signal_15371) ) ;
    buf_clk cell_10491 ( .C (clk), .D (signal_15378), .Q (signal_15379) ) ;
    buf_clk cell_10499 ( .C (clk), .D (signal_15386), .Q (signal_15387) ) ;
    buf_clk cell_10507 ( .C (clk), .D (signal_15394), .Q (signal_15395) ) ;
    buf_clk cell_10515 ( .C (clk), .D (signal_15402), .Q (signal_15403) ) ;
    buf_clk cell_10523 ( .C (clk), .D (signal_15410), .Q (signal_15411) ) ;
    buf_clk cell_10531 ( .C (clk), .D (signal_15418), .Q (signal_15419) ) ;
    buf_clk cell_10539 ( .C (clk), .D (signal_15426), .Q (signal_15427) ) ;
    buf_clk cell_10547 ( .C (clk), .D (signal_15434), .Q (signal_15435) ) ;
    buf_clk cell_10555 ( .C (clk), .D (signal_15442), .Q (signal_15443) ) ;
    buf_clk cell_10563 ( .C (clk), .D (signal_15450), .Q (signal_15451) ) ;
    buf_clk cell_10571 ( .C (clk), .D (signal_15458), .Q (signal_15459) ) ;
    buf_clk cell_10579 ( .C (clk), .D (signal_15466), .Q (signal_15467) ) ;
    buf_clk cell_10587 ( .C (clk), .D (signal_15474), .Q (signal_15475) ) ;
    buf_clk cell_10595 ( .C (clk), .D (signal_15482), .Q (signal_15483) ) ;
    buf_clk cell_10603 ( .C (clk), .D (signal_15490), .Q (signal_15491) ) ;
    buf_clk cell_10611 ( .C (clk), .D (signal_15498), .Q (signal_15499) ) ;
    buf_clk cell_10619 ( .C (clk), .D (signal_15506), .Q (signal_15507) ) ;
    buf_clk cell_10627 ( .C (clk), .D (signal_15514), .Q (signal_15515) ) ;
    buf_clk cell_10635 ( .C (clk), .D (signal_15522), .Q (signal_15523) ) ;
    buf_clk cell_10643 ( .C (clk), .D (signal_15530), .Q (signal_15531) ) ;
    buf_clk cell_10651 ( .C (clk), .D (signal_15538), .Q (signal_15539) ) ;
    buf_clk cell_10659 ( .C (clk), .D (signal_15546), .Q (signal_15547) ) ;
    buf_clk cell_10667 ( .C (clk), .D (signal_15554), .Q (signal_15555) ) ;
    buf_clk cell_10675 ( .C (clk), .D (signal_15562), .Q (signal_15563) ) ;
    buf_clk cell_10683 ( .C (clk), .D (signal_15570), .Q (signal_15571) ) ;
    buf_clk cell_10691 ( .C (clk), .D (signal_15578), .Q (signal_15579) ) ;
    buf_clk cell_10699 ( .C (clk), .D (signal_15586), .Q (signal_15587) ) ;
    buf_clk cell_10707 ( .C (clk), .D (signal_15594), .Q (signal_15595) ) ;
    buf_clk cell_10715 ( .C (clk), .D (signal_15602), .Q (signal_15603) ) ;
    buf_clk cell_10723 ( .C (clk), .D (signal_15610), .Q (signal_15611) ) ;
    buf_clk cell_10731 ( .C (clk), .D (signal_15618), .Q (signal_15619) ) ;
    buf_clk cell_10739 ( .C (clk), .D (signal_15626), .Q (signal_15627) ) ;
    buf_clk cell_10747 ( .C (clk), .D (signal_15634), .Q (signal_15635) ) ;
    buf_clk cell_10755 ( .C (clk), .D (signal_15642), .Q (signal_15643) ) ;
    buf_clk cell_10763 ( .C (clk), .D (signal_15650), .Q (signal_15651) ) ;
    buf_clk cell_10771 ( .C (clk), .D (signal_15658), .Q (signal_15659) ) ;
    buf_clk cell_10779 ( .C (clk), .D (signal_15666), .Q (signal_15667) ) ;
    buf_clk cell_10787 ( .C (clk), .D (signal_15674), .Q (signal_15675) ) ;
    buf_clk cell_10795 ( .C (clk), .D (signal_15682), .Q (signal_15683) ) ;
    buf_clk cell_10803 ( .C (clk), .D (signal_15690), .Q (signal_15691) ) ;
    buf_clk cell_10811 ( .C (clk), .D (signal_15698), .Q (signal_15699) ) ;
    buf_clk cell_10819 ( .C (clk), .D (signal_15706), .Q (signal_15707) ) ;
    buf_clk cell_10827 ( .C (clk), .D (signal_15714), .Q (signal_15715) ) ;
    buf_clk cell_10835 ( .C (clk), .D (signal_15722), .Q (signal_15723) ) ;
    buf_clk cell_10843 ( .C (clk), .D (signal_15730), .Q (signal_15731) ) ;
    buf_clk cell_10851 ( .C (clk), .D (signal_15738), .Q (signal_15739) ) ;
    buf_clk cell_10859 ( .C (clk), .D (signal_15746), .Q (signal_15747) ) ;
    buf_clk cell_10867 ( .C (clk), .D (signal_15754), .Q (signal_15755) ) ;
    buf_clk cell_10875 ( .C (clk), .D (signal_15762), .Q (signal_15763) ) ;
    buf_clk cell_10883 ( .C (clk), .D (signal_15770), .Q (signal_15771) ) ;
    buf_clk cell_10891 ( .C (clk), .D (signal_15778), .Q (signal_15779) ) ;
    buf_clk cell_10899 ( .C (clk), .D (signal_15786), .Q (signal_15787) ) ;
    buf_clk cell_10907 ( .C (clk), .D (signal_15794), .Q (signal_15795) ) ;
    buf_clk cell_10915 ( .C (clk), .D (signal_15802), .Q (signal_15803) ) ;
    buf_clk cell_10923 ( .C (clk), .D (signal_15810), .Q (signal_15811) ) ;
    buf_clk cell_10931 ( .C (clk), .D (signal_15818), .Q (signal_15819) ) ;
    buf_clk cell_10939 ( .C (clk), .D (signal_15826), .Q (signal_15827) ) ;
    buf_clk cell_10947 ( .C (clk), .D (signal_15834), .Q (signal_15835) ) ;
    buf_clk cell_10955 ( .C (clk), .D (signal_15842), .Q (signal_15843) ) ;
    buf_clk cell_10963 ( .C (clk), .D (signal_15850), .Q (signal_15851) ) ;
    buf_clk cell_10971 ( .C (clk), .D (signal_15858), .Q (signal_15859) ) ;
    buf_clk cell_10979 ( .C (clk), .D (signal_15866), .Q (signal_15867) ) ;
    buf_clk cell_10987 ( .C (clk), .D (signal_15874), .Q (signal_15875) ) ;
    buf_clk cell_10995 ( .C (clk), .D (signal_15882), .Q (signal_15883) ) ;
    buf_clk cell_11003 ( .C (clk), .D (signal_15890), .Q (signal_15891) ) ;
    buf_clk cell_11011 ( .C (clk), .D (signal_15898), .Q (signal_15899) ) ;
    buf_clk cell_11019 ( .C (clk), .D (signal_15906), .Q (signal_15907) ) ;
    buf_clk cell_11027 ( .C (clk), .D (signal_15914), .Q (signal_15915) ) ;
    buf_clk cell_11035 ( .C (clk), .D (signal_15922), .Q (signal_15923) ) ;
    buf_clk cell_11043 ( .C (clk), .D (signal_15930), .Q (signal_15931) ) ;
    buf_clk cell_11051 ( .C (clk), .D (signal_15938), .Q (signal_15939) ) ;
    buf_clk cell_11059 ( .C (clk), .D (signal_15946), .Q (signal_15947) ) ;
    buf_clk cell_11067 ( .C (clk), .D (signal_15954), .Q (signal_15955) ) ;
    buf_clk cell_11075 ( .C (clk), .D (signal_15962), .Q (signal_15963) ) ;
    buf_clk cell_11083 ( .C (clk), .D (signal_15970), .Q (signal_15971) ) ;
    buf_clk cell_11091 ( .C (clk), .D (signal_15978), .Q (signal_15979) ) ;
    buf_clk cell_11099 ( .C (clk), .D (signal_15986), .Q (signal_15987) ) ;
    buf_clk cell_11107 ( .C (clk), .D (signal_15994), .Q (signal_15995) ) ;
    buf_clk cell_11115 ( .C (clk), .D (signal_16002), .Q (signal_16003) ) ;
    buf_clk cell_11123 ( .C (clk), .D (signal_16010), .Q (signal_16011) ) ;
    buf_clk cell_11131 ( .C (clk), .D (signal_16018), .Q (signal_16019) ) ;
    buf_clk cell_11139 ( .C (clk), .D (signal_16026), .Q (signal_16027) ) ;
    buf_clk cell_11147 ( .C (clk), .D (signal_16034), .Q (signal_16035) ) ;
    buf_clk cell_11155 ( .C (clk), .D (signal_16042), .Q (signal_16043) ) ;
    buf_clk cell_11163 ( .C (clk), .D (signal_16050), .Q (signal_16051) ) ;
    buf_clk cell_11171 ( .C (clk), .D (signal_16058), .Q (signal_16059) ) ;
    buf_clk cell_11179 ( .C (clk), .D (signal_16066), .Q (signal_16067) ) ;
    buf_clk cell_11187 ( .C (clk), .D (signal_16074), .Q (signal_16075) ) ;
    buf_clk cell_11195 ( .C (clk), .D (signal_16082), .Q (signal_16083) ) ;
    buf_clk cell_11203 ( .C (clk), .D (signal_16090), .Q (signal_16091) ) ;
    buf_clk cell_11211 ( .C (clk), .D (signal_16098), .Q (signal_16099) ) ;
    buf_clk cell_11219 ( .C (clk), .D (signal_16106), .Q (signal_16107) ) ;
    buf_clk cell_11227 ( .C (clk), .D (signal_16114), .Q (signal_16115) ) ;
    buf_clk cell_11235 ( .C (clk), .D (signal_16122), .Q (signal_16123) ) ;
    buf_clk cell_11243 ( .C (clk), .D (signal_16130), .Q (signal_16131) ) ;
    buf_clk cell_11251 ( .C (clk), .D (signal_16138), .Q (signal_16139) ) ;
    buf_clk cell_11259 ( .C (clk), .D (signal_16146), .Q (signal_16147) ) ;
    buf_clk cell_11267 ( .C (clk), .D (signal_16154), .Q (signal_16155) ) ;
    buf_clk cell_11275 ( .C (clk), .D (signal_16162), .Q (signal_16163) ) ;
    buf_clk cell_11283 ( .C (clk), .D (signal_16170), .Q (signal_16171) ) ;
    buf_clk cell_11291 ( .C (clk), .D (signal_16178), .Q (signal_16179) ) ;
    buf_clk cell_11299 ( .C (clk), .D (signal_16186), .Q (signal_16187) ) ;
    buf_clk cell_11307 ( .C (clk), .D (signal_16194), .Q (signal_16195) ) ;
    buf_clk cell_11315 ( .C (clk), .D (signal_16202), .Q (signal_16203) ) ;
    buf_clk cell_11323 ( .C (clk), .D (signal_16210), .Q (signal_16211) ) ;
    buf_clk cell_11331 ( .C (clk), .D (signal_16218), .Q (signal_16219) ) ;
    buf_clk cell_11339 ( .C (clk), .D (signal_16226), .Q (signal_16227) ) ;
    buf_clk cell_11347 ( .C (clk), .D (signal_16234), .Q (signal_16235) ) ;
    buf_clk cell_11355 ( .C (clk), .D (signal_16242), .Q (signal_16243) ) ;
    buf_clk cell_11363 ( .C (clk), .D (signal_16250), .Q (signal_16251) ) ;
    buf_clk cell_11371 ( .C (clk), .D (signal_16258), .Q (signal_16259) ) ;
    buf_clk cell_11379 ( .C (clk), .D (signal_16266), .Q (signal_16267) ) ;
    buf_clk cell_11387 ( .C (clk), .D (signal_16274), .Q (signal_16275) ) ;
    buf_clk cell_11395 ( .C (clk), .D (signal_16282), .Q (signal_16283) ) ;
    buf_clk cell_11403 ( .C (clk), .D (signal_16290), .Q (signal_16291) ) ;
    buf_clk cell_11411 ( .C (clk), .D (signal_16298), .Q (signal_16299) ) ;
    buf_clk cell_11419 ( .C (clk), .D (signal_16306), .Q (signal_16307) ) ;
    buf_clk cell_11427 ( .C (clk), .D (signal_16314), .Q (signal_16315) ) ;
    buf_clk cell_11435 ( .C (clk), .D (signal_16322), .Q (signal_16323) ) ;
    buf_clk cell_11443 ( .C (clk), .D (signal_16330), .Q (signal_16331) ) ;
    buf_clk cell_11451 ( .C (clk), .D (signal_16338), .Q (signal_16339) ) ;
    buf_clk cell_11459 ( .C (clk), .D (signal_16346), .Q (signal_16347) ) ;
    buf_clk cell_11467 ( .C (clk), .D (signal_16354), .Q (signal_16355) ) ;
    buf_clk cell_11475 ( .C (clk), .D (signal_16362), .Q (signal_16363) ) ;
    buf_clk cell_11483 ( .C (clk), .D (signal_16370), .Q (signal_16371) ) ;
    buf_clk cell_11491 ( .C (clk), .D (signal_16378), .Q (signal_16379) ) ;
    buf_clk cell_11499 ( .C (clk), .D (signal_16386), .Q (signal_16387) ) ;
    buf_clk cell_11507 ( .C (clk), .D (signal_16394), .Q (signal_16395) ) ;
    buf_clk cell_11515 ( .C (clk), .D (signal_16402), .Q (signal_16403) ) ;
    buf_clk cell_11523 ( .C (clk), .D (signal_16410), .Q (signal_16411) ) ;
    buf_clk cell_11531 ( .C (clk), .D (signal_16418), .Q (signal_16419) ) ;
    buf_clk cell_11539 ( .C (clk), .D (signal_16426), .Q (signal_16427) ) ;
    buf_clk cell_11547 ( .C (clk), .D (signal_16434), .Q (signal_16435) ) ;
    buf_clk cell_11555 ( .C (clk), .D (signal_16442), .Q (signal_16443) ) ;
    buf_clk cell_11563 ( .C (clk), .D (signal_16450), .Q (signal_16451) ) ;
    buf_clk cell_11571 ( .C (clk), .D (signal_16458), .Q (signal_16459) ) ;
    buf_clk cell_11579 ( .C (clk), .D (signal_16466), .Q (signal_16467) ) ;
    buf_clk cell_11587 ( .C (clk), .D (signal_16474), .Q (signal_16475) ) ;
    buf_clk cell_11595 ( .C (clk), .D (signal_16482), .Q (signal_16483) ) ;
    buf_clk cell_11603 ( .C (clk), .D (signal_16490), .Q (signal_16491) ) ;
    buf_clk cell_11611 ( .C (clk), .D (signal_16498), .Q (signal_16499) ) ;
    buf_clk cell_11619 ( .C (clk), .D (signal_16506), .Q (signal_16507) ) ;
    buf_clk cell_11627 ( .C (clk), .D (signal_16514), .Q (signal_16515) ) ;
    buf_clk cell_11635 ( .C (clk), .D (signal_16522), .Q (signal_16523) ) ;
    buf_clk cell_11643 ( .C (clk), .D (signal_16530), .Q (signal_16531) ) ;
    buf_clk cell_11651 ( .C (clk), .D (signal_16538), .Q (signal_16539) ) ;
    buf_clk cell_11659 ( .C (clk), .D (signal_16546), .Q (signal_16547) ) ;
    buf_clk cell_11667 ( .C (clk), .D (signal_16554), .Q (signal_16555) ) ;
    buf_clk cell_11675 ( .C (clk), .D (signal_16562), .Q (signal_16563) ) ;
    buf_clk cell_11683 ( .C (clk), .D (signal_16570), .Q (signal_16571) ) ;
    buf_clk cell_11691 ( .C (clk), .D (signal_16578), .Q (signal_16579) ) ;
    buf_clk cell_11699 ( .C (clk), .D (signal_16586), .Q (signal_16587) ) ;
    buf_clk cell_11707 ( .C (clk), .D (signal_16594), .Q (signal_16595) ) ;
    buf_clk cell_11715 ( .C (clk), .D (signal_16602), .Q (signal_16603) ) ;
    buf_clk cell_11723 ( .C (clk), .D (signal_16610), .Q (signal_16611) ) ;
    buf_clk cell_11731 ( .C (clk), .D (signal_16618), .Q (signal_16619) ) ;
    buf_clk cell_11739 ( .C (clk), .D (signal_16626), .Q (signal_16627) ) ;
    buf_clk cell_11747 ( .C (clk), .D (signal_16634), .Q (signal_16635) ) ;
    buf_clk cell_11755 ( .C (clk), .D (signal_16642), .Q (signal_16643) ) ;
    buf_clk cell_11763 ( .C (clk), .D (signal_16650), .Q (signal_16651) ) ;
    buf_clk cell_11771 ( .C (clk), .D (signal_16658), .Q (signal_16659) ) ;
    buf_clk cell_11779 ( .C (clk), .D (signal_16666), .Q (signal_16667) ) ;
    buf_clk cell_11787 ( .C (clk), .D (signal_16674), .Q (signal_16675) ) ;
    buf_clk cell_11795 ( .C (clk), .D (signal_16682), .Q (signal_16683) ) ;
    buf_clk cell_11803 ( .C (clk), .D (signal_16690), .Q (signal_16691) ) ;
    buf_clk cell_11811 ( .C (clk), .D (signal_16698), .Q (signal_16699) ) ;
    buf_clk cell_11819 ( .C (clk), .D (signal_16706), .Q (signal_16707) ) ;
    buf_clk cell_11827 ( .C (clk), .D (signal_16714), .Q (signal_16715) ) ;
    buf_clk cell_11835 ( .C (clk), .D (signal_16722), .Q (signal_16723) ) ;
    buf_clk cell_11843 ( .C (clk), .D (signal_16730), .Q (signal_16731) ) ;
    buf_clk cell_11851 ( .C (clk), .D (signal_16738), .Q (signal_16739) ) ;
    buf_clk cell_11859 ( .C (clk), .D (signal_16746), .Q (signal_16747) ) ;
    buf_clk cell_11867 ( .C (clk), .D (signal_16754), .Q (signal_16755) ) ;
    buf_clk cell_11875 ( .C (clk), .D (signal_16762), .Q (signal_16763) ) ;
    buf_clk cell_11883 ( .C (clk), .D (signal_16770), .Q (signal_16771) ) ;
    buf_clk cell_11891 ( .C (clk), .D (signal_16778), .Q (signal_16779) ) ;
    buf_clk cell_11899 ( .C (clk), .D (signal_16786), .Q (signal_16787) ) ;
    buf_clk cell_11907 ( .C (clk), .D (signal_16794), .Q (signal_16795) ) ;
    buf_clk cell_11915 ( .C (clk), .D (signal_16802), .Q (signal_16803) ) ;
    buf_clk cell_11923 ( .C (clk), .D (signal_16810), .Q (signal_16811) ) ;
    buf_clk cell_11931 ( .C (clk), .D (signal_16818), .Q (signal_16819) ) ;
    buf_clk cell_11939 ( .C (clk), .D (signal_16826), .Q (signal_16827) ) ;
    buf_clk cell_11947 ( .C (clk), .D (signal_16834), .Q (signal_16835) ) ;
    buf_clk cell_11955 ( .C (clk), .D (signal_16842), .Q (signal_16843) ) ;
    buf_clk cell_11963 ( .C (clk), .D (signal_16850), .Q (signal_16851) ) ;
    buf_clk cell_11971 ( .C (clk), .D (signal_16858), .Q (signal_16859) ) ;
    buf_clk cell_11979 ( .C (clk), .D (signal_16866), .Q (signal_16867) ) ;
    buf_clk cell_11987 ( .C (clk), .D (signal_16874), .Q (signal_16875) ) ;
    buf_clk cell_11995 ( .C (clk), .D (signal_16882), .Q (signal_16883) ) ;
    buf_clk cell_12003 ( .C (clk), .D (signal_16890), .Q (signal_16891) ) ;
    buf_clk cell_12011 ( .C (clk), .D (signal_16898), .Q (signal_16899) ) ;
    buf_clk cell_12019 ( .C (clk), .D (signal_16906), .Q (signal_16907) ) ;
    buf_clk cell_12027 ( .C (clk), .D (signal_16914), .Q (signal_16915) ) ;
    buf_clk cell_12035 ( .C (clk), .D (signal_16922), .Q (signal_16923) ) ;
    buf_clk cell_12043 ( .C (clk), .D (signal_16930), .Q (signal_16931) ) ;
    buf_clk cell_12051 ( .C (clk), .D (signal_16938), .Q (signal_16939) ) ;
    buf_clk cell_12059 ( .C (clk), .D (signal_16946), .Q (signal_16947) ) ;
    buf_clk cell_12067 ( .C (clk), .D (signal_16954), .Q (signal_16955) ) ;
    buf_clk cell_12075 ( .C (clk), .D (signal_16962), .Q (signal_16963) ) ;
    buf_clk cell_12083 ( .C (clk), .D (signal_16970), .Q (signal_16971) ) ;
    buf_clk cell_12091 ( .C (clk), .D (signal_16978), .Q (signal_16979) ) ;
    buf_clk cell_12099 ( .C (clk), .D (signal_16986), .Q (signal_16987) ) ;
    buf_clk cell_12107 ( .C (clk), .D (signal_16994), .Q (signal_16995) ) ;
    buf_clk cell_12115 ( .C (clk), .D (signal_17002), .Q (signal_17003) ) ;
    buf_clk cell_12123 ( .C (clk), .D (signal_17010), .Q (signal_17011) ) ;
    buf_clk cell_12131 ( .C (clk), .D (signal_17018), .Q (signal_17019) ) ;
    buf_clk cell_12139 ( .C (clk), .D (signal_17026), .Q (signal_17027) ) ;
    buf_clk cell_12147 ( .C (clk), .D (signal_17034), .Q (signal_17035) ) ;
    buf_clk cell_12155 ( .C (clk), .D (signal_17042), .Q (signal_17043) ) ;
    buf_clk cell_12163 ( .C (clk), .D (signal_17050), .Q (signal_17051) ) ;
    buf_clk cell_12171 ( .C (clk), .D (signal_17058), .Q (signal_17059) ) ;
    buf_clk cell_12179 ( .C (clk), .D (signal_17066), .Q (signal_17067) ) ;
    buf_clk cell_12187 ( .C (clk), .D (signal_17074), .Q (signal_17075) ) ;
    buf_clk cell_12195 ( .C (clk), .D (signal_17082), .Q (signal_17083) ) ;
    buf_clk cell_12203 ( .C (clk), .D (signal_17090), .Q (signal_17091) ) ;
    buf_clk cell_12211 ( .C (clk), .D (signal_17098), .Q (signal_17099) ) ;
    buf_clk cell_12219 ( .C (clk), .D (signal_17106), .Q (signal_17107) ) ;
    buf_clk cell_12227 ( .C (clk), .D (signal_17114), .Q (signal_17115) ) ;
    buf_clk cell_12235 ( .C (clk), .D (signal_17122), .Q (signal_17123) ) ;
    buf_clk cell_12243 ( .C (clk), .D (signal_17130), .Q (signal_17131) ) ;
    buf_clk cell_12251 ( .C (clk), .D (signal_17138), .Q (signal_17139) ) ;
    buf_clk cell_12259 ( .C (clk), .D (signal_17146), .Q (signal_17147) ) ;
    buf_clk cell_12267 ( .C (clk), .D (signal_17154), .Q (signal_17155) ) ;
    buf_clk cell_12275 ( .C (clk), .D (signal_17162), .Q (signal_17163) ) ;
    buf_clk cell_12283 ( .C (clk), .D (signal_17170), .Q (signal_17171) ) ;
    buf_clk cell_12291 ( .C (clk), .D (signal_17178), .Q (signal_17179) ) ;
    buf_clk cell_12299 ( .C (clk), .D (signal_17186), .Q (signal_17187) ) ;
    buf_clk cell_12307 ( .C (clk), .D (signal_17194), .Q (signal_17195) ) ;
    buf_clk cell_12315 ( .C (clk), .D (signal_17202), .Q (signal_17203) ) ;
    buf_clk cell_12323 ( .C (clk), .D (signal_17210), .Q (signal_17211) ) ;
    buf_clk cell_12331 ( .C (clk), .D (signal_17218), .Q (signal_17219) ) ;
    buf_clk cell_12339 ( .C (clk), .D (signal_17226), .Q (signal_17227) ) ;
    buf_clk cell_12347 ( .C (clk), .D (signal_17234), .Q (signal_17235) ) ;
    buf_clk cell_12355 ( .C (clk), .D (signal_17242), .Q (signal_17243) ) ;
    buf_clk cell_12363 ( .C (clk), .D (signal_17250), .Q (signal_17251) ) ;
    buf_clk cell_12371 ( .C (clk), .D (signal_17258), .Q (signal_17259) ) ;
    buf_clk cell_12379 ( .C (clk), .D (signal_17266), .Q (signal_17267) ) ;
    buf_clk cell_12387 ( .C (clk), .D (signal_17274), .Q (signal_17275) ) ;
    buf_clk cell_12395 ( .C (clk), .D (signal_17282), .Q (signal_17283) ) ;
    buf_clk cell_12403 ( .C (clk), .D (signal_17290), .Q (signal_17291) ) ;
    buf_clk cell_12411 ( .C (clk), .D (signal_17298), .Q (signal_17299) ) ;
    buf_clk cell_12419 ( .C (clk), .D (signal_17306), .Q (signal_17307) ) ;
    buf_clk cell_12427 ( .C (clk), .D (signal_17314), .Q (signal_17315) ) ;
    buf_clk cell_12435 ( .C (clk), .D (signal_17322), .Q (signal_17323) ) ;
    buf_clk cell_12443 ( .C (clk), .D (signal_17330), .Q (signal_17331) ) ;
    buf_clk cell_12451 ( .C (clk), .D (signal_17338), .Q (signal_17339) ) ;
    buf_clk cell_12459 ( .C (clk), .D (signal_17346), .Q (signal_17347) ) ;
    buf_clk cell_12467 ( .C (clk), .D (signal_17354), .Q (signal_17355) ) ;
    buf_clk cell_12475 ( .C (clk), .D (signal_17362), .Q (signal_17363) ) ;
    buf_clk cell_12483 ( .C (clk), .D (signal_17370), .Q (signal_17371) ) ;
    buf_clk cell_12491 ( .C (clk), .D (signal_17378), .Q (signal_17379) ) ;
    buf_clk cell_12499 ( .C (clk), .D (signal_17386), .Q (signal_17387) ) ;
    buf_clk cell_12507 ( .C (clk), .D (signal_17394), .Q (signal_17395) ) ;
    buf_clk cell_12515 ( .C (clk), .D (signal_17402), .Q (signal_17403) ) ;
    buf_clk cell_12523 ( .C (clk), .D (signal_17410), .Q (signal_17411) ) ;
    buf_clk cell_12531 ( .C (clk), .D (signal_17418), .Q (signal_17419) ) ;
    buf_clk cell_12539 ( .C (clk), .D (signal_17426), .Q (signal_17427) ) ;
    buf_clk cell_12547 ( .C (clk), .D (signal_17434), .Q (signal_17435) ) ;
    buf_clk cell_12555 ( .C (clk), .D (signal_17442), .Q (signal_17443) ) ;
    buf_clk cell_12563 ( .C (clk), .D (signal_17450), .Q (signal_17451) ) ;
    buf_clk cell_12571 ( .C (clk), .D (signal_17458), .Q (signal_17459) ) ;
    buf_clk cell_12579 ( .C (clk), .D (signal_17466), .Q (signal_17467) ) ;
    buf_clk cell_12587 ( .C (clk), .D (signal_17474), .Q (signal_17475) ) ;
    buf_clk cell_12595 ( .C (clk), .D (signal_17482), .Q (signal_17483) ) ;
    buf_clk cell_12603 ( .C (clk), .D (signal_17490), .Q (signal_17491) ) ;
    buf_clk cell_12611 ( .C (clk), .D (signal_17498), .Q (signal_17499) ) ;
    buf_clk cell_12619 ( .C (clk), .D (signal_17506), .Q (signal_17507) ) ;
    buf_clk cell_12627 ( .C (clk), .D (signal_17514), .Q (signal_17515) ) ;
    buf_clk cell_12635 ( .C (clk), .D (signal_17522), .Q (signal_17523) ) ;
    buf_clk cell_12643 ( .C (clk), .D (signal_17530), .Q (signal_17531) ) ;
    buf_clk cell_12651 ( .C (clk), .D (signal_17538), .Q (signal_17539) ) ;
    buf_clk cell_12659 ( .C (clk), .D (signal_17546), .Q (signal_17547) ) ;
    buf_clk cell_12667 ( .C (clk), .D (signal_17554), .Q (signal_17555) ) ;
    buf_clk cell_12675 ( .C (clk), .D (signal_17562), .Q (signal_17563) ) ;
    buf_clk cell_12683 ( .C (clk), .D (signal_17570), .Q (signal_17571) ) ;
    buf_clk cell_12691 ( .C (clk), .D (signal_17578), .Q (signal_17579) ) ;
    buf_clk cell_12699 ( .C (clk), .D (signal_17586), .Q (signal_17587) ) ;
    buf_clk cell_12707 ( .C (clk), .D (signal_17594), .Q (signal_17595) ) ;
    buf_clk cell_12715 ( .C (clk), .D (signal_17602), .Q (signal_17603) ) ;
    buf_clk cell_12723 ( .C (clk), .D (signal_17610), .Q (signal_17611) ) ;
    buf_clk cell_12731 ( .C (clk), .D (signal_17618), .Q (signal_17619) ) ;
    buf_clk cell_12739 ( .C (clk), .D (signal_17626), .Q (signal_17627) ) ;
    buf_clk cell_12747 ( .C (clk), .D (signal_17634), .Q (signal_17635) ) ;
    buf_clk cell_12755 ( .C (clk), .D (signal_17642), .Q (signal_17643) ) ;
    buf_clk cell_12763 ( .C (clk), .D (signal_17650), .Q (signal_17651) ) ;
    buf_clk cell_12771 ( .C (clk), .D (signal_17658), .Q (signal_17659) ) ;
    buf_clk cell_12779 ( .C (clk), .D (signal_17666), .Q (signal_17667) ) ;
    buf_clk cell_12787 ( .C (clk), .D (signal_17674), .Q (signal_17675) ) ;
    buf_clk cell_12795 ( .C (clk), .D (signal_17682), .Q (signal_17683) ) ;
    buf_clk cell_12803 ( .C (clk), .D (signal_17690), .Q (signal_17691) ) ;
    buf_clk cell_12811 ( .C (clk), .D (signal_17698), .Q (signal_17699) ) ;
    buf_clk cell_12819 ( .C (clk), .D (signal_17706), .Q (signal_17707) ) ;
    buf_clk cell_12827 ( .C (clk), .D (signal_17714), .Q (signal_17715) ) ;
    buf_clk cell_12835 ( .C (clk), .D (signal_17722), .Q (signal_17723) ) ;
    buf_clk cell_12843 ( .C (clk), .D (signal_17730), .Q (signal_17731) ) ;
    buf_clk cell_12851 ( .C (clk), .D (signal_17738), .Q (signal_17739) ) ;
    buf_clk cell_12859 ( .C (clk), .D (signal_17746), .Q (signal_17747) ) ;
    buf_clk cell_12867 ( .C (clk), .D (signal_17754), .Q (signal_17755) ) ;
    buf_clk cell_12875 ( .C (clk), .D (signal_17762), .Q (signal_17763) ) ;
    buf_clk cell_12883 ( .C (clk), .D (signal_17770), .Q (signal_17771) ) ;
    buf_clk cell_12891 ( .C (clk), .D (signal_17778), .Q (signal_17779) ) ;
    buf_clk cell_12899 ( .C (clk), .D (signal_17786), .Q (signal_17787) ) ;
    buf_clk cell_12907 ( .C (clk), .D (signal_17794), .Q (signal_17795) ) ;
    buf_clk cell_12915 ( .C (clk), .D (signal_17802), .Q (signal_17803) ) ;
    buf_clk cell_12923 ( .C (clk), .D (signal_17810), .Q (signal_17811) ) ;
    buf_clk cell_12931 ( .C (clk), .D (signal_17818), .Q (signal_17819) ) ;
    buf_clk cell_12939 ( .C (clk), .D (signal_17826), .Q (signal_17827) ) ;
    buf_clk cell_12947 ( .C (clk), .D (signal_17834), .Q (signal_17835) ) ;
    buf_clk cell_12955 ( .C (clk), .D (signal_17842), .Q (signal_17843) ) ;
    buf_clk cell_12963 ( .C (clk), .D (signal_17850), .Q (signal_17851) ) ;
    buf_clk cell_12971 ( .C (clk), .D (signal_17858), .Q (signal_17859) ) ;
    buf_clk cell_12979 ( .C (clk), .D (signal_17866), .Q (signal_17867) ) ;
    buf_clk cell_12987 ( .C (clk), .D (signal_17874), .Q (signal_17875) ) ;
    buf_clk cell_12995 ( .C (clk), .D (signal_17882), .Q (signal_17883) ) ;
    buf_clk cell_13003 ( .C (clk), .D (signal_17890), .Q (signal_17891) ) ;
    buf_clk cell_13011 ( .C (clk), .D (signal_17898), .Q (signal_17899) ) ;
    buf_clk cell_13019 ( .C (clk), .D (signal_17906), .Q (signal_17907) ) ;
    buf_clk cell_13027 ( .C (clk), .D (signal_17914), .Q (signal_17915) ) ;
    buf_clk cell_13035 ( .C (clk), .D (signal_17922), .Q (signal_17923) ) ;
    buf_clk cell_13043 ( .C (clk), .D (signal_17930), .Q (signal_17931) ) ;
    buf_clk cell_13051 ( .C (clk), .D (signal_17938), .Q (signal_17939) ) ;
    buf_clk cell_13059 ( .C (clk), .D (signal_17946), .Q (signal_17947) ) ;
    buf_clk cell_13067 ( .C (clk), .D (signal_17954), .Q (signal_17955) ) ;
    buf_clk cell_13075 ( .C (clk), .D (signal_17962), .Q (signal_17963) ) ;
    buf_clk cell_13083 ( .C (clk), .D (signal_17970), .Q (signal_17971) ) ;
    buf_clk cell_13091 ( .C (clk), .D (signal_17978), .Q (signal_17979) ) ;
    buf_clk cell_13099 ( .C (clk), .D (signal_17986), .Q (signal_17987) ) ;
    buf_clk cell_13107 ( .C (clk), .D (signal_17994), .Q (signal_17995) ) ;
    buf_clk cell_13115 ( .C (clk), .D (signal_18002), .Q (signal_18003) ) ;
    buf_clk cell_13123 ( .C (clk), .D (signal_18010), .Q (signal_18011) ) ;
    buf_clk cell_13131 ( .C (clk), .D (signal_18018), .Q (signal_18019) ) ;
    buf_clk cell_13139 ( .C (clk), .D (signal_18026), .Q (signal_18027) ) ;
    buf_clk cell_13147 ( .C (clk), .D (signal_18034), .Q (signal_18035) ) ;
    buf_clk cell_13155 ( .C (clk), .D (signal_18042), .Q (signal_18043) ) ;
    buf_clk cell_13163 ( .C (clk), .D (signal_18050), .Q (signal_18051) ) ;
    buf_clk cell_13171 ( .C (clk), .D (signal_18058), .Q (signal_18059) ) ;
    buf_clk cell_13179 ( .C (clk), .D (signal_18066), .Q (signal_18067) ) ;
    buf_clk cell_13187 ( .C (clk), .D (signal_18074), .Q (signal_18075) ) ;
    buf_clk cell_13195 ( .C (clk), .D (signal_18082), .Q (signal_18083) ) ;
    buf_clk cell_13203 ( .C (clk), .D (signal_18090), .Q (signal_18091) ) ;
    buf_clk cell_13211 ( .C (clk), .D (signal_18098), .Q (signal_18099) ) ;
    buf_clk cell_13219 ( .C (clk), .D (signal_18106), .Q (signal_18107) ) ;
    buf_clk cell_13227 ( .C (clk), .D (signal_18114), .Q (signal_18115) ) ;
    buf_clk cell_13235 ( .C (clk), .D (signal_18122), .Q (signal_18123) ) ;
    buf_clk cell_13243 ( .C (clk), .D (signal_18130), .Q (signal_18131) ) ;
    buf_clk cell_13251 ( .C (clk), .D (signal_18138), .Q (signal_18139) ) ;
    buf_clk cell_13259 ( .C (clk), .D (signal_18146), .Q (signal_18147) ) ;
    buf_clk cell_13267 ( .C (clk), .D (signal_18154), .Q (signal_18155) ) ;
    buf_clk cell_13275 ( .C (clk), .D (signal_18162), .Q (signal_18163) ) ;
    buf_clk cell_17591 ( .C (clk), .D (signal_22478), .Q (signal_22479) ) ;
    buf_clk cell_17599 ( .C (clk), .D (signal_22486), .Q (signal_22487) ) ;
    buf_clk cell_17607 ( .C (clk), .D (signal_22494), .Q (signal_22495) ) ;
    buf_clk cell_17615 ( .C (clk), .D (signal_22502), .Q (signal_22503) ) ;
    buf_clk cell_17623 ( .C (clk), .D (signal_22510), .Q (signal_22511) ) ;
    buf_clk cell_17631 ( .C (clk), .D (signal_22518), .Q (signal_22519) ) ;
    buf_clk cell_17639 ( .C (clk), .D (signal_22526), .Q (signal_22527) ) ;
    buf_clk cell_17647 ( .C (clk), .D (signal_22534), .Q (signal_22535) ) ;
    buf_clk cell_17655 ( .C (clk), .D (signal_22542), .Q (signal_22543) ) ;
    buf_clk cell_17663 ( .C (clk), .D (signal_22550), .Q (signal_22551) ) ;
    buf_clk cell_17671 ( .C (clk), .D (signal_22558), .Q (signal_22559) ) ;
    buf_clk cell_17679 ( .C (clk), .D (signal_22566), .Q (signal_22567) ) ;
    buf_clk cell_17687 ( .C (clk), .D (signal_22574), .Q (signal_22575) ) ;
    buf_clk cell_17695 ( .C (clk), .D (signal_22582), .Q (signal_22583) ) ;
    buf_clk cell_17703 ( .C (clk), .D (signal_22590), .Q (signal_22591) ) ;
    buf_clk cell_17711 ( .C (clk), .D (signal_22598), .Q (signal_22599) ) ;
    buf_clk cell_17719 ( .C (clk), .D (signal_22606), .Q (signal_22607) ) ;
    buf_clk cell_17727 ( .C (clk), .D (signal_22614), .Q (signal_22615) ) ;
    buf_clk cell_17735 ( .C (clk), .D (signal_22622), .Q (signal_22623) ) ;
    buf_clk cell_17743 ( .C (clk), .D (signal_22630), .Q (signal_22631) ) ;
    buf_clk cell_17751 ( .C (clk), .D (signal_22638), .Q (signal_22639) ) ;
    buf_clk cell_17759 ( .C (clk), .D (signal_22646), .Q (signal_22647) ) ;
    buf_clk cell_17767 ( .C (clk), .D (signal_22654), .Q (signal_22655) ) ;
    buf_clk cell_17775 ( .C (clk), .D (signal_22662), .Q (signal_22663) ) ;
    buf_clk cell_17783 ( .C (clk), .D (signal_22670), .Q (signal_22671) ) ;
    buf_clk cell_17791 ( .C (clk), .D (signal_22678), .Q (signal_22679) ) ;
    buf_clk cell_17799 ( .C (clk), .D (signal_22686), .Q (signal_22687) ) ;
    buf_clk cell_17807 ( .C (clk), .D (signal_22694), .Q (signal_22695) ) ;
    buf_clk cell_17815 ( .C (clk), .D (signal_22702), .Q (signal_22703) ) ;
    buf_clk cell_17823 ( .C (clk), .D (signal_22710), .Q (signal_22711) ) ;
    buf_clk cell_17831 ( .C (clk), .D (signal_22718), .Q (signal_22719) ) ;
    buf_clk cell_17839 ( .C (clk), .D (signal_22726), .Q (signal_22727) ) ;
    buf_clk cell_17847 ( .C (clk), .D (signal_22734), .Q (signal_22735) ) ;
    buf_clk cell_17855 ( .C (clk), .D (signal_22742), .Q (signal_22743) ) ;
    buf_clk cell_17863 ( .C (clk), .D (signal_22750), .Q (signal_22751) ) ;
    buf_clk cell_17871 ( .C (clk), .D (signal_22758), .Q (signal_22759) ) ;
    buf_clk cell_17879 ( .C (clk), .D (signal_22766), .Q (signal_22767) ) ;
    buf_clk cell_17887 ( .C (clk), .D (signal_22774), .Q (signal_22775) ) ;
    buf_clk cell_17895 ( .C (clk), .D (signal_22782), .Q (signal_22783) ) ;
    buf_clk cell_17903 ( .C (clk), .D (signal_22790), .Q (signal_22791) ) ;
    buf_clk cell_17911 ( .C (clk), .D (signal_22798), .Q (signal_22799) ) ;
    buf_clk cell_17919 ( .C (clk), .D (signal_22806), .Q (signal_22807) ) ;
    buf_clk cell_17927 ( .C (clk), .D (signal_22814), .Q (signal_22815) ) ;
    buf_clk cell_17935 ( .C (clk), .D (signal_22822), .Q (signal_22823) ) ;
    buf_clk cell_17943 ( .C (clk), .D (signal_22830), .Q (signal_22831) ) ;
    buf_clk cell_17951 ( .C (clk), .D (signal_22838), .Q (signal_22839) ) ;
    buf_clk cell_17959 ( .C (clk), .D (signal_22846), .Q (signal_22847) ) ;
    buf_clk cell_17967 ( .C (clk), .D (signal_22854), .Q (signal_22855) ) ;
    buf_clk cell_17975 ( .C (clk), .D (signal_22862), .Q (signal_22863) ) ;
    buf_clk cell_17983 ( .C (clk), .D (signal_22870), .Q (signal_22871) ) ;
    buf_clk cell_17991 ( .C (clk), .D (signal_22878), .Q (signal_22879) ) ;
    buf_clk cell_17999 ( .C (clk), .D (signal_22886), .Q (signal_22887) ) ;
    buf_clk cell_18007 ( .C (clk), .D (signal_22894), .Q (signal_22895) ) ;
    buf_clk cell_18015 ( .C (clk), .D (signal_22902), .Q (signal_22903) ) ;
    buf_clk cell_18023 ( .C (clk), .D (signal_22910), .Q (signal_22911) ) ;
    buf_clk cell_18031 ( .C (clk), .D (signal_22918), .Q (signal_22919) ) ;
    buf_clk cell_18039 ( .C (clk), .D (signal_22926), .Q (signal_22927) ) ;
    buf_clk cell_18047 ( .C (clk), .D (signal_22934), .Q (signal_22935) ) ;
    buf_clk cell_18055 ( .C (clk), .D (signal_22942), .Q (signal_22943) ) ;
    buf_clk cell_18063 ( .C (clk), .D (signal_22950), .Q (signal_22951) ) ;
    buf_clk cell_18071 ( .C (clk), .D (signal_22958), .Q (signal_22959) ) ;
    buf_clk cell_18079 ( .C (clk), .D (signal_22966), .Q (signal_22967) ) ;
    buf_clk cell_18087 ( .C (clk), .D (signal_22974), .Q (signal_22975) ) ;
    buf_clk cell_18095 ( .C (clk), .D (signal_22982), .Q (signal_22983) ) ;
    buf_clk cell_18103 ( .C (clk), .D (signal_22990), .Q (signal_22991) ) ;
    buf_clk cell_18111 ( .C (clk), .D (signal_22998), .Q (signal_22999) ) ;
    buf_clk cell_18119 ( .C (clk), .D (signal_23006), .Q (signal_23007) ) ;
    buf_clk cell_18127 ( .C (clk), .D (signal_23014), .Q (signal_23015) ) ;
    buf_clk cell_18135 ( .C (clk), .D (signal_23022), .Q (signal_23023) ) ;
    buf_clk cell_18143 ( .C (clk), .D (signal_23030), .Q (signal_23031) ) ;
    buf_clk cell_18151 ( .C (clk), .D (signal_23038), .Q (signal_23039) ) ;
    buf_clk cell_18159 ( .C (clk), .D (signal_23046), .Q (signal_23047) ) ;
    buf_clk cell_18167 ( .C (clk), .D (signal_23054), .Q (signal_23055) ) ;
    buf_clk cell_18175 ( .C (clk), .D (signal_23062), .Q (signal_23063) ) ;
    buf_clk cell_18183 ( .C (clk), .D (signal_23070), .Q (signal_23071) ) ;
    buf_clk cell_18191 ( .C (clk), .D (signal_23078), .Q (signal_23079) ) ;
    buf_clk cell_18199 ( .C (clk), .D (signal_23086), .Q (signal_23087) ) ;
    buf_clk cell_18207 ( .C (clk), .D (signal_23094), .Q (signal_23095) ) ;
    buf_clk cell_18215 ( .C (clk), .D (signal_23102), .Q (signal_23103) ) ;
    buf_clk cell_18223 ( .C (clk), .D (signal_23110), .Q (signal_23111) ) ;
    buf_clk cell_18231 ( .C (clk), .D (signal_23118), .Q (signal_23119) ) ;
    buf_clk cell_18239 ( .C (clk), .D (signal_23126), .Q (signal_23127) ) ;
    buf_clk cell_18247 ( .C (clk), .D (signal_23134), .Q (signal_23135) ) ;
    buf_clk cell_18255 ( .C (clk), .D (signal_23142), .Q (signal_23143) ) ;
    buf_clk cell_18263 ( .C (clk), .D (signal_23150), .Q (signal_23151) ) ;
    buf_clk cell_18271 ( .C (clk), .D (signal_23158), .Q (signal_23159) ) ;
    buf_clk cell_18279 ( .C (clk), .D (signal_23166), .Q (signal_23167) ) ;
    buf_clk cell_18287 ( .C (clk), .D (signal_23174), .Q (signal_23175) ) ;
    buf_clk cell_18295 ( .C (clk), .D (signal_23182), .Q (signal_23183) ) ;
    buf_clk cell_18303 ( .C (clk), .D (signal_23190), .Q (signal_23191) ) ;
    buf_clk cell_18311 ( .C (clk), .D (signal_23198), .Q (signal_23199) ) ;
    buf_clk cell_18319 ( .C (clk), .D (signal_23206), .Q (signal_23207) ) ;
    buf_clk cell_18327 ( .C (clk), .D (signal_23214), .Q (signal_23215) ) ;
    buf_clk cell_18335 ( .C (clk), .D (signal_23222), .Q (signal_23223) ) ;
    buf_clk cell_18343 ( .C (clk), .D (signal_23230), .Q (signal_23231) ) ;
    buf_clk cell_18351 ( .C (clk), .D (signal_23238), .Q (signal_23239) ) ;
    buf_clk cell_18359 ( .C (clk), .D (signal_23246), .Q (signal_23247) ) ;
    buf_clk cell_18367 ( .C (clk), .D (signal_23254), .Q (signal_23255) ) ;
    buf_clk cell_18375 ( .C (clk), .D (signal_23262), .Q (signal_23263) ) ;
    buf_clk cell_18383 ( .C (clk), .D (signal_23270), .Q (signal_23271) ) ;
    buf_clk cell_18391 ( .C (clk), .D (signal_23278), .Q (signal_23279) ) ;
    buf_clk cell_18399 ( .C (clk), .D (signal_23286), .Q (signal_23287) ) ;
    buf_clk cell_18401 ( .C (clk), .D (signal_18566), .Q (signal_23289) ) ;
    buf_clk cell_18403 ( .C (clk), .D (signal_18572), .Q (signal_23291) ) ;
    buf_clk cell_18411 ( .C (clk), .D (signal_23298), .Q (signal_23299) ) ;
    buf_clk cell_18419 ( .C (clk), .D (signal_23306), .Q (signal_23307) ) ;
    buf_clk cell_18427 ( .C (clk), .D (signal_23314), .Q (signal_23315) ) ;
    buf_clk cell_18435 ( .C (clk), .D (signal_23322), .Q (signal_23323) ) ;
    buf_clk cell_18443 ( .C (clk), .D (signal_23330), .Q (signal_23331) ) ;
    buf_clk cell_18451 ( .C (clk), .D (signal_23338), .Q (signal_23339) ) ;
    buf_clk cell_18459 ( .C (clk), .D (signal_23346), .Q (signal_23347) ) ;
    buf_clk cell_18467 ( .C (clk), .D (signal_23354), .Q (signal_23355) ) ;
    buf_clk cell_18475 ( .C (clk), .D (signal_23362), .Q (signal_23363) ) ;
    buf_clk cell_18483 ( .C (clk), .D (signal_23370), .Q (signal_23371) ) ;
    buf_clk cell_18491 ( .C (clk), .D (signal_23378), .Q (signal_23379) ) ;
    buf_clk cell_18499 ( .C (clk), .D (signal_23386), .Q (signal_23387) ) ;
    buf_clk cell_18507 ( .C (clk), .D (signal_23394), .Q (signal_23395) ) ;
    buf_clk cell_18515 ( .C (clk), .D (signal_23402), .Q (signal_23403) ) ;
    buf_clk cell_18523 ( .C (clk), .D (signal_23410), .Q (signal_23411) ) ;
    buf_clk cell_18531 ( .C (clk), .D (signal_23418), .Q (signal_23419) ) ;
    buf_clk cell_18539 ( .C (clk), .D (signal_23426), .Q (signal_23427) ) ;
    buf_clk cell_18547 ( .C (clk), .D (signal_23434), .Q (signal_23435) ) ;
    buf_clk cell_18555 ( .C (clk), .D (signal_23442), .Q (signal_23443) ) ;
    buf_clk cell_18563 ( .C (clk), .D (signal_23450), .Q (signal_23451) ) ;
    buf_clk cell_18571 ( .C (clk), .D (signal_23458), .Q (signal_23459) ) ;
    buf_clk cell_18579 ( .C (clk), .D (signal_23466), .Q (signal_23467) ) ;
    buf_clk cell_18587 ( .C (clk), .D (signal_23474), .Q (signal_23475) ) ;
    buf_clk cell_18595 ( .C (clk), .D (signal_23482), .Q (signal_23483) ) ;
    buf_clk cell_18603 ( .C (clk), .D (signal_23490), .Q (signal_23491) ) ;
    buf_clk cell_18611 ( .C (clk), .D (signal_23498), .Q (signal_23499) ) ;
    buf_clk cell_18619 ( .C (clk), .D (signal_23506), .Q (signal_23507) ) ;
    buf_clk cell_18627 ( .C (clk), .D (signal_23514), .Q (signal_23515) ) ;
    buf_clk cell_18635 ( .C (clk), .D (signal_23522), .Q (signal_23523) ) ;
    buf_clk cell_18643 ( .C (clk), .D (signal_23530), .Q (signal_23531) ) ;
    buf_clk cell_18645 ( .C (clk), .D (signal_18470), .Q (signal_23533) ) ;
    buf_clk cell_18647 ( .C (clk), .D (signal_18476), .Q (signal_23535) ) ;
    buf_clk cell_18655 ( .C (clk), .D (signal_23542), .Q (signal_23543) ) ;
    buf_clk cell_18663 ( .C (clk), .D (signal_23550), .Q (signal_23551) ) ;
    buf_clk cell_18671 ( .C (clk), .D (signal_23558), .Q (signal_23559) ) ;
    buf_clk cell_18679 ( .C (clk), .D (signal_23566), .Q (signal_23567) ) ;
    buf_clk cell_18687 ( .C (clk), .D (signal_23574), .Q (signal_23575) ) ;
    buf_clk cell_18695 ( .C (clk), .D (signal_23582), .Q (signal_23583) ) ;
    buf_clk cell_18703 ( .C (clk), .D (signal_23590), .Q (signal_23591) ) ;
    buf_clk cell_18711 ( .C (clk), .D (signal_23598), .Q (signal_23599) ) ;
    buf_clk cell_18719 ( .C (clk), .D (signal_23606), .Q (signal_23607) ) ;
    buf_clk cell_18727 ( .C (clk), .D (signal_23614), .Q (signal_23615) ) ;
    buf_clk cell_18735 ( .C (clk), .D (signal_23622), .Q (signal_23623) ) ;
    buf_clk cell_18743 ( .C (clk), .D (signal_23630), .Q (signal_23631) ) ;
    buf_clk cell_18745 ( .C (clk), .D (signal_18662), .Q (signal_23633) ) ;
    buf_clk cell_18747 ( .C (clk), .D (signal_18668), .Q (signal_23635) ) ;
    buf_clk cell_18755 ( .C (clk), .D (signal_23642), .Q (signal_23643) ) ;
    buf_clk cell_18763 ( .C (clk), .D (signal_23650), .Q (signal_23651) ) ;
    buf_clk cell_18771 ( .C (clk), .D (signal_23658), .Q (signal_23659) ) ;
    buf_clk cell_18779 ( .C (clk), .D (signal_23666), .Q (signal_23667) ) ;
    buf_clk cell_18787 ( .C (clk), .D (signal_23674), .Q (signal_23675) ) ;
    buf_clk cell_18795 ( .C (clk), .D (signal_23682), .Q (signal_23683) ) ;
    buf_clk cell_18803 ( .C (clk), .D (signal_23690), .Q (signal_23691) ) ;
    buf_clk cell_18811 ( .C (clk), .D (signal_23698), .Q (signal_23699) ) ;
    buf_clk cell_18819 ( .C (clk), .D (signal_23706), .Q (signal_23707) ) ;
    buf_clk cell_18827 ( .C (clk), .D (signal_23714), .Q (signal_23715) ) ;
    buf_clk cell_18835 ( .C (clk), .D (signal_23722), .Q (signal_23723) ) ;
    buf_clk cell_18843 ( .C (clk), .D (signal_23730), .Q (signal_23731) ) ;
    buf_clk cell_18851 ( .C (clk), .D (signal_23738), .Q (signal_23739) ) ;
    buf_clk cell_18859 ( .C (clk), .D (signal_23746), .Q (signal_23747) ) ;
    buf_clk cell_18867 ( .C (clk), .D (signal_23754), .Q (signal_23755) ) ;
    buf_clk cell_18875 ( .C (clk), .D (signal_23762), .Q (signal_23763) ) ;
    buf_clk cell_18883 ( .C (clk), .D (signal_23770), .Q (signal_23771) ) ;
    buf_clk cell_18891 ( .C (clk), .D (signal_23778), .Q (signal_23779) ) ;
    buf_clk cell_18899 ( .C (clk), .D (signal_23786), .Q (signal_23787) ) ;
    buf_clk cell_18907 ( .C (clk), .D (signal_23794), .Q (signal_23795) ) ;
    buf_clk cell_18915 ( .C (clk), .D (signal_23802), .Q (signal_23803) ) ;
    buf_clk cell_18923 ( .C (clk), .D (signal_23810), .Q (signal_23811) ) ;
    buf_clk cell_18931 ( .C (clk), .D (signal_23818), .Q (signal_23819) ) ;
    buf_clk cell_18939 ( .C (clk), .D (signal_23826), .Q (signal_23827) ) ;
    buf_clk cell_18947 ( .C (clk), .D (signal_23834), .Q (signal_23835) ) ;
    buf_clk cell_18955 ( .C (clk), .D (signal_23842), .Q (signal_23843) ) ;
    buf_clk cell_18963 ( .C (clk), .D (signal_23850), .Q (signal_23851) ) ;
    buf_clk cell_18971 ( .C (clk), .D (signal_23858), .Q (signal_23859) ) ;
    buf_clk cell_18979 ( .C (clk), .D (signal_23866), .Q (signal_23867) ) ;
    buf_clk cell_18987 ( .C (clk), .D (signal_23874), .Q (signal_23875) ) ;
    buf_clk cell_18995 ( .C (clk), .D (signal_23882), .Q (signal_23883) ) ;
    buf_clk cell_19003 ( .C (clk), .D (signal_23890), .Q (signal_23891) ) ;
    buf_clk cell_19011 ( .C (clk), .D (signal_23898), .Q (signal_23899) ) ;
    buf_clk cell_19019 ( .C (clk), .D (signal_23906), .Q (signal_23907) ) ;
    buf_clk cell_19027 ( .C (clk), .D (signal_23914), .Q (signal_23915) ) ;
    buf_clk cell_19035 ( .C (clk), .D (signal_23922), .Q (signal_23923) ) ;
    buf_clk cell_19043 ( .C (clk), .D (signal_23930), .Q (signal_23931) ) ;
    buf_clk cell_19051 ( .C (clk), .D (signal_23938), .Q (signal_23939) ) ;
    buf_clk cell_19059 ( .C (clk), .D (signal_23946), .Q (signal_23947) ) ;
    buf_clk cell_19067 ( .C (clk), .D (signal_23954), .Q (signal_23955) ) ;
    buf_clk cell_19075 ( .C (clk), .D (signal_23962), .Q (signal_23963) ) ;
    buf_clk cell_19083 ( .C (clk), .D (signal_23970), .Q (signal_23971) ) ;
    buf_clk cell_19091 ( .C (clk), .D (signal_23978), .Q (signal_23979) ) ;
    buf_clk cell_19099 ( .C (clk), .D (signal_23986), .Q (signal_23987) ) ;
    buf_clk cell_19107 ( .C (clk), .D (signal_23994), .Q (signal_23995) ) ;
    buf_clk cell_19115 ( .C (clk), .D (signal_24002), .Q (signal_24003) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_28 ( .s (signal_13436), .b ({signal_10326, signal_3994}), .a ({signal_11320, signal_4122}), .c ({signal_11378, signal_3742}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_29 ( .s (signal_13436), .b ({signal_10344, signal_4415}), .a ({signal_11331, signal_4022}), .c ({signal_11379, signal_3642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_30 ( .s (signal_13436), .b ({signal_10516, signal_4414}), .a ({signal_11278, signal_4021}), .c ({signal_11380, signal_3641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_31 ( .s (signal_13436), .b ({signal_10515, signal_4413}), .a ({signal_11277, signal_4020}), .c ({signal_11381, signal_3640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_32 ( .s (signal_13436), .b ({signal_10341, signal_4420}), .a ({signal_11025, signal_4019}), .c ({signal_11169, signal_3639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_33 ( .s (signal_13436), .b ({signal_10327, signal_3890}), .a ({signal_11276, signal_4018}), .c ({signal_11382, signal_3638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_34 ( .s (signal_13436), .b ({signal_10532, signal_4410}), .a ({signal_11559, signal_4017}), .c ({signal_11575, signal_3637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_35 ( .s (signal_13436), .b ({signal_10381, signal_3888}), .a ({signal_11052, signal_4016}), .c ({signal_11170, signal_3636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_36 ( .s (signal_13444), .b ({signal_10380, signal_3887}), .a ({signal_11341, signal_4015}), .c ({signal_11383, signal_3635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_37 ( .s (signal_13452), .b ({signal_10379, signal_4407}), .a ({signal_11340, signal_4014}), .c ({signal_11384, signal_3634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_38 ( .s (signal_13460), .b ({signal_10531, signal_4406}), .a ({signal_11285, signal_4013}), .c ({signal_11385, signal_3633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_39 ( .s (signal_13468), .b ({signal_10402, signal_3984}), .a ({signal_11146, signal_4112}), .c ({signal_11171, signal_3732}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_40 ( .s (signal_13476), .b ({signal_10530, signal_4405}), .a ({signal_11284, signal_4012}), .c ({signal_11386, signal_3632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_41 ( .s (signal_13484), .b ({signal_10376, signal_4412}), .a ({signal_11047, signal_4011}), .c ({signal_11172, signal_3631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_42 ( .s (signal_13476), .b ({signal_10331, signal_3882}), .a ({signal_11283, signal_4010}), .c ({signal_11387, signal_3630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_43 ( .s (signal_13468), .b ({signal_10544, signal_4402}), .a ({signal_11562, signal_4009}), .c ({signal_11576, signal_3629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_44 ( .s (signal_13468), .b ({signal_10409, signal_3880}), .a ({signal_11044, signal_4008}), .c ({signal_11173, signal_3628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_45 ( .s (signal_13444), .b ({signal_10408, signal_3879}), .a ({signal_11338, signal_4007}), .c ({signal_11388, signal_3627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_46 ( .s (signal_13452), .b ({signal_10407, signal_4399}), .a ({signal_11336, signal_4006}), .c ({signal_11389, signal_3626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_47 ( .s (signal_13460), .b ({signal_10543, signal_4398}), .a ({signal_11282, signal_4005}), .c ({signal_11390, signal_3625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_48 ( .s (signal_13476), .b ({signal_10542, signal_4397}), .a ({signal_11281, signal_4004}), .c ({signal_11391, signal_3624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_49 ( .s (signal_13484), .b ({signal_10404, signal_4404}), .a ({signal_11038, signal_4003}), .c ({signal_11174, signal_3623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_50 ( .s (signal_13484), .b ({signal_10401, signal_3983}), .a ({signal_11377, signal_4111}), .c ({signal_11392, signal_3731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_51 ( .s (signal_13476), .b ({signal_10300, signal_3874}), .a ({signal_11273, signal_4002}), .c ({signal_11393, signal_3622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_52 ( .s (signal_13468), .b ({signal_10502, signal_4394}), .a ({signal_11560, signal_4001}), .c ({signal_11577, signal_3621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_53 ( .s (signal_13476), .b ({signal_10320, signal_3872}), .a ({signal_11036, signal_4000}), .c ({signal_11175, signal_3620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_54 ( .s (signal_13484), .b ({signal_10319, signal_3871}), .a ({signal_11334, signal_3999}), .c ({signal_11394, signal_3619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_55 ( .s (signal_13452), .b ({signal_10318, signal_4391}), .a ({signal_11333, signal_3998}), .c ({signal_11395, signal_3618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_13484), .b ({signal_10501, signal_4390}), .a ({signal_11280, signal_3997}), .c ({signal_11396, signal_3617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_13452), .b ({signal_10500, signal_4389}), .a ({signal_11279, signal_3996}), .c ({signal_11397, signal_3616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_13460), .b ({signal_10315, signal_4396}), .a ({signal_11030, signal_3995}), .c ({signal_11176, signal_3615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_13444), .b ({signal_10400, signal_4503}), .a ({signal_11376, signal_4110}), .c ({signal_11398, signal_3730}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_13460), .b ({signal_10540, signal_4502}), .a ({signal_11319, signal_4109}), .c ({signal_11399, signal_3729}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_13452), .b ({signal_10539, signal_4501}), .a ({signal_11318, signal_4108}), .c ({signal_11400, signal_3728}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_13460), .b ({signal_10397, signal_4508}), .a ({signal_11141, signal_4107}), .c ({signal_11177, signal_3727}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_13444), .b ({signal_10334, signal_3978}), .a ({signal_11317, signal_4106}), .c ({signal_11401, signal_3726}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_64 ( .s (signal_13468), .b ({signal_10553, signal_4498}), .a ({signal_11574, signal_4105}), .c ({signal_11578, signal_3725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_65 ( .s (signal_13476), .b ({signal_10430, signal_3976}), .a ({signal_11138, signal_4104}), .c ({signal_11178, signal_3724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_66 ( .s (signal_13484), .b ({signal_10429, signal_3975}), .a ({signal_11374, signal_4103}), .c ({signal_11402, signal_3723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_67 ( .s (signal_13468), .b ({signal_10529, signal_4514}), .a ({signal_11573, signal_4121}), .c ({signal_11579, signal_3741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_68 ( .s (signal_13476), .b ({signal_10428, signal_4495}), .a ({signal_11372, signal_4102}), .c ({signal_11403, signal_3722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_69 ( .s (signal_13452), .b ({signal_10552, signal_4494}), .a ({signal_11316, signal_4101}), .c ({signal_11404, signal_3721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_70 ( .s (signal_13460), .b ({signal_10551, signal_4493}), .a ({signal_11315, signal_4100}), .c ({signal_11405, signal_3720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_71 ( .s (signal_13444), .b ({signal_10425, signal_4500}), .a ({signal_11132, signal_4099}), .c ({signal_11179, signal_3719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_72 ( .s (signal_13484), .b ({signal_10325, signal_3970}), .a ({signal_11314, signal_4098}), .c ({signal_11406, signal_3718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_73 ( .s (signal_13468), .b ({signal_10526, signal_4490}), .a ({signal_11572, signal_4097}), .c ({signal_11580, signal_3717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_74 ( .s (signal_13452), .b ({signal_10367, signal_3968}), .a ({signal_11129, signal_4096}), .c ({signal_11180, signal_3716}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_75 ( .s (signal_13460), .b ({signal_10366, signal_3967}), .a ({signal_11370, signal_4095}), .c ({signal_11407, signal_3715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_76 ( .s (signal_13444), .b ({signal_10365, signal_4487}), .a ({signal_11369, signal_4094}), .c ({signal_11408, signal_3714}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_77 ( .s (signal_13476), .b ({signal_10525, signal_4486}), .a ({signal_11313, signal_4093}), .c ({signal_11409, signal_3713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_78 ( .s (signal_13444), .b ({signal_10374, signal_3992}), .a ({signal_11125, signal_4120}), .c ({signal_11181, signal_3740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_79 ( .s (signal_13484), .b ({signal_10524, signal_4485}), .a ({signal_11312, signal_4092}), .c ({signal_11410, signal_3712}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_80 ( .s (signal_13468), .b ({signal_10362, signal_4492}), .a ({signal_11123, signal_4091}), .c ({signal_11182, signal_3711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_81 ( .s (signal_13452), .b ({signal_10329, signal_3962}), .a ({signal_11308, signal_4090}), .c ({signal_11411, signal_3710}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_82 ( .s (signal_13460), .b ({signal_10538, signal_4482}), .a ({signal_11569, signal_4089}), .c ({signal_11581, signal_3709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_83 ( .s (signal_13444), .b ({signal_10395, signal_3960}), .a ({signal_11094, signal_4088}), .c ({signal_11183, signal_3708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_84 ( .s (signal_13484), .b ({signal_10394, signal_3959}), .a ({signal_11356, signal_4087}), .c ({signal_11412, signal_3707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_85 ( .s (signal_13484), .b ({signal_10393, signal_4479}), .a ({signal_11355, signal_4086}), .c ({signal_11413, signal_3706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_86 ( .s (signal_13484), .b ({signal_10537, signal_4478}), .a ({signal_11300, signal_4085}), .c ({signal_11414, signal_3705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_87 ( .s (signal_13484), .b ({signal_10536, signal_4477}), .a ({signal_11299, signal_4084}), .c ({signal_11415, signal_3704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_88 ( .s (signal_13484), .b ({signal_10390, signal_4484}), .a ({signal_11087, signal_4083}), .c ({signal_11184, signal_3703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_89 ( .s (signal_13484), .b ({signal_10373, signal_3991}), .a ({signal_11368, signal_4119}), .c ({signal_11416, signal_3739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_90 ( .s (signal_13484), .b ({signal_10333, signal_3954}), .a ({signal_11298, signal_4082}), .c ({signal_11417, signal_3702}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_13484), .b ({signal_10550, signal_4474}), .a ({signal_11567, signal_4081}), .c ({signal_11582, signal_3701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_92 ( .s (signal_13484), .b ({signal_10423, signal_3952}), .a ({signal_11114, signal_4080}), .c ({signal_11185, signal_3700}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_93 ( .s (signal_13484), .b ({signal_10422, signal_3951}), .a ({signal_11365, signal_4079}), .c ({signal_11418, signal_3699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_94 ( .s (signal_13484), .b ({signal_10421, signal_4471}), .a ({signal_11364, signal_4078}), .c ({signal_11419, signal_3698}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_95 ( .s (signal_13484), .b ({signal_10549, signal_4470}), .a ({signal_11307, signal_4077}), .c ({signal_11420, signal_3697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_96 ( .s (signal_13476), .b ({signal_10548, signal_4469}), .a ({signal_11306, signal_4076}), .c ({signal_11421, signal_3696}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_97 ( .s (signal_13476), .b ({signal_10418, signal_4476}), .a ({signal_11109, signal_4075}), .c ({signal_11186, signal_3695}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_98 ( .s (signal_13476), .b ({signal_10324, signal_3946}), .a ({signal_11305, signal_4074}), .c ({signal_11422, signal_3694}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_99 ( .s (signal_13476), .b ({signal_10523, signal_4466}), .a ({signal_11570, signal_4073}), .c ({signal_11583, signal_3693}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_100 ( .s (signal_13476), .b ({signal_10372, signal_4511}), .a ({signal_11367, signal_4118}), .c ({signal_11423, signal_3738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_101 ( .s (signal_13476), .b ({signal_10360, signal_3944}), .a ({signal_11106, signal_4072}), .c ({signal_11187, signal_3692}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_102 ( .s (signal_13476), .b ({signal_10359, signal_3943}), .a ({signal_11362, signal_4071}), .c ({signal_11424, signal_3691}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_103 ( .s (signal_13476), .b ({signal_10358, signal_4463}), .a ({signal_11360, signal_4070}), .c ({signal_11425, signal_3690}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_104 ( .s (signal_13476), .b ({signal_10522, signal_4462}), .a ({signal_11304, signal_4069}), .c ({signal_11426, signal_3689}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_105 ( .s (signal_13476), .b ({signal_10521, signal_4461}), .a ({signal_11303, signal_4068}), .c ({signal_11427, signal_3688}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_106 ( .s (signal_13476), .b ({signal_10355, signal_4468}), .a ({signal_11100, signal_4067}), .c ({signal_11188, signal_3687}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_107 ( .s (signal_13476), .b ({signal_10298, signal_3938}), .a ({signal_11275, signal_4066}), .c ({signal_11428, signal_3686}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_108 ( .s (signal_13468), .b ({signal_10496, signal_4458}), .a ({signal_11568, signal_4065}), .c ({signal_11584, signal_3685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_13468), .b ({signal_10306, signal_3936}), .a ({signal_11098, signal_4064}), .c ({signal_11189, signal_3684}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_110 ( .s (signal_13468), .b ({signal_10305, signal_3935}), .a ({signal_11358, signal_4063}), .c ({signal_11429, signal_3683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_111 ( .s (signal_13468), .b ({signal_10528, signal_4510}), .a ({signal_11311, signal_4117}), .c ({signal_11430, signal_3737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_13468), .b ({signal_10304, signal_4455}), .a ({signal_11357, signal_4062}), .c ({signal_11431, signal_3682}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_113 ( .s (signal_13468), .b ({signal_10495, signal_4454}), .a ({signal_11302, signal_4061}), .c ({signal_11432, signal_3681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_114 ( .s (signal_13468), .b ({signal_10494, signal_4453}), .a ({signal_11301, signal_4060}), .c ({signal_11433, signal_3680}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_115 ( .s (signal_13468), .b ({signal_10301, signal_4460}), .a ({signal_11092, signal_4059}), .c ({signal_11190, signal_3679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_116 ( .s (signal_13468), .b ({signal_10332, signal_3930}), .a ({signal_11297, signal_4058}), .c ({signal_11434, signal_3678}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_117 ( .s (signal_13468), .b ({signal_10547, signal_4450}), .a ({signal_11565, signal_4057}), .c ({signal_11585, signal_3677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_118 ( .s (signal_13468), .b ({signal_10416, signal_3928}), .a ({signal_11063, signal_4056}), .c ({signal_11191, signal_3676}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_119 ( .s (signal_13468), .b ({signal_10415, signal_3927}), .a ({signal_11344, signal_4055}), .c ({signal_11435, signal_3675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_120 ( .s (signal_13460), .b ({signal_10414, signal_4447}), .a ({signal_11343, signal_4054}), .c ({signal_11436, signal_3674}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_13460), .b ({signal_10546, signal_4446}), .a ({signal_11289, signal_4053}), .c ({signal_11437, signal_3673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_122 ( .s (signal_13460), .b ({signal_10527, signal_4509}), .a ({signal_11310, signal_4116}), .c ({signal_11438, signal_3736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_123 ( .s (signal_13460), .b ({signal_10545, signal_4445}), .a ({signal_11288, signal_4052}), .c ({signal_11439, signal_3672}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_13460), .b ({signal_10411, signal_4452}), .a ({signal_11056, signal_4051}), .c ({signal_11192, signal_3671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_125 ( .s (signal_13460), .b ({signal_10323, signal_3922}), .a ({signal_11287, signal_4050}), .c ({signal_11440, signal_3670}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_126 ( .s (signal_13460), .b ({signal_10520, signal_4442}), .a ({signal_11563, signal_4049}), .c ({signal_11586, signal_3669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_127 ( .s (signal_13460), .b ({signal_10353, signal_3920}), .a ({signal_11083, signal_4048}), .c ({signal_11193, signal_3668}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_128 ( .s (signal_13460), .b ({signal_10352, signal_3919}), .a ({signal_11353, signal_4047}), .c ({signal_11441, signal_3667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_129 ( .s (signal_13460), .b ({signal_10351, signal_4439}), .a ({signal_11352, signal_4046}), .c ({signal_11442, signal_3666}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_130 ( .s (signal_13460), .b ({signal_10519, signal_4438}), .a ({signal_11296, signal_4045}), .c ({signal_11443, signal_3665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_131 ( .s (signal_13460), .b ({signal_10518, signal_4437}), .a ({signal_11295, signal_4044}), .c ({signal_11444, signal_3664}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_132 ( .s (signal_13452), .b ({signal_10348, signal_4444}), .a ({signal_11078, signal_4043}), .c ({signal_11194, signal_3663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_13452), .b ({signal_10369, signal_4516}), .a ({signal_11118, signal_4115}), .c ({signal_11195, signal_3735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_134 ( .s (signal_13452), .b ({signal_10328, signal_3914}), .a ({signal_11294, signal_4042}), .c ({signal_11445, signal_3662}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_135 ( .s (signal_13452), .b ({signal_10535, signal_4434}), .a ({signal_11566, signal_4041}), .c ({signal_11587, signal_3661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_13452), .b ({signal_10388, signal_3912}), .a ({signal_11075, signal_4040}), .c ({signal_11196, signal_3660}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_137 ( .s (signal_13452), .b ({signal_10387, signal_3911}), .a ({signal_11350, signal_4039}), .c ({signal_11446, signal_3659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_138 ( .s (signal_13452), .b ({signal_10386, signal_4431}), .a ({signal_11348, signal_4038}), .c ({signal_11447, signal_3658}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_139 ( .s (signal_13452), .b ({signal_10534, signal_4430}), .a ({signal_11293, signal_4037}), .c ({signal_11448, signal_3657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_140 ( .s (signal_13452), .b ({signal_10533, signal_4429}), .a ({signal_11292, signal_4036}), .c ({signal_11449, signal_3656}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_141 ( .s (signal_13452), .b ({signal_10383, signal_4436}), .a ({signal_11069, signal_4035}), .c ({signal_11197, signal_3655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_142 ( .s (signal_13452), .b ({signal_10299, signal_3906}), .a ({signal_11274, signal_4034}), .c ({signal_11450, signal_3654}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_143 ( .s (signal_13452), .b ({signal_10499, signal_4426}), .a ({signal_11564, signal_4033}), .c ({signal_11588, signal_3653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_144 ( .s (signal_13444), .b ({signal_10330, signal_3986}), .a ({signal_11309, signal_4114}), .c ({signal_11451, signal_3734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_13444), .b ({signal_10313, signal_3904}), .a ({signal_11067, signal_4032}), .c ({signal_11198, signal_3652}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_146 ( .s (signal_13444), .b ({signal_10312, signal_3903}), .a ({signal_11346, signal_4031}), .c ({signal_11452, signal_3651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_147 ( .s (signal_13444), .b ({signal_10311, signal_4423}), .a ({signal_11345, signal_4030}), .c ({signal_11453, signal_3650}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_13444), .b ({signal_10498, signal_4422}), .a ({signal_11291, signal_4029}), .c ({signal_11454, signal_3649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_149 ( .s (signal_13444), .b ({signal_10497, signal_4421}), .a ({signal_11290, signal_4028}), .c ({signal_11455, signal_3648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_150 ( .s (signal_13444), .b ({signal_10308, signal_4428}), .a ({signal_11061, signal_4027}), .c ({signal_11199, signal_3647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_151 ( .s (signal_13444), .b ({signal_10322, signal_3898}), .a ({signal_11286, signal_4026}), .c ({signal_11456, signal_3646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_152 ( .s (signal_13444), .b ({signal_10517, signal_4418}), .a ({signal_11561, signal_4025}), .c ({signal_11589, signal_3645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_153 ( .s (signal_13444), .b ({signal_10346, signal_3896}), .a ({signal_11032, signal_4024}), .c ({signal_11200, signal_3644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_154 ( .s (signal_13444), .b ({signal_10345, signal_3895}), .a ({signal_11332, signal_4023}), .c ({signal_11457, signal_3643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_155 ( .s (signal_13444), .b ({signal_10541, signal_4506}), .a ({signal_11571, signal_4113}), .c ({signal_11590, signal_3733}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_291 ( .s (signal_13492), .b ({signal_11378, signal_3742}), .a ({signal_13508, signal_13500}), .c ({signal_11592, signal_421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_294 ( .s (signal_13492), .b ({signal_11579, signal_3741}), .a ({signal_13524, signal_13516}), .c ({signal_11758, signal_423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_297 ( .s (signal_13492), .b ({signal_11181, signal_3740}), .a ({signal_13540, signal_13532}), .c ({signal_11459, signal_425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_300 ( .s (signal_13492), .b ({signal_11416, signal_3739}), .a ({signal_13556, signal_13548}), .c ({signal_11594, signal_427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_303 ( .s (signal_13492), .b ({signal_11423, signal_3738}), .a ({signal_13572, signal_13564}), .c ({signal_11596, signal_429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_306 ( .s (signal_13492), .b ({signal_11430, signal_3737}), .a ({signal_13588, signal_13580}), .c ({signal_11598, signal_431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_309 ( .s (signal_13492), .b ({signal_11438, signal_3736}), .a ({signal_13604, signal_13596}), .c ({signal_11600, signal_433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_312 ( .s (signal_13492), .b ({signal_11195, signal_3735}), .a ({signal_13620, signal_13612}), .c ({signal_11461, signal_435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_315 ( .s (signal_13492), .b ({signal_11451, signal_3734}), .a ({signal_13636, signal_13628}), .c ({signal_11602, signal_437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_318 ( .s (signal_13492), .b ({signal_11590, signal_3733}), .a ({signal_13652, signal_13644}), .c ({signal_11760, signal_439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_321 ( .s (signal_13492), .b ({signal_11171, signal_3732}), .a ({signal_13668, signal_13660}), .c ({signal_11463, signal_441}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_324 ( .s (signal_13492), .b ({signal_11392, signal_3731}), .a ({signal_13684, signal_13676}), .c ({signal_11604, signal_443}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_327 ( .s (signal_13492), .b ({signal_11398, signal_3730}), .a ({signal_13700, signal_13692}), .c ({signal_11606, signal_445}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_330 ( .s (signal_13492), .b ({signal_11399, signal_3729}), .a ({signal_13716, signal_13708}), .c ({signal_11608, signal_447}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_333 ( .s (signal_13492), .b ({signal_11400, signal_3728}), .a ({signal_13732, signal_13724}), .c ({signal_11610, signal_449}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_336 ( .s (signal_13492), .b ({signal_11177, signal_3727}), .a ({signal_13748, signal_13740}), .c ({signal_11465, signal_451}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_339 ( .s (signal_13492), .b ({signal_11401, signal_3726}), .a ({signal_13764, signal_13756}), .c ({signal_11612, signal_453}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_342 ( .s (signal_13492), .b ({signal_11578, signal_3725}), .a ({signal_13780, signal_13772}), .c ({signal_11762, signal_455}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_345 ( .s (signal_13492), .b ({signal_11178, signal_3724}), .a ({signal_13796, signal_13788}), .c ({signal_11467, signal_457}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_348 ( .s (signal_13492), .b ({signal_11402, signal_3723}), .a ({signal_13812, signal_13804}), .c ({signal_11614, signal_459}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_351 ( .s (signal_13492), .b ({signal_11403, signal_3722}), .a ({signal_13828, signal_13820}), .c ({signal_11616, signal_461}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_354 ( .s (signal_13492), .b ({signal_11404, signal_3721}), .a ({signal_13844, signal_13836}), .c ({signal_11618, signal_463}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_357 ( .s (signal_13492), .b ({signal_11405, signal_3720}), .a ({signal_13860, signal_13852}), .c ({signal_11620, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_360 ( .s (signal_13492), .b ({signal_11179, signal_3719}), .a ({signal_13876, signal_13868}), .c ({signal_11469, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_363 ( .s (signal_13492), .b ({signal_11406, signal_3718}), .a ({signal_13892, signal_13884}), .c ({signal_11622, signal_469}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_366 ( .s (signal_13492), .b ({signal_11580, signal_3717}), .a ({signal_13908, signal_13900}), .c ({signal_11764, signal_471}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_369 ( .s (signal_13492), .b ({signal_11180, signal_3716}), .a ({signal_13924, signal_13916}), .c ({signal_11471, signal_473}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_372 ( .s (signal_13492), .b ({signal_11407, signal_3715}), .a ({signal_13940, signal_13932}), .c ({signal_11624, signal_475}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_375 ( .s (signal_13492), .b ({signal_11408, signal_3714}), .a ({signal_13956, signal_13948}), .c ({signal_11626, signal_477}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_378 ( .s (signal_13492), .b ({signal_11409, signal_3713}), .a ({signal_13972, signal_13964}), .c ({signal_11628, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_381 ( .s (signal_13492), .b ({signal_11410, signal_3712}), .a ({signal_13988, signal_13980}), .c ({signal_11630, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_384 ( .s (signal_13492), .b ({signal_11182, signal_3711}), .a ({signal_14004, signal_13996}), .c ({signal_11473, signal_483}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_387 ( .s (signal_13492), .b ({signal_11411, signal_3710}), .a ({signal_14020, signal_14012}), .c ({signal_11632, signal_485}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_390 ( .s (signal_13492), .b ({signal_11581, signal_3709}), .a ({signal_14036, signal_14028}), .c ({signal_11766, signal_487}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_393 ( .s (signal_13492), .b ({signal_11183, signal_3708}), .a ({signal_14052, signal_14044}), .c ({signal_11475, signal_489}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_396 ( .s (signal_13492), .b ({signal_11412, signal_3707}), .a ({signal_14068, signal_14060}), .c ({signal_11634, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_399 ( .s (signal_13492), .b ({signal_11413, signal_3706}), .a ({signal_14084, signal_14076}), .c ({signal_11636, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_402 ( .s (signal_13492), .b ({signal_11414, signal_3705}), .a ({signal_14100, signal_14092}), .c ({signal_11638, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_405 ( .s (signal_13492), .b ({signal_11415, signal_3704}), .a ({signal_14116, signal_14108}), .c ({signal_11640, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_408 ( .s (signal_13492), .b ({signal_11184, signal_3703}), .a ({signal_14132, signal_14124}), .c ({signal_11477, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_411 ( .s (signal_13492), .b ({signal_11417, signal_3702}), .a ({signal_14148, signal_14140}), .c ({signal_11642, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_414 ( .s (signal_13492), .b ({signal_11582, signal_3701}), .a ({signal_14164, signal_14156}), .c ({signal_11768, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_417 ( .s (signal_13492), .b ({signal_11185, signal_3700}), .a ({signal_14180, signal_14172}), .c ({signal_11479, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_420 ( .s (signal_13492), .b ({signal_11418, signal_3699}), .a ({signal_14196, signal_14188}), .c ({signal_11644, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_423 ( .s (signal_13492), .b ({signal_11419, signal_3698}), .a ({signal_14212, signal_14204}), .c ({signal_11646, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_426 ( .s (signal_13492), .b ({signal_11420, signal_3697}), .a ({signal_14228, signal_14220}), .c ({signal_11648, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_429 ( .s (signal_13492), .b ({signal_11421, signal_3696}), .a ({signal_14244, signal_14236}), .c ({signal_11650, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_432 ( .s (signal_13492), .b ({signal_11186, signal_3695}), .a ({signal_14260, signal_14252}), .c ({signal_11481, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_435 ( .s (signal_13492), .b ({signal_11422, signal_3694}), .a ({signal_14276, signal_14268}), .c ({signal_11652, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_438 ( .s (signal_13492), .b ({signal_11583, signal_3693}), .a ({signal_14292, signal_14284}), .c ({signal_11770, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_441 ( .s (signal_13492), .b ({signal_11187, signal_3692}), .a ({signal_14308, signal_14300}), .c ({signal_11483, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_444 ( .s (signal_13492), .b ({signal_11424, signal_3691}), .a ({signal_14324, signal_14316}), .c ({signal_11654, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_447 ( .s (signal_13492), .b ({signal_11425, signal_3690}), .a ({signal_14340, signal_14332}), .c ({signal_11656, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_450 ( .s (signal_13492), .b ({signal_11426, signal_3689}), .a ({signal_14356, signal_14348}), .c ({signal_11658, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_453 ( .s (signal_13492), .b ({signal_11427, signal_3688}), .a ({signal_14372, signal_14364}), .c ({signal_11660, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_456 ( .s (signal_13492), .b ({signal_11188, signal_3687}), .a ({signal_14388, signal_14380}), .c ({signal_11485, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_459 ( .s (signal_13492), .b ({signal_11428, signal_3686}), .a ({signal_14404, signal_14396}), .c ({signal_11662, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_462 ( .s (signal_13492), .b ({signal_11584, signal_3685}), .a ({signal_14420, signal_14412}), .c ({signal_11772, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_465 ( .s (signal_13492), .b ({signal_11189, signal_3684}), .a ({signal_14436, signal_14428}), .c ({signal_11487, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_468 ( .s (signal_13492), .b ({signal_11429, signal_3683}), .a ({signal_14452, signal_14444}), .c ({signal_11664, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_471 ( .s (signal_13492), .b ({signal_11431, signal_3682}), .a ({signal_14468, signal_14460}), .c ({signal_11666, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_474 ( .s (signal_13492), .b ({signal_11432, signal_3681}), .a ({signal_14484, signal_14476}), .c ({signal_11668, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_477 ( .s (signal_13492), .b ({signal_11433, signal_3680}), .a ({signal_14500, signal_14492}), .c ({signal_11670, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_480 ( .s (signal_13492), .b ({signal_11190, signal_3679}), .a ({signal_14516, signal_14508}), .c ({signal_11489, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_483 ( .s (signal_13492), .b ({signal_11434, signal_3678}), .a ({signal_14532, signal_14524}), .c ({signal_11672, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_486 ( .s (signal_13492), .b ({signal_11585, signal_3677}), .a ({signal_14548, signal_14540}), .c ({signal_11774, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_489 ( .s (signal_13492), .b ({signal_11191, signal_3676}), .a ({signal_14564, signal_14556}), .c ({signal_11491, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_492 ( .s (signal_13492), .b ({signal_11435, signal_3675}), .a ({signal_14580, signal_14572}), .c ({signal_11674, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_495 ( .s (signal_13492), .b ({signal_11436, signal_3674}), .a ({signal_14596, signal_14588}), .c ({signal_11676, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_498 ( .s (signal_13492), .b ({signal_11437, signal_3673}), .a ({signal_14612, signal_14604}), .c ({signal_11678, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_501 ( .s (signal_13492), .b ({signal_11439, signal_3672}), .a ({signal_14628, signal_14620}), .c ({signal_11680, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_504 ( .s (signal_13492), .b ({signal_11192, signal_3671}), .a ({signal_14644, signal_14636}), .c ({signal_11493, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_507 ( .s (signal_13492), .b ({signal_11440, signal_3670}), .a ({signal_14660, signal_14652}), .c ({signal_11682, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_510 ( .s (signal_13492), .b ({signal_11586, signal_3669}), .a ({signal_14676, signal_14668}), .c ({signal_11776, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_513 ( .s (signal_13492), .b ({signal_11193, signal_3668}), .a ({signal_14692, signal_14684}), .c ({signal_11495, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_516 ( .s (signal_13492), .b ({signal_11441, signal_3667}), .a ({signal_14708, signal_14700}), .c ({signal_11684, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_519 ( .s (signal_13492), .b ({signal_11442, signal_3666}), .a ({signal_14724, signal_14716}), .c ({signal_11686, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_522 ( .s (signal_13492), .b ({signal_11443, signal_3665}), .a ({signal_14740, signal_14732}), .c ({signal_11688, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_525 ( .s (signal_13492), .b ({signal_11444, signal_3664}), .a ({signal_14756, signal_14748}), .c ({signal_11690, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_528 ( .s (signal_13492), .b ({signal_11194, signal_3663}), .a ({signal_14772, signal_14764}), .c ({signal_11497, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_531 ( .s (signal_13492), .b ({signal_11445, signal_3662}), .a ({signal_14788, signal_14780}), .c ({signal_11692, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_534 ( .s (signal_13492), .b ({signal_11587, signal_3661}), .a ({signal_14804, signal_14796}), .c ({signal_11778, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_537 ( .s (signal_13492), .b ({signal_11196, signal_3660}), .a ({signal_14820, signal_14812}), .c ({signal_11499, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_540 ( .s (signal_13492), .b ({signal_11446, signal_3659}), .a ({signal_14836, signal_14828}), .c ({signal_11694, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_543 ( .s (signal_13492), .b ({signal_11447, signal_3658}), .a ({signal_14852, signal_14844}), .c ({signal_11696, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_546 ( .s (signal_13492), .b ({signal_11448, signal_3657}), .a ({signal_14868, signal_14860}), .c ({signal_11698, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_549 ( .s (signal_13492), .b ({signal_11449, signal_3656}), .a ({signal_14884, signal_14876}), .c ({signal_11700, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_552 ( .s (signal_13492), .b ({signal_11197, signal_3655}), .a ({signal_14900, signal_14892}), .c ({signal_11501, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_555 ( .s (signal_13492), .b ({signal_11450, signal_3654}), .a ({signal_14916, signal_14908}), .c ({signal_11702, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_558 ( .s (signal_13492), .b ({signal_11588, signal_3653}), .a ({signal_14932, signal_14924}), .c ({signal_11780, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_561 ( .s (signal_13492), .b ({signal_11198, signal_3652}), .a ({signal_14948, signal_14940}), .c ({signal_11503, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_564 ( .s (signal_13492), .b ({signal_11452, signal_3651}), .a ({signal_14964, signal_14956}), .c ({signal_11704, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_567 ( .s (signal_13492), .b ({signal_11453, signal_3650}), .a ({signal_14980, signal_14972}), .c ({signal_11706, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_570 ( .s (signal_13492), .b ({signal_11454, signal_3649}), .a ({signal_14996, signal_14988}), .c ({signal_11708, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_573 ( .s (signal_13492), .b ({signal_11455, signal_3648}), .a ({signal_15012, signal_15004}), .c ({signal_11710, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_576 ( .s (signal_13492), .b ({signal_11199, signal_3647}), .a ({signal_15028, signal_15020}), .c ({signal_11505, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_579 ( .s (signal_13492), .b ({signal_11456, signal_3646}), .a ({signal_15044, signal_15036}), .c ({signal_11712, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_582 ( .s (signal_13492), .b ({signal_11589, signal_3645}), .a ({signal_15060, signal_15052}), .c ({signal_11782, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_585 ( .s (signal_13492), .b ({signal_11200, signal_3644}), .a ({signal_15076, signal_15068}), .c ({signal_11507, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_588 ( .s (signal_13492), .b ({signal_11457, signal_3643}), .a ({signal_15092, signal_15084}), .c ({signal_11714, signal_619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_591 ( .s (signal_13492), .b ({signal_11379, signal_3642}), .a ({signal_15108, signal_15100}), .c ({signal_11716, signal_621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_594 ( .s (signal_13492), .b ({signal_11380, signal_3641}), .a ({signal_15124, signal_15116}), .c ({signal_11718, signal_623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_597 ( .s (signal_13492), .b ({signal_11381, signal_3640}), .a ({signal_15140, signal_15132}), .c ({signal_11720, signal_625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_600 ( .s (signal_13492), .b ({signal_11169, signal_3639}), .a ({signal_15156, signal_15148}), .c ({signal_11509, signal_627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_603 ( .s (signal_13492), .b ({signal_11382, signal_3638}), .a ({signal_15172, signal_15164}), .c ({signal_11722, signal_629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_606 ( .s (signal_13492), .b ({signal_11575, signal_3637}), .a ({signal_15188, signal_15180}), .c ({signal_11784, signal_631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_609 ( .s (signal_13492), .b ({signal_11170, signal_3636}), .a ({signal_15204, signal_15196}), .c ({signal_11511, signal_633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_612 ( .s (signal_13492), .b ({signal_11383, signal_3635}), .a ({signal_15220, signal_15212}), .c ({signal_11724, signal_635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_615 ( .s (signal_13492), .b ({signal_11384, signal_3634}), .a ({signal_15236, signal_15228}), .c ({signal_11726, signal_637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_618 ( .s (signal_13492), .b ({signal_11385, signal_3633}), .a ({signal_15252, signal_15244}), .c ({signal_11728, signal_639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_621 ( .s (signal_13492), .b ({signal_11386, signal_3632}), .a ({signal_15268, signal_15260}), .c ({signal_11730, signal_641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_624 ( .s (signal_13492), .b ({signal_11172, signal_3631}), .a ({signal_15284, signal_15276}), .c ({signal_11513, signal_643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_627 ( .s (signal_13492), .b ({signal_11387, signal_3630}), .a ({signal_15300, signal_15292}), .c ({signal_11732, signal_645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_630 ( .s (signal_13492), .b ({signal_11576, signal_3629}), .a ({signal_15316, signal_15308}), .c ({signal_11786, signal_647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_633 ( .s (signal_13492), .b ({signal_11173, signal_3628}), .a ({signal_15332, signal_15324}), .c ({signal_11515, signal_649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_636 ( .s (signal_13492), .b ({signal_11388, signal_3627}), .a ({signal_15348, signal_15340}), .c ({signal_11734, signal_651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_639 ( .s (signal_13492), .b ({signal_11389, signal_3626}), .a ({signal_15364, signal_15356}), .c ({signal_11736, signal_653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_642 ( .s (signal_13492), .b ({signal_11390, signal_3625}), .a ({signal_15380, signal_15372}), .c ({signal_11738, signal_655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_645 ( .s (signal_13492), .b ({signal_11391, signal_3624}), .a ({signal_15396, signal_15388}), .c ({signal_11740, signal_657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_648 ( .s (signal_13492), .b ({signal_11174, signal_3623}), .a ({signal_15412, signal_15404}), .c ({signal_11517, signal_659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_651 ( .s (signal_13492), .b ({signal_11393, signal_3622}), .a ({signal_15428, signal_15420}), .c ({signal_11742, signal_661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_654 ( .s (signal_13492), .b ({signal_11577, signal_3621}), .a ({signal_15444, signal_15436}), .c ({signal_11788, signal_663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_657 ( .s (signal_13492), .b ({signal_11175, signal_3620}), .a ({signal_15460, signal_15452}), .c ({signal_11519, signal_665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_660 ( .s (signal_13492), .b ({signal_11394, signal_3619}), .a ({signal_15476, signal_15468}), .c ({signal_11744, signal_667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_663 ( .s (signal_13492), .b ({signal_11395, signal_3618}), .a ({signal_15492, signal_15484}), .c ({signal_11746, signal_669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_666 ( .s (signal_13492), .b ({signal_11396, signal_3617}), .a ({signal_15508, signal_15500}), .c ({signal_11748, signal_671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_669 ( .s (signal_13492), .b ({signal_11397, signal_3616}), .a ({signal_15524, signal_15516}), .c ({signal_11750, signal_673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_672 ( .s (signal_13492), .b ({signal_11176, signal_3615}), .a ({signal_15540, signal_15532}), .c ({signal_11521, signal_675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3155 ( .s (signal_13492), .b ({signal_11022, signal_4250}), .a ({signal_15556, signal_15548}), .c ({signal_11202, signal_2853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3158 ( .s (signal_13492), .b ({signal_11326, signal_4249}), .a ({signal_15572, signal_15564}), .c ({signal_11523, signal_2855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3161 ( .s (signal_13492), .b ({signal_11154, signal_4248}), .a ({signal_15588, signal_15580}), .c ({signal_11204, signal_2857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3164 ( .s (signal_13492), .b ({signal_11153, signal_4247}), .a ({signal_15604, signal_15596}), .c ({signal_11206, signal_2859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3167 ( .s (signal_13492), .b ({signal_11152, signal_4246}), .a ({signal_15620, signal_15612}), .c ({signal_11208, signal_2861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3170 ( .s (signal_13492), .b ({signal_11323, signal_4245}), .a ({signal_15636, signal_15628}), .c ({signal_11525, signal_2863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3173 ( .s (signal_13492), .b ({signal_11322, signal_4244}), .a ({signal_15652, signal_15644}), .c ({signal_11527, signal_2865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3176 ( .s (signal_13492), .b ({signal_11149, signal_4243}), .a ({signal_15668, signal_15660}), .c ({signal_11210, signal_2867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3179 ( .s (signal_13492), .b ({signal_11011, signal_4242}), .a ({signal_15684, signal_15676}), .c ({signal_11212, signal_2869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3182 ( .s (signal_13492), .b ({signal_11321, signal_4241}), .a ({signal_15700, signal_15692}), .c ({signal_11529, signal_2871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3185 ( .s (signal_13492), .b ({signal_11168, signal_4240}), .a ({signal_15716, signal_15708}), .c ({signal_11214, signal_2873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3188 ( .s (signal_13492), .b ({signal_11167, signal_4239}), .a ({signal_15732, signal_15724}), .c ({signal_11216, signal_2875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3191 ( .s (signal_13492), .b ({signal_11166, signal_4238}), .a ({signal_15748, signal_15740}), .c ({signal_11218, signal_2877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3194 ( .s (signal_13492), .b ({signal_11329, signal_4237}), .a ({signal_15764, signal_15756}), .c ({signal_11531, signal_2879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3197 ( .s (signal_13492), .b ({signal_11328, signal_4236}), .a ({signal_15780, signal_15772}), .c ({signal_11533, signal_2881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3200 ( .s (signal_13492), .b ({signal_11163, signal_4235}), .a ({signal_15796, signal_15788}), .c ({signal_11220, signal_2883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3203 ( .s (signal_13492), .b ({signal_11019, signal_4234}), .a ({signal_15812, signal_15804}), .c ({signal_11222, signal_2885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3206 ( .s (signal_13492), .b ({signal_11327, signal_4233}), .a ({signal_15828, signal_15820}), .c ({signal_11535, signal_2887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3209 ( .s (signal_13492), .b ({signal_11161, signal_4232}), .a ({signal_15844, signal_15836}), .c ({signal_11224, signal_2889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3212 ( .s (signal_13492), .b ({signal_11160, signal_4231}), .a ({signal_15860, signal_15852}), .c ({signal_11226, signal_2891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3215 ( .s (signal_13492), .b ({signal_11158, signal_4230}), .a ({signal_15876, signal_15868}), .c ({signal_11228, signal_2893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3218 ( .s (signal_13492), .b ({signal_11325, signal_4229}), .a ({signal_15892, signal_15884}), .c ({signal_11537, signal_2895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3221 ( .s (signal_13492), .b ({signal_11324, signal_4228}), .a ({signal_15908, signal_15900}), .c ({signal_11539, signal_2897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3224 ( .s (signal_13492), .b ({signal_11155, signal_4227}), .a ({signal_15924, signal_15916}), .c ({signal_11230, signal_2899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3227 ( .s (signal_13492), .b ({signal_11272, signal_4226}), .a ({signal_15940, signal_15932}), .c ({signal_11541, signal_2901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3230 ( .s (signal_13492), .b ({signal_11558, signal_4225}), .a ({signal_15956, signal_15948}), .c ({signal_11752, signal_2903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3233 ( .s (signal_13492), .b ({signal_11270, signal_4224}), .a ({signal_15972, signal_15964}), .c ({signal_11543, signal_2905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3236 ( .s (signal_13492), .b ({signal_11269, signal_4223}), .a ({signal_15988, signal_15980}), .c ({signal_11545, signal_2907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3239 ( .s (signal_13492), .b ({signal_11268, signal_4222}), .a ({signal_16004, signal_15996}), .c ({signal_11547, signal_2909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3242 ( .s (signal_13492), .b ({signal_11557, signal_4221}), .a ({signal_16020, signal_16012}), .c ({signal_11754, signal_2911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3245 ( .s (signal_13492), .b ({signal_11556, signal_4220}), .a ({signal_16036, signal_16028}), .c ({signal_11756, signal_2913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3248 ( .s (signal_13492), .b ({signal_11265, signal_4219}), .a ({signal_16052, signal_16044}), .c ({signal_11549, signal_2915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3251 ( .s (signal_13492), .b ({signal_10795, signal_4218}), .a ({signal_16068, signal_16060}), .c ({signal_10937, signal_2917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3254 ( .s (signal_13492), .b ({signal_11017, signal_4217}), .a ({signal_16084, signal_16076}), .c ({signal_11232, signal_2919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3257 ( .s (signal_13492), .b ({signal_10919, signal_4216}), .a ({signal_16100, signal_16092}), .c ({signal_10939, signal_2921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3260 ( .s (signal_13492), .b ({signal_10918, signal_4215}), .a ({signal_16116, signal_16108}), .c ({signal_10941, signal_2923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3263 ( .s (signal_13492), .b ({signal_10917, signal_4214}), .a ({signal_16132, signal_16124}), .c ({signal_10943, signal_2925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3266 ( .s (signal_13492), .b ({signal_11014, signal_4213}), .a ({signal_16148, signal_16140}), .c ({signal_11234, signal_2927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3269 ( .s (signal_13492), .b ({signal_11013, signal_4212}), .a ({signal_16164, signal_16156}), .c ({signal_11236, signal_2929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3272 ( .s (signal_13492), .b ({signal_10914, signal_4211}), .a ({signal_16180, signal_16172}), .c ({signal_10945, signal_2931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3275 ( .s (signal_13492), .b ({signal_10785, signal_4210}), .a ({signal_16196, signal_16188}), .c ({signal_10947, signal_2933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3278 ( .s (signal_13492), .b ({signal_11012, signal_4209}), .a ({signal_16212, signal_16204}), .c ({signal_11238, signal_2935}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3281 ( .s (signal_13492), .b ({signal_10934, signal_4208}), .a ({signal_16228, signal_16220}), .c ({signal_10949, signal_2937}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3284 ( .s (signal_13492), .b ({signal_10933, signal_4207}), .a ({signal_16244, signal_16236}), .c ({signal_10951, signal_2939}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3287 ( .s (signal_13492), .b ({signal_10932, signal_4206}), .a ({signal_16260, signal_16252}), .c ({signal_10953, signal_2941}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3290 ( .s (signal_13492), .b ({signal_11021, signal_4205}), .a ({signal_16276, signal_16268}), .c ({signal_11240, signal_2943}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3293 ( .s (signal_13492), .b ({signal_11020, signal_4204}), .a ({signal_16292, signal_16284}), .c ({signal_11242, signal_2945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3296 ( .s (signal_13492), .b ({signal_10929, signal_4203}), .a ({signal_16308, signal_16300}), .c ({signal_10955, signal_2947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3299 ( .s (signal_13492), .b ({signal_10792, signal_4202}), .a ({signal_16324, signal_16316}), .c ({signal_10957, signal_2949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3302 ( .s (signal_13492), .b ({signal_11018, signal_4201}), .a ({signal_16340, signal_16332}), .c ({signal_11244, signal_2951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3305 ( .s (signal_13492), .b ({signal_10926, signal_4200}), .a ({signal_16356, signal_16348}), .c ({signal_10959, signal_2953}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3308 ( .s (signal_13492), .b ({signal_10925, signal_4199}), .a ({signal_16372, signal_16364}), .c ({signal_10961, signal_2955}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3311 ( .s (signal_13492), .b ({signal_10923, signal_4198}), .a ({signal_16388, signal_16380}), .c ({signal_10963, signal_2957}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3314 ( .s (signal_13492), .b ({signal_11016, signal_4197}), .a ({signal_16404, signal_16396}), .c ({signal_11246, signal_2959}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3317 ( .s (signal_13492), .b ({signal_11015, signal_4196}), .a ({signal_16420, signal_16412}), .c ({signal_11248, signal_2961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3320 ( .s (signal_13492), .b ({signal_10920, signal_4195}), .a ({signal_16436, signal_16428}), .c ({signal_10965, signal_2963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3323 ( .s (signal_13492), .b ({signal_11007, signal_4194}), .a ({signal_16452, signal_16444}), .c ({signal_11250, signal_2965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3326 ( .s (signal_13492), .b ({signal_11271, signal_4193}), .a ({signal_16468, signal_16460}), .c ({signal_11551, signal_2967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3329 ( .s (signal_13492), .b ({signal_11005, signal_4192}), .a ({signal_16484, signal_16476}), .c ({signal_11252, signal_2969}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3332 ( .s (signal_13492), .b ({signal_11004, signal_4191}), .a ({signal_16500, signal_16492}), .c ({signal_11254, signal_2971}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3335 ( .s (signal_13492), .b ({signal_11003, signal_4190}), .a ({signal_16516, signal_16508}), .c ({signal_11256, signal_2973}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3338 ( .s (signal_13492), .b ({signal_11267, signal_4189}), .a ({signal_16532, signal_16524}), .c ({signal_11553, signal_2975}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3341 ( .s (signal_13492), .b ({signal_11266, signal_4188}), .a ({signal_16548, signal_16540}), .c ({signal_11555, signal_2977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3344 ( .s (signal_13492), .b ({signal_11000, signal_4187}), .a ({signal_16564, signal_16556}), .c ({signal_11258, signal_2979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3347 ( .s (signal_13492), .b ({signal_10565, signal_4186}), .a ({signal_16580, signal_16572}), .c ({signal_10707, signal_2981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3350 ( .s (signal_13492), .b ({signal_10790, signal_4185}), .a ({signal_16596, signal_16588}), .c ({signal_10967, signal_2983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3353 ( .s (signal_13492), .b ({signal_10689, signal_4184}), .a ({signal_16612, signal_16604}), .c ({signal_10709, signal_2985}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3356 ( .s (signal_13492), .b ({signal_10688, signal_4183}), .a ({signal_16628, signal_16620}), .c ({signal_10711, signal_2987}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3359 ( .s (signal_13492), .b ({signal_10687, signal_4182}), .a ({signal_16644, signal_16636}), .c ({signal_10713, signal_2989}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3362 ( .s (signal_13492), .b ({signal_10787, signal_4181}), .a ({signal_16660, signal_16652}), .c ({signal_10969, signal_2991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3365 ( .s (signal_13492), .b ({signal_10786, signal_4180}), .a ({signal_16676, signal_16668}), .c ({signal_10971, signal_2993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3368 ( .s (signal_13492), .b ({signal_10684, signal_4179}), .a ({signal_16692, signal_16684}), .c ({signal_10715, signal_2995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3371 ( .s (signal_13492), .b ({signal_10554, signal_4178}), .a ({signal_16708, signal_16700}), .c ({signal_10717, signal_2997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3374 ( .s (signal_13492), .b ({signal_10784, signal_4177}), .a ({signal_16724, signal_16716}), .c ({signal_10973, signal_2999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3377 ( .s (signal_13492), .b ({signal_10704, signal_4176}), .a ({signal_16740, signal_16732}), .c ({signal_10719, signal_3001}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3380 ( .s (signal_13492), .b ({signal_10703, signal_4175}), .a ({signal_16756, signal_16748}), .c ({signal_10721, signal_3003}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3383 ( .s (signal_13492), .b ({signal_10702, signal_4174}), .a ({signal_16772, signal_16764}), .c ({signal_10723, signal_3005}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3386 ( .s (signal_13492), .b ({signal_10794, signal_4173}), .a ({signal_16788, signal_16780}), .c ({signal_10975, signal_3007}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3389 ( .s (signal_13492), .b ({signal_10793, signal_4172}), .a ({signal_16804, signal_16796}), .c ({signal_10977, signal_3009}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3392 ( .s (signal_13492), .b ({signal_10699, signal_4171}), .a ({signal_16820, signal_16812}), .c ({signal_10725, signal_3011}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3395 ( .s (signal_13492), .b ({signal_10556, signal_4170}), .a ({signal_16836, signal_16828}), .c ({signal_10727, signal_3013}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3398 ( .s (signal_13492), .b ({signal_10791, signal_4169}), .a ({signal_16852, signal_16844}), .c ({signal_10979, signal_3015}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3401 ( .s (signal_13492), .b ({signal_10696, signal_4168}), .a ({signal_16868, signal_16860}), .c ({signal_10729, signal_3017}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3404 ( .s (signal_13492), .b ({signal_10695, signal_4167}), .a ({signal_16884, signal_16876}), .c ({signal_10731, signal_3019}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3407 ( .s (signal_13492), .b ({signal_10693, signal_4166}), .a ({signal_16900, signal_16892}), .c ({signal_10733, signal_3021}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3410 ( .s (signal_13492), .b ({signal_10789, signal_4165}), .a ({signal_16916, signal_16908}), .c ({signal_10981, signal_3023}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3413 ( .s (signal_13492), .b ({signal_10788, signal_4164}), .a ({signal_16932, signal_16924}), .c ({signal_10983, signal_3025}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3416 ( .s (signal_13492), .b ({signal_10690, signal_4163}), .a ({signal_16948, signal_16940}), .c ({signal_10735, signal_3027}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3419 ( .s (signal_13492), .b ({signal_10768, signal_4162}), .a ({signal_16964, signal_16956}), .c ({signal_10985, signal_3029}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3422 ( .s (signal_13492), .b ({signal_11006, signal_4161}), .a ({signal_16980, signal_16972}), .c ({signal_11260, signal_3031}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3425 ( .s (signal_13492), .b ({signal_10767, signal_4160}), .a ({signal_16996, signal_16988}), .c ({signal_10987, signal_3033}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3428 ( .s (signal_13492), .b ({signal_10766, signal_4159}), .a ({signal_17012, signal_17004}), .c ({signal_10989, signal_3035}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3431 ( .s (signal_13492), .b ({signal_10765, signal_4158}), .a ({signal_17028, signal_17020}), .c ({signal_10991, signal_3037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3434 ( .s (signal_13492), .b ({signal_11002, signal_4157}), .a ({signal_17044, signal_17036}), .c ({signal_11262, signal_3039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3437 ( .s (signal_13492), .b ({signal_11001, signal_4156}), .a ({signal_17060, signal_17052}), .c ({signal_11264, signal_3041}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3440 ( .s (signal_13492), .b ({signal_10764, signal_4155}), .a ({signal_17076, signal_17068}), .c ({signal_10993, signal_3043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3443 ( .s (signal_13492), .b ({signal_10337, signal_4154}), .a ({signal_17092, signal_17084}), .c ({signal_10457, signal_3045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3446 ( .s (signal_13492), .b ({signal_10555, signal_4153}), .a ({signal_17108, signal_17100}), .c ({signal_10737, signal_3047}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3449 ( .s (signal_13492), .b ({signal_10434, signal_4152}), .a ({signal_17124, signal_17116}), .c ({signal_10459, signal_3049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3452 ( .s (signal_13492), .b ({signal_10433, signal_4151}), .a ({signal_17140, signal_17132}), .c ({signal_10461, signal_3051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3455 ( .s (signal_13492), .b ({signal_10454, signal_4150}), .a ({signal_17156, signal_17148}), .c ({signal_10463, signal_3053}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3458 ( .s (signal_13492), .b ({signal_10564, signal_4149}), .a ({signal_17172, signal_17164}), .c ({signal_10739, signal_3055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3461 ( .s (signal_13492), .b ({signal_10563, signal_4148}), .a ({signal_17188, signal_17180}), .c ({signal_10741, signal_3057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3464 ( .s (signal_13492), .b ({signal_10451, signal_4147}), .a ({signal_17204, signal_17196}), .c ({signal_10465, signal_3059}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3467 ( .s (signal_13492), .b ({signal_10336, signal_4146}), .a ({signal_17220, signal_17212}), .c ({signal_10467, signal_3061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3470 ( .s (signal_13492), .b ({signal_10562, signal_4145}), .a ({signal_17236, signal_17228}), .c ({signal_10743, signal_3063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3473 ( .s (signal_13492), .b ({signal_10449, signal_4144}), .a ({signal_17252, signal_17244}), .c ({signal_10469, signal_3065}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3476 ( .s (signal_13492), .b ({signal_10448, signal_4143}), .a ({signal_17268, signal_17260}), .c ({signal_10471, signal_3067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3479 ( .s (signal_13492), .b ({signal_10447, signal_4142}), .a ({signal_17284, signal_17276}), .c ({signal_10473, signal_3069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3482 ( .s (signal_13492), .b ({signal_10561, signal_4141}), .a ({signal_17300, signal_17292}), .c ({signal_10745, signal_3071}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3485 ( .s (signal_13492), .b ({signal_10560, signal_4140}), .a ({signal_17316, signal_17308}), .c ({signal_10747, signal_3073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3488 ( .s (signal_13492), .b ({signal_10444, signal_4139}), .a ({signal_17332, signal_17324}), .c ({signal_10475, signal_3075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3491 ( .s (signal_13492), .b ({signal_10335, signal_4138}), .a ({signal_17348, signal_17340}), .c ({signal_10477, signal_3077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3494 ( .s (signal_13492), .b ({signal_10559, signal_4137}), .a ({signal_17364, signal_17356}), .c ({signal_10749, signal_3079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3497 ( .s (signal_13492), .b ({signal_10442, signal_4136}), .a ({signal_17380, signal_17372}), .c ({signal_10479, signal_3081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3500 ( .s (signal_13492), .b ({signal_10441, signal_4135}), .a ({signal_17396, signal_17388}), .c ({signal_10481, signal_3083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3503 ( .s (signal_13492), .b ({signal_10440, signal_4134}), .a ({signal_17412, signal_17404}), .c ({signal_10483, signal_3085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3506 ( .s (signal_13492), .b ({signal_10558, signal_4133}), .a ({signal_17428, signal_17420}), .c ({signal_10751, signal_3087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3509 ( .s (signal_13492), .b ({signal_10557, signal_4132}), .a ({signal_17444, signal_17436}), .c ({signal_10753, signal_3089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3512 ( .s (signal_13492), .b ({signal_10437, signal_4131}), .a ({signal_17460, signal_17452}), .c ({signal_10485, signal_3091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3515 ( .s (signal_13492), .b ({signal_10490, signal_4130}), .a ({signal_17476, signal_17468}), .c ({signal_10755, signal_3093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3518 ( .s (signal_13492), .b ({signal_10771, signal_4129}), .a ({signal_17492, signal_17484}), .c ({signal_10995, signal_3095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3521 ( .s (signal_13492), .b ({signal_10489, signal_4128}), .a ({signal_17508, signal_17500}), .c ({signal_10757, signal_3097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3524 ( .s (signal_13492), .b ({signal_10488, signal_4127}), .a ({signal_17524, signal_17516}), .c ({signal_10759, signal_3099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3527 ( .s (signal_13492), .b ({signal_10487, signal_4126}), .a ({signal_17540, signal_17532}), .c ({signal_10761, signal_3101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3530 ( .s (signal_13492), .b ({signal_10770, signal_4125}), .a ({signal_17556, signal_17548}), .c ({signal_10997, signal_3103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3533 ( .s (signal_13492), .b ({signal_10769, signal_4124}), .a ({signal_17572, signal_17564}), .c ({signal_10999, signal_3105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3536 ( .s (signal_13492), .b ({signal_10486, signal_4123}), .a ({signal_17588, signal_17580}), .c ({signal_10763, signal_3107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3561 ( .a ({signal_17604, signal_17596}), .b ({signal_11000, signal_4187}), .c ({signal_11265, signal_4219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3562 ( .a ({signal_17620, signal_17612}), .b ({signal_10764, signal_4155}), .c ({signal_11000, signal_4187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3563 ( .a ({signal_17636, signal_17628}), .b ({signal_10486, signal_4123}), .c ({signal_10764, signal_4155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3564 ( .a ({signal_17652, signal_17644}), .b ({signal_11266, signal_4188}), .c ({signal_11556, signal_4220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3565 ( .a ({signal_17668, signal_17660}), .b ({signal_11001, signal_4156}), .c ({signal_11266, signal_4188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3566 ( .a ({signal_17684, signal_17676}), .b ({signal_10769, signal_4124}), .c ({signal_11001, signal_4156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3571 ( .a ({signal_17700, signal_17692}), .b ({signal_11267, signal_4189}), .c ({signal_11557, signal_4221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3572 ( .a ({signal_17716, signal_17708}), .b ({signal_11002, signal_4157}), .c ({signal_11267, signal_4189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3573 ( .a ({signal_17732, signal_17724}), .b ({signal_10770, signal_4125}), .c ({signal_11002, signal_4157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3574 ( .a ({signal_17748, signal_17740}), .b ({signal_11003, signal_4190}), .c ({signal_11268, signal_4222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3575 ( .a ({signal_17764, signal_17756}), .b ({signal_10765, signal_4158}), .c ({signal_11003, signal_4190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3576 ( .a ({signal_17780, signal_17772}), .b ({signal_10487, signal_4126}), .c ({signal_10765, signal_4158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3577 ( .a ({signal_17796, signal_17788}), .b ({signal_11004, signal_4191}), .c ({signal_11269, signal_4223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3578 ( .a ({signal_17812, signal_17804}), .b ({signal_10766, signal_4159}), .c ({signal_11004, signal_4191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3579 ( .a ({signal_17828, signal_17820}), .b ({signal_10488, signal_4127}), .c ({signal_10766, signal_4159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3580 ( .a ({signal_17844, signal_17836}), .b ({signal_11005, signal_4192}), .c ({signal_11270, signal_4224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3581 ( .a ({signal_17860, signal_17852}), .b ({signal_10767, signal_4160}), .c ({signal_11005, signal_4192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3582 ( .a ({signal_17876, signal_17868}), .b ({signal_10489, signal_4128}), .c ({signal_10767, signal_4160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3583 ( .a ({signal_17892, signal_17884}), .b ({signal_11271, signal_4193}), .c ({signal_11558, signal_4225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3584 ( .a ({signal_17908, signal_17900}), .b ({signal_11006, signal_4161}), .c ({signal_11271, signal_4193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3585 ( .a ({signal_17924, signal_17916}), .b ({signal_10771, signal_4129}), .c ({signal_11006, signal_4161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3586 ( .a ({signal_17940, signal_17932}), .b ({signal_11007, signal_4194}), .c ({signal_11272, signal_4226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3587 ( .a ({signal_17956, signal_17948}), .b ({signal_10768, signal_4162}), .c ({signal_11007, signal_4194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3588 ( .a ({signal_17972, signal_17964}), .b ({signal_10490, signal_4130}), .c ({signal_10768, signal_4162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3629 ( .a ({signal_17988, signal_17980}), .b ({signal_10293, signal_4517}), .c ({signal_10486, signal_4123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3630 ( .a ({signal_18004, signal_17996}), .b ({signal_10491, signal_4518}), .c ({signal_10769, signal_4124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3631 ( .a ({signal_18020, signal_18012}), .b ({signal_10492, signal_4519}), .c ({signal_10770, signal_4125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3632 ( .a ({signal_18036, signal_18028}), .b ({signal_10294, signal_4520}), .c ({signal_10487, signal_4126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3633 ( .a ({signal_18052, signal_18044}), .b ({signal_10295, signal_4521}), .c ({signal_10488, signal_4127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3634 ( .a ({signal_18068, signal_18060}), .b ({signal_10296, signal_4522}), .c ({signal_10489, signal_4128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3635 ( .a ({signal_18084, signal_18076}), .b ({signal_10493, signal_4523}), .c ({signal_10771, signal_4129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3636 ( .a ({signal_18100, signal_18092}), .b ({signal_10297, signal_4524}), .c ({signal_10490, signal_4130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3667 ( .a ({signal_10265, signal_3116}), .b ({1'b0, signal_18108}), .c ({signal_10293, signal_4517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3668 ( .a ({signal_10338, signal_3115}), .b ({1'b0, signal_18116}), .c ({signal_10491, signal_4518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3669 ( .a ({signal_10339, signal_3114}), .b ({1'b0, signal_18124}), .c ({signal_10492, signal_4519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3670 ( .a ({signal_10268, signal_3113}), .b ({1'b0, signal_18132}), .c ({signal_10294, signal_4520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3671 ( .a ({signal_10269, signal_3112}), .b ({1'b0, signal_18140}), .c ({signal_10295, signal_4521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3672 ( .a ({signal_10270, signal_3111}), .b ({1'b0, signal_18148}), .c ({signal_10296, signal_4522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3673 ( .a ({signal_10340, signal_3110}), .b ({1'b0, signal_18156}), .c ({signal_10493, signal_4523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3674 ( .a ({signal_10118, signal_3109}), .b ({1'b0, signal_18164}), .c ({signal_10297, signal_4524}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5601 ( .a ({signal_18176, signal_18170}), .b ({signal_9120, signal_5806}), .clk (clk), .r (Fresh[320]), .c ({signal_9229, signal_5837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5602 ( .a ({signal_18188, signal_18182}), .b ({signal_9119, signal_5805}), .clk (clk), .r (Fresh[321]), .c ({signal_9230, signal_5838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5603 ( .a ({signal_18200, signal_18194}), .b ({signal_9118, signal_5804}), .clk (clk), .r (Fresh[322]), .c ({signal_9231, signal_5839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5604 ( .a ({signal_18212, signal_18206}), .b ({signal_9117, signal_5803}), .clk (clk), .r (Fresh[323]), .c ({signal_9232, signal_5840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5605 ( .a ({signal_18224, signal_18218}), .b ({signal_9120, signal_5806}), .clk (clk), .r (Fresh[324]), .c ({signal_9233, signal_5841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5606 ( .a ({signal_18236, signal_18230}), .b ({signal_9119, signal_5805}), .clk (clk), .r (Fresh[325]), .c ({signal_9234, signal_5842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5607 ( .a ({signal_18248, signal_18242}), .b ({signal_9118, signal_5804}), .clk (clk), .r (Fresh[326]), .c ({signal_9235, signal_5843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5608 ( .a ({signal_18260, signal_18254}), .b ({signal_9117, signal_5803}), .clk (clk), .r (Fresh[327]), .c ({signal_9236, signal_5844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5609 ( .a ({signal_18272, signal_18266}), .b ({signal_9124, signal_5813}), .clk (clk), .r (Fresh[328]), .c ({signal_9237, signal_5845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5610 ( .a ({signal_18284, signal_18278}), .b ({signal_9123, signal_5812}), .clk (clk), .r (Fresh[329]), .c ({signal_9238, signal_5846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5611 ( .a ({signal_18296, signal_18290}), .b ({signal_9122, signal_5811}), .clk (clk), .r (Fresh[330]), .c ({signal_9239, signal_5847}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5612 ( .a ({signal_18308, signal_18302}), .b ({signal_9121, signal_5810}), .clk (clk), .r (Fresh[331]), .c ({signal_9240, signal_5848}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5613 ( .a ({signal_18320, signal_18314}), .b ({signal_9124, signal_5813}), .clk (clk), .r (Fresh[332]), .c ({signal_9241, signal_5849}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5614 ( .a ({signal_18332, signal_18326}), .b ({signal_9123, signal_5812}), .clk (clk), .r (Fresh[333]), .c ({signal_9242, signal_5850}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5615 ( .a ({signal_18344, signal_18338}), .b ({signal_9122, signal_5811}), .clk (clk), .r (Fresh[334]), .c ({signal_9243, signal_5851}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5616 ( .a ({signal_18356, signal_18350}), .b ({signal_9121, signal_5810}), .clk (clk), .r (Fresh[335]), .c ({signal_9244, signal_5852}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5617 ( .a ({signal_18368, signal_18362}), .b ({signal_9128, signal_5820}), .clk (clk), .r (Fresh[336]), .c ({signal_9245, signal_5853}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5618 ( .a ({signal_18380, signal_18374}), .b ({signal_9127, signal_5819}), .clk (clk), .r (Fresh[337]), .c ({signal_9246, signal_5854}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5619 ( .a ({signal_18392, signal_18386}), .b ({signal_9126, signal_5818}), .clk (clk), .r (Fresh[338]), .c ({signal_9247, signal_5855}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5620 ( .a ({signal_18404, signal_18398}), .b ({signal_9125, signal_5817}), .clk (clk), .r (Fresh[339]), .c ({signal_9248, signal_5856}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5621 ( .a ({signal_18416, signal_18410}), .b ({signal_9128, signal_5820}), .clk (clk), .r (Fresh[340]), .c ({signal_9249, signal_5857}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5622 ( .a ({signal_18428, signal_18422}), .b ({signal_9127, signal_5819}), .clk (clk), .r (Fresh[341]), .c ({signal_9250, signal_5858}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5623 ( .a ({signal_18440, signal_18434}), .b ({signal_9126, signal_5818}), .clk (clk), .r (Fresh[342]), .c ({signal_9251, signal_5859}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5624 ( .a ({signal_18452, signal_18446}), .b ({signal_9125, signal_5817}), .clk (clk), .r (Fresh[343]), .c ({signal_9252, signal_5860}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5625 ( .a ({signal_18464, signal_18458}), .b ({signal_9104, signal_5824}), .clk (clk), .r (Fresh[344]), .c ({signal_9129, signal_5861}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5626 ( .a ({signal_18476, signal_18470}), .b ({signal_9103, signal_5823}), .clk (clk), .r (Fresh[345]), .c ({signal_9130, signal_5862}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5627 ( .a ({signal_18488, signal_18482}), .b ({signal_9102, signal_5822}), .clk (clk), .r (Fresh[346]), .c ({signal_9131, signal_5863}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5628 ( .a ({signal_18500, signal_18494}), .b ({signal_9101, signal_5821}), .clk (clk), .r (Fresh[347]), .c ({signal_9132, signal_5864}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5629 ( .a ({signal_18512, signal_18506}), .b ({signal_9104, signal_5824}), .clk (clk), .r (Fresh[348]), .c ({signal_9133, signal_5865}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5630 ( .a ({signal_18524, signal_18518}), .b ({signal_9103, signal_5823}), .clk (clk), .r (Fresh[349]), .c ({signal_9134, signal_5866}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5631 ( .a ({signal_18536, signal_18530}), .b ({signal_9102, signal_5822}), .clk (clk), .r (Fresh[350]), .c ({signal_9135, signal_5867}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5632 ( .a ({signal_18548, signal_18542}), .b ({signal_9101, signal_5821}), .clk (clk), .r (Fresh[351]), .c ({signal_9136, signal_5868}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5633 ( .a ({signal_18560, signal_18554}), .b ({signal_9108, signal_5828}), .clk (clk), .r (Fresh[352]), .c ({signal_9137, signal_5869}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5634 ( .a ({signal_18572, signal_18566}), .b ({signal_9107, signal_5827}), .clk (clk), .r (Fresh[353]), .c ({signal_9138, signal_5870}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5635 ( .a ({signal_18584, signal_18578}), .b ({signal_9106, signal_5826}), .clk (clk), .r (Fresh[354]), .c ({signal_9139, signal_5871}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5636 ( .a ({signal_18596, signal_18590}), .b ({signal_9105, signal_5825}), .clk (clk), .r (Fresh[355]), .c ({signal_9140, signal_5872}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5637 ( .a ({signal_18608, signal_18602}), .b ({signal_9108, signal_5828}), .clk (clk), .r (Fresh[356]), .c ({signal_9141, signal_5873}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5638 ( .a ({signal_18620, signal_18614}), .b ({signal_9107, signal_5827}), .clk (clk), .r (Fresh[357]), .c ({signal_9142, signal_5874}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5639 ( .a ({signal_18632, signal_18626}), .b ({signal_9106, signal_5826}), .clk (clk), .r (Fresh[358]), .c ({signal_9143, signal_5875}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5640 ( .a ({signal_18644, signal_18638}), .b ({signal_9105, signal_5825}), .clk (clk), .r (Fresh[359]), .c ({signal_9144, signal_5876}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5641 ( .a ({signal_18656, signal_18650}), .b ({signal_9112, signal_5832}), .clk (clk), .r (Fresh[360]), .c ({signal_9145, signal_5877}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5642 ( .a ({signal_18668, signal_18662}), .b ({signal_9111, signal_5831}), .clk (clk), .r (Fresh[361]), .c ({signal_9146, signal_5878}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5643 ( .a ({signal_18680, signal_18674}), .b ({signal_9110, signal_5830}), .clk (clk), .r (Fresh[362]), .c ({signal_9147, signal_5879}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5644 ( .a ({signal_18692, signal_18686}), .b ({signal_9109, signal_5829}), .clk (clk), .r (Fresh[363]), .c ({signal_9148, signal_5880}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5645 ( .a ({signal_18704, signal_18698}), .b ({signal_9112, signal_5832}), .clk (clk), .r (Fresh[364]), .c ({signal_9149, signal_5881}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5646 ( .a ({signal_18716, signal_18710}), .b ({signal_9111, signal_5831}), .clk (clk), .r (Fresh[365]), .c ({signal_9150, signal_5882}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5647 ( .a ({signal_18728, signal_18722}), .b ({signal_9110, signal_5830}), .clk (clk), .r (Fresh[366]), .c ({signal_9151, signal_5883}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5648 ( .a ({signal_18740, signal_18734}), .b ({signal_9109, signal_5829}), .clk (clk), .r (Fresh[367]), .c ({signal_9152, signal_5884}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5649 ( .a ({signal_18752, signal_18746}), .b ({signal_9116, signal_5836}), .clk (clk), .r (Fresh[368]), .c ({signal_9153, signal_5885}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5650 ( .a ({signal_17938, signal_17930}), .b ({signal_9115, signal_5835}), .clk (clk), .r (Fresh[369]), .c ({signal_9154, signal_5886}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5651 ( .a ({signal_18764, signal_18758}), .b ({signal_9114, signal_5834}), .clk (clk), .r (Fresh[370]), .c ({signal_9155, signal_5887}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5652 ( .a ({signal_18776, signal_18770}), .b ({signal_9113, signal_5833}), .clk (clk), .r (Fresh[371]), .c ({signal_9156, signal_5888}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5653 ( .a ({signal_18788, signal_18782}), .b ({signal_9116, signal_5836}), .clk (clk), .r (Fresh[372]), .c ({signal_9157, signal_5889}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5654 ( .a ({signal_18800, signal_18794}), .b ({signal_9115, signal_5835}), .clk (clk), .r (Fresh[373]), .c ({signal_9158, signal_5890}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5655 ( .a ({signal_18812, signal_18806}), .b ({signal_9114, signal_5834}), .clk (clk), .r (Fresh[374]), .c ({signal_9159, signal_5891}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5656 ( .a ({signal_18824, signal_18818}), .b ({signal_9113, signal_5833}), .clk (clk), .r (Fresh[375]), .c ({signal_9160, signal_5892}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5737 ( .a ({signal_18836, signal_18830}), .b ({signal_9164, signal_5896}), .clk (clk), .r (Fresh[376]), .c ({signal_9265, signal_5973}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5738 ( .a ({signal_18848, signal_18842}), .b ({signal_9163, signal_5895}), .clk (clk), .r (Fresh[377]), .c ({signal_9266, signal_5974}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5739 ( .a ({signal_18860, signal_18854}), .b ({signal_9162, signal_5894}), .clk (clk), .r (Fresh[378]), .c ({signal_9267, signal_5975}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5740 ( .a ({signal_18872, signal_18866}), .b ({signal_9161, signal_5893}), .clk (clk), .r (Fresh[379]), .c ({signal_9268, signal_5976}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5741 ( .a ({signal_18884, signal_18878}), .b ({signal_9164, signal_5896}), .clk (clk), .r (Fresh[380]), .c ({signal_9269, signal_5977}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5742 ( .a ({signal_18896, signal_18890}), .b ({signal_9163, signal_5895}), .clk (clk), .r (Fresh[381]), .c ({signal_9270, signal_5978}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5743 ( .a ({signal_18908, signal_18902}), .b ({signal_9162, signal_5894}), .clk (clk), .r (Fresh[382]), .c ({signal_9271, signal_5979}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5744 ( .a ({signal_18920, signal_18914}), .b ({signal_9161, signal_5893}), .clk (clk), .r (Fresh[383]), .c ({signal_9272, signal_5980}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5745 ( .a ({signal_18932, signal_18926}), .b ({signal_9168, signal_5900}), .clk (clk), .r (Fresh[384]), .c ({signal_9273, signal_5981}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5746 ( .a ({signal_18944, signal_18938}), .b ({signal_9167, signal_5899}), .clk (clk), .r (Fresh[385]), .c ({signal_9274, signal_5982}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5747 ( .a ({signal_18956, signal_18950}), .b ({signal_9166, signal_5898}), .clk (clk), .r (Fresh[386]), .c ({signal_9275, signal_5983}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5748 ( .a ({signal_18968, signal_18962}), .b ({signal_9165, signal_5897}), .clk (clk), .r (Fresh[387]), .c ({signal_9276, signal_5984}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5749 ( .a ({signal_18980, signal_18974}), .b ({signal_9168, signal_5900}), .clk (clk), .r (Fresh[388]), .c ({signal_9277, signal_5985}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5750 ( .a ({signal_18992, signal_18986}), .b ({signal_9167, signal_5899}), .clk (clk), .r (Fresh[389]), .c ({signal_9278, signal_5986}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5751 ( .a ({signal_19004, signal_18998}), .b ({signal_9166, signal_5898}), .clk (clk), .r (Fresh[390]), .c ({signal_9279, signal_5987}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5752 ( .a ({signal_19016, signal_19010}), .b ({signal_9165, signal_5897}), .clk (clk), .r (Fresh[391]), .c ({signal_9280, signal_5988}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5753 ( .a ({signal_19028, signal_19022}), .b ({signal_9172, signal_5904}), .clk (clk), .r (Fresh[392]), .c ({signal_9281, signal_5989}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5754 ( .a ({signal_19040, signal_19034}), .b ({signal_9171, signal_5903}), .clk (clk), .r (Fresh[393]), .c ({signal_9282, signal_5990}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5755 ( .a ({signal_19052, signal_19046}), .b ({signal_9170, signal_5902}), .clk (clk), .r (Fresh[394]), .c ({signal_9283, signal_5991}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5756 ( .a ({signal_19064, signal_19058}), .b ({signal_9169, signal_5901}), .clk (clk), .r (Fresh[395]), .c ({signal_9284, signal_5992}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5757 ( .a ({signal_19076, signal_19070}), .b ({signal_9172, signal_5904}), .clk (clk), .r (Fresh[396]), .c ({signal_9285, signal_5993}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5758 ( .a ({signal_19088, signal_19082}), .b ({signal_9171, signal_5903}), .clk (clk), .r (Fresh[397]), .c ({signal_9286, signal_5994}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5759 ( .a ({signal_19100, signal_19094}), .b ({signal_9170, signal_5902}), .clk (clk), .r (Fresh[398]), .c ({signal_9287, signal_5995}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5760 ( .a ({signal_19112, signal_19106}), .b ({signal_9169, signal_5901}), .clk (clk), .r (Fresh[399]), .c ({signal_9288, signal_5996}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5761 ( .a ({signal_19124, signal_19118}), .b ({signal_9176, signal_5908}), .clk (clk), .r (Fresh[400]), .c ({signal_9289, signal_5997}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5762 ( .a ({signal_19136, signal_19130}), .b ({signal_9175, signal_5907}), .clk (clk), .r (Fresh[401]), .c ({signal_9290, signal_5998}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5763 ( .a ({signal_19148, signal_19142}), .b ({signal_9174, signal_5906}), .clk (clk), .r (Fresh[402]), .c ({signal_9291, signal_5999}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5764 ( .a ({signal_19160, signal_19154}), .b ({signal_9173, signal_5905}), .clk (clk), .r (Fresh[403]), .c ({signal_9292, signal_6000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5765 ( .a ({signal_19172, signal_19166}), .b ({signal_9176, signal_5908}), .clk (clk), .r (Fresh[404]), .c ({signal_9293, signal_6001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5766 ( .a ({signal_19184, signal_19178}), .b ({signal_9175, signal_5907}), .clk (clk), .r (Fresh[405]), .c ({signal_9294, signal_6002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5767 ( .a ({signal_19196, signal_19190}), .b ({signal_9174, signal_5906}), .clk (clk), .r (Fresh[406]), .c ({signal_9295, signal_6003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5768 ( .a ({signal_19208, signal_19202}), .b ({signal_9173, signal_5905}), .clk (clk), .r (Fresh[407]), .c ({signal_9296, signal_6004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5769 ( .a ({signal_19220, signal_19214}), .b ({signal_9180, signal_5912}), .clk (clk), .r (Fresh[408]), .c ({signal_9297, signal_6005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5770 ( .a ({signal_19232, signal_19226}), .b ({signal_9179, signal_5911}), .clk (clk), .r (Fresh[409]), .c ({signal_9298, signal_6006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5771 ( .a ({signal_19244, signal_19238}), .b ({signal_9178, signal_5910}), .clk (clk), .r (Fresh[410]), .c ({signal_9299, signal_6007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5772 ( .a ({signal_19256, signal_19250}), .b ({signal_9177, signal_5909}), .clk (clk), .r (Fresh[411]), .c ({signal_9300, signal_6008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5773 ( .a ({signal_19268, signal_19262}), .b ({signal_9180, signal_5912}), .clk (clk), .r (Fresh[412]), .c ({signal_9301, signal_6009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5774 ( .a ({signal_19280, signal_19274}), .b ({signal_9179, signal_5911}), .clk (clk), .r (Fresh[413]), .c ({signal_9302, signal_6010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5775 ( .a ({signal_19292, signal_19286}), .b ({signal_9178, signal_5910}), .clk (clk), .r (Fresh[414]), .c ({signal_9303, signal_6011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5776 ( .a ({signal_19304, signal_19298}), .b ({signal_9177, signal_5909}), .clk (clk), .r (Fresh[415]), .c ({signal_9304, signal_6012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5777 ( .a ({signal_19316, signal_19310}), .b ({signal_9184, signal_5916}), .clk (clk), .r (Fresh[416]), .c ({signal_9305, signal_6013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5778 ( .a ({signal_19328, signal_19322}), .b ({signal_9183, signal_5915}), .clk (clk), .r (Fresh[417]), .c ({signal_9306, signal_6014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5779 ( .a ({signal_19340, signal_19334}), .b ({signal_9182, signal_5914}), .clk (clk), .r (Fresh[418]), .c ({signal_9307, signal_6015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5780 ( .a ({signal_19352, signal_19346}), .b ({signal_9181, signal_5913}), .clk (clk), .r (Fresh[419]), .c ({signal_9308, signal_6016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5781 ( .a ({signal_19364, signal_19358}), .b ({signal_9184, signal_5916}), .clk (clk), .r (Fresh[420]), .c ({signal_9309, signal_6017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5782 ( .a ({signal_19376, signal_19370}), .b ({signal_9183, signal_5915}), .clk (clk), .r (Fresh[421]), .c ({signal_9310, signal_6018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5783 ( .a ({signal_19388, signal_19382}), .b ({signal_9182, signal_5914}), .clk (clk), .r (Fresh[422]), .c ({signal_9311, signal_6019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5784 ( .a ({signal_19400, signal_19394}), .b ({signal_9181, signal_5913}), .clk (clk), .r (Fresh[423]), .c ({signal_9312, signal_6020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5785 ( .a ({signal_19412, signal_19406}), .b ({signal_9188, signal_5920}), .clk (clk), .r (Fresh[424]), .c ({signal_9313, signal_6021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5786 ( .a ({signal_19424, signal_19418}), .b ({signal_9187, signal_5919}), .clk (clk), .r (Fresh[425]), .c ({signal_9314, signal_6022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5787 ( .a ({signal_19436, signal_19430}), .b ({signal_9186, signal_5918}), .clk (clk), .r (Fresh[426]), .c ({signal_9315, signal_6023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5788 ( .a ({signal_19448, signal_19442}), .b ({signal_9185, signal_5917}), .clk (clk), .r (Fresh[427]), .c ({signal_9316, signal_6024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5789 ( .a ({signal_19460, signal_19454}), .b ({signal_9188, signal_5920}), .clk (clk), .r (Fresh[428]), .c ({signal_9317, signal_6025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5790 ( .a ({signal_19472, signal_19466}), .b ({signal_9187, signal_5919}), .clk (clk), .r (Fresh[429]), .c ({signal_9318, signal_6026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5791 ( .a ({signal_19484, signal_19478}), .b ({signal_9186, signal_5918}), .clk (clk), .r (Fresh[430]), .c ({signal_9319, signal_6027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5792 ( .a ({signal_19496, signal_19490}), .b ({signal_9185, signal_5917}), .clk (clk), .r (Fresh[431]), .c ({signal_9320, signal_6028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5793 ( .a ({signal_19508, signal_19502}), .b ({signal_9256, signal_5924}), .clk (clk), .r (Fresh[432]), .c ({signal_9469, signal_6029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5794 ( .a ({signal_19520, signal_19514}), .b ({signal_9255, signal_5923}), .clk (clk), .r (Fresh[433]), .c ({signal_9470, signal_6030}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5795 ( .a ({signal_19532, signal_19526}), .b ({signal_9254, signal_5922}), .clk (clk), .r (Fresh[434]), .c ({signal_9471, signal_6031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5796 ( .a ({signal_19544, signal_19538}), .b ({signal_9253, signal_5921}), .clk (clk), .r (Fresh[435]), .c ({signal_9472, signal_6032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5797 ( .a ({signal_19556, signal_19550}), .b ({signal_9256, signal_5924}), .clk (clk), .r (Fresh[436]), .c ({signal_9473, signal_6033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5798 ( .a ({signal_19568, signal_19562}), .b ({signal_9255, signal_5923}), .clk (clk), .r (Fresh[437]), .c ({signal_9474, signal_6034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5799 ( .a ({signal_19580, signal_19574}), .b ({signal_9254, signal_5922}), .clk (clk), .r (Fresh[438]), .c ({signal_9475, signal_6035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5800 ( .a ({signal_19592, signal_19586}), .b ({signal_9253, signal_5921}), .clk (clk), .r (Fresh[439]), .c ({signal_9476, signal_6036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5801 ( .a ({signal_19604, signal_19598}), .b ({signal_9192, signal_5928}), .clk (clk), .r (Fresh[440]), .c ({signal_9321, signal_6037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5802 ( .a ({signal_19616, signal_19610}), .b ({signal_9191, signal_5927}), .clk (clk), .r (Fresh[441]), .c ({signal_9322, signal_6038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5803 ( .a ({signal_19628, signal_19622}), .b ({signal_9190, signal_5926}), .clk (clk), .r (Fresh[442]), .c ({signal_9323, signal_6039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5804 ( .a ({signal_19640, signal_19634}), .b ({signal_9189, signal_5925}), .clk (clk), .r (Fresh[443]), .c ({signal_9324, signal_6040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5805 ( .a ({signal_19652, signal_19646}), .b ({signal_9192, signal_5928}), .clk (clk), .r (Fresh[444]), .c ({signal_9325, signal_6041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5806 ( .a ({signal_19664, signal_19658}), .b ({signal_9191, signal_5927}), .clk (clk), .r (Fresh[445]), .c ({signal_9326, signal_6042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5807 ( .a ({signal_19676, signal_19670}), .b ({signal_9190, signal_5926}), .clk (clk), .r (Fresh[446]), .c ({signal_9327, signal_6043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5808 ( .a ({signal_19688, signal_19682}), .b ({signal_9189, signal_5925}), .clk (clk), .r (Fresh[447]), .c ({signal_9328, signal_6044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5809 ( .a ({signal_19700, signal_19694}), .b ({signal_9196, signal_5932}), .clk (clk), .r (Fresh[448]), .c ({signal_9329, signal_6045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5810 ( .a ({signal_19712, signal_19706}), .b ({signal_9195, signal_5931}), .clk (clk), .r (Fresh[449]), .c ({signal_9330, signal_6046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5811 ( .a ({signal_19724, signal_19718}), .b ({signal_9194, signal_5930}), .clk (clk), .r (Fresh[450]), .c ({signal_9331, signal_6047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5812 ( .a ({signal_19736, signal_19730}), .b ({signal_9193, signal_5929}), .clk (clk), .r (Fresh[451]), .c ({signal_9332, signal_6048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5813 ( .a ({signal_19748, signal_19742}), .b ({signal_9196, signal_5932}), .clk (clk), .r (Fresh[452]), .c ({signal_9333, signal_6049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5814 ( .a ({signal_19760, signal_19754}), .b ({signal_9195, signal_5931}), .clk (clk), .r (Fresh[453]), .c ({signal_9334, signal_6050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5815 ( .a ({signal_19772, signal_19766}), .b ({signal_9194, signal_5930}), .clk (clk), .r (Fresh[454]), .c ({signal_9335, signal_6051}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5816 ( .a ({signal_19784, signal_19778}), .b ({signal_9193, signal_5929}), .clk (clk), .r (Fresh[455]), .c ({signal_9336, signal_6052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5817 ( .a ({signal_19796, signal_19790}), .b ({signal_9200, signal_5936}), .clk (clk), .r (Fresh[456]), .c ({signal_9337, signal_6053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5818 ( .a ({signal_19808, signal_19802}), .b ({signal_9199, signal_5935}), .clk (clk), .r (Fresh[457]), .c ({signal_9338, signal_6054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5819 ( .a ({signal_19820, signal_19814}), .b ({signal_9198, signal_5934}), .clk (clk), .r (Fresh[458]), .c ({signal_9339, signal_6055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5820 ( .a ({signal_19832, signal_19826}), .b ({signal_9197, signal_5933}), .clk (clk), .r (Fresh[459]), .c ({signal_9340, signal_6056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5821 ( .a ({signal_19844, signal_19838}), .b ({signal_9200, signal_5936}), .clk (clk), .r (Fresh[460]), .c ({signal_9341, signal_6057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5822 ( .a ({signal_19856, signal_19850}), .b ({signal_9199, signal_5935}), .clk (clk), .r (Fresh[461]), .c ({signal_9342, signal_6058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5823 ( .a ({signal_19868, signal_19862}), .b ({signal_9198, signal_5934}), .clk (clk), .r (Fresh[462]), .c ({signal_9343, signal_6059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5824 ( .a ({signal_19880, signal_19874}), .b ({signal_9197, signal_5933}), .clk (clk), .r (Fresh[463]), .c ({signal_9344, signal_6060}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5825 ( .a ({signal_19892, signal_19886}), .b ({signal_9260, signal_5940}), .clk (clk), .r (Fresh[464]), .c ({signal_9477, signal_6061}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5826 ( .a ({signal_19904, signal_19898}), .b ({signal_9259, signal_5939}), .clk (clk), .r (Fresh[465]), .c ({signal_9478, signal_6062}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5827 ( .a ({signal_19916, signal_19910}), .b ({signal_9258, signal_5938}), .clk (clk), .r (Fresh[466]), .c ({signal_9479, signal_6063}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5828 ( .a ({signal_19928, signal_19922}), .b ({signal_9257, signal_5937}), .clk (clk), .r (Fresh[467]), .c ({signal_9480, signal_6064}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5829 ( .a ({signal_19940, signal_19934}), .b ({signal_9260, signal_5940}), .clk (clk), .r (Fresh[468]), .c ({signal_9481, signal_6065}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5830 ( .a ({signal_19952, signal_19946}), .b ({signal_9259, signal_5939}), .clk (clk), .r (Fresh[469]), .c ({signal_9482, signal_6066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5831 ( .a ({signal_19964, signal_19958}), .b ({signal_9258, signal_5938}), .clk (clk), .r (Fresh[470]), .c ({signal_9483, signal_6067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5832 ( .a ({signal_19976, signal_19970}), .b ({signal_9257, signal_5937}), .clk (clk), .r (Fresh[471]), .c ({signal_9484, signal_6068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5833 ( .a ({signal_19988, signal_19982}), .b ({signal_9204, signal_5944}), .clk (clk), .r (Fresh[472]), .c ({signal_9345, signal_6069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5834 ( .a ({signal_20000, signal_19994}), .b ({signal_9203, signal_5943}), .clk (clk), .r (Fresh[473]), .c ({signal_9346, signal_6070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5835 ( .a ({signal_20012, signal_20006}), .b ({signal_9202, signal_5942}), .clk (clk), .r (Fresh[474]), .c ({signal_9347, signal_6071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5836 ( .a ({signal_20024, signal_20018}), .b ({signal_9201, signal_5941}), .clk (clk), .r (Fresh[475]), .c ({signal_9348, signal_6072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5837 ( .a ({signal_20036, signal_20030}), .b ({signal_9204, signal_5944}), .clk (clk), .r (Fresh[476]), .c ({signal_9349, signal_6073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5838 ( .a ({signal_20048, signal_20042}), .b ({signal_9203, signal_5943}), .clk (clk), .r (Fresh[477]), .c ({signal_9350, signal_6074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5839 ( .a ({signal_20060, signal_20054}), .b ({signal_9202, signal_5942}), .clk (clk), .r (Fresh[478]), .c ({signal_9351, signal_6075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5840 ( .a ({signal_20072, signal_20066}), .b ({signal_9201, signal_5941}), .clk (clk), .r (Fresh[479]), .c ({signal_9352, signal_6076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5841 ( .a ({signal_20084, signal_20078}), .b ({signal_9208, signal_5948}), .clk (clk), .r (Fresh[480]), .c ({signal_9353, signal_6077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5842 ( .a ({signal_20096, signal_20090}), .b ({signal_9207, signal_5947}), .clk (clk), .r (Fresh[481]), .c ({signal_9354, signal_6078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5843 ( .a ({signal_20108, signal_20102}), .b ({signal_9206, signal_5946}), .clk (clk), .r (Fresh[482]), .c ({signal_9355, signal_6079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5844 ( .a ({signal_20120, signal_20114}), .b ({signal_9205, signal_5945}), .clk (clk), .r (Fresh[483]), .c ({signal_9356, signal_6080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5845 ( .a ({signal_20132, signal_20126}), .b ({signal_9208, signal_5948}), .clk (clk), .r (Fresh[484]), .c ({signal_9357, signal_6081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5846 ( .a ({signal_20144, signal_20138}), .b ({signal_9207, signal_5947}), .clk (clk), .r (Fresh[485]), .c ({signal_9358, signal_6082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5847 ( .a ({signal_20156, signal_20150}), .b ({signal_9206, signal_5946}), .clk (clk), .r (Fresh[486]), .c ({signal_9359, signal_6083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5848 ( .a ({signal_20168, signal_20162}), .b ({signal_9205, signal_5945}), .clk (clk), .r (Fresh[487]), .c ({signal_9360, signal_6084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5849 ( .a ({signal_20180, signal_20174}), .b ({signal_9212, signal_5952}), .clk (clk), .r (Fresh[488]), .c ({signal_9361, signal_6085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5850 ( .a ({signal_20192, signal_20186}), .b ({signal_9211, signal_5951}), .clk (clk), .r (Fresh[489]), .c ({signal_9362, signal_6086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5851 ( .a ({signal_20204, signal_20198}), .b ({signal_9210, signal_5950}), .clk (clk), .r (Fresh[490]), .c ({signal_9363, signal_6087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5852 ( .a ({signal_20216, signal_20210}), .b ({signal_9209, signal_5949}), .clk (clk), .r (Fresh[491]), .c ({signal_9364, signal_6088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5853 ( .a ({signal_20228, signal_20222}), .b ({signal_9212, signal_5952}), .clk (clk), .r (Fresh[492]), .c ({signal_9365, signal_6089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5854 ( .a ({signal_20240, signal_20234}), .b ({signal_9211, signal_5951}), .clk (clk), .r (Fresh[493]), .c ({signal_9366, signal_6090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5855 ( .a ({signal_20252, signal_20246}), .b ({signal_9210, signal_5950}), .clk (clk), .r (Fresh[494]), .c ({signal_9367, signal_6091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5856 ( .a ({signal_20264, signal_20258}), .b ({signal_9209, signal_5949}), .clk (clk), .r (Fresh[495]), .c ({signal_9368, signal_6092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5857 ( .a ({signal_20276, signal_20270}), .b ({signal_9264, signal_5956}), .clk (clk), .r (Fresh[496]), .c ({signal_9485, signal_6093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5858 ( .a ({signal_20288, signal_20282}), .b ({signal_9263, signal_5955}), .clk (clk), .r (Fresh[497]), .c ({signal_9486, signal_6094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5859 ( .a ({signal_20300, signal_20294}), .b ({signal_9262, signal_5954}), .clk (clk), .r (Fresh[498]), .c ({signal_9487, signal_6095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5860 ( .a ({signal_20312, signal_20306}), .b ({signal_9261, signal_5953}), .clk (clk), .r (Fresh[499]), .c ({signal_9488, signal_6096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5861 ( .a ({signal_20324, signal_20318}), .b ({signal_9264, signal_5956}), .clk (clk), .r (Fresh[500]), .c ({signal_9489, signal_6097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5862 ( .a ({signal_20336, signal_20330}), .b ({signal_9263, signal_5955}), .clk (clk), .r (Fresh[501]), .c ({signal_9490, signal_6098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5863 ( .a ({signal_20348, signal_20342}), .b ({signal_9262, signal_5954}), .clk (clk), .r (Fresh[502]), .c ({signal_9491, signal_6099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5864 ( .a ({signal_20360, signal_20354}), .b ({signal_9261, signal_5953}), .clk (clk), .r (Fresh[503]), .c ({signal_9492, signal_6100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5865 ( .a ({signal_20372, signal_20366}), .b ({signal_9216, signal_5960}), .clk (clk), .r (Fresh[504]), .c ({signal_9369, signal_6101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5866 ( .a ({signal_20384, signal_20378}), .b ({signal_9215, signal_5959}), .clk (clk), .r (Fresh[505]), .c ({signal_9370, signal_6102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5867 ( .a ({signal_20396, signal_20390}), .b ({signal_9214, signal_5958}), .clk (clk), .r (Fresh[506]), .c ({signal_9371, signal_6103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5868 ( .a ({signal_20408, signal_20402}), .b ({signal_9213, signal_5957}), .clk (clk), .r (Fresh[507]), .c ({signal_9372, signal_6104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5869 ( .a ({signal_20420, signal_20414}), .b ({signal_9216, signal_5960}), .clk (clk), .r (Fresh[508]), .c ({signal_9373, signal_6105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5870 ( .a ({signal_20432, signal_20426}), .b ({signal_9215, signal_5959}), .clk (clk), .r (Fresh[509]), .c ({signal_9374, signal_6106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5871 ( .a ({signal_20444, signal_20438}), .b ({signal_9214, signal_5958}), .clk (clk), .r (Fresh[510]), .c ({signal_9375, signal_6107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5872 ( .a ({signal_20456, signal_20450}), .b ({signal_9213, signal_5957}), .clk (clk), .r (Fresh[511]), .c ({signal_9376, signal_6108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5873 ( .a ({signal_20468, signal_20462}), .b ({signal_9220, signal_5964}), .clk (clk), .r (Fresh[512]), .c ({signal_9377, signal_6109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5874 ( .a ({signal_20480, signal_20474}), .b ({signal_9219, signal_5963}), .clk (clk), .r (Fresh[513]), .c ({signal_9378, signal_6110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5875 ( .a ({signal_20492, signal_20486}), .b ({signal_9218, signal_5962}), .clk (clk), .r (Fresh[514]), .c ({signal_9379, signal_6111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5876 ( .a ({signal_20504, signal_20498}), .b ({signal_9217, signal_5961}), .clk (clk), .r (Fresh[515]), .c ({signal_9380, signal_6112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5877 ( .a ({signal_20516, signal_20510}), .b ({signal_9220, signal_5964}), .clk (clk), .r (Fresh[516]), .c ({signal_9381, signal_6113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5878 ( .a ({signal_20528, signal_20522}), .b ({signal_9219, signal_5963}), .clk (clk), .r (Fresh[517]), .c ({signal_9382, signal_6114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5879 ( .a ({signal_20540, signal_20534}), .b ({signal_9218, signal_5962}), .clk (clk), .r (Fresh[518]), .c ({signal_9383, signal_6115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5880 ( .a ({signal_20552, signal_20546}), .b ({signal_9217, signal_5961}), .clk (clk), .r (Fresh[519]), .c ({signal_9384, signal_6116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5881 ( .a ({signal_20564, signal_20558}), .b ({signal_9224, signal_5968}), .clk (clk), .r (Fresh[520]), .c ({signal_9385, signal_6117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5882 ( .a ({signal_20576, signal_20570}), .b ({signal_9223, signal_5967}), .clk (clk), .r (Fresh[521]), .c ({signal_9386, signal_6118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5883 ( .a ({signal_20588, signal_20582}), .b ({signal_9222, signal_5966}), .clk (clk), .r (Fresh[522]), .c ({signal_9387, signal_6119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5884 ( .a ({signal_20600, signal_20594}), .b ({signal_9221, signal_5965}), .clk (clk), .r (Fresh[523]), .c ({signal_9388, signal_6120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5885 ( .a ({signal_20612, signal_20606}), .b ({signal_9224, signal_5968}), .clk (clk), .r (Fresh[524]), .c ({signal_9389, signal_6121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5886 ( .a ({signal_20624, signal_20618}), .b ({signal_9223, signal_5967}), .clk (clk), .r (Fresh[525]), .c ({signal_9390, signal_6122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5887 ( .a ({signal_20636, signal_20630}), .b ({signal_9222, signal_5966}), .clk (clk), .r (Fresh[526]), .c ({signal_9391, signal_6123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5888 ( .a ({signal_20648, signal_20642}), .b ({signal_9221, signal_5965}), .clk (clk), .r (Fresh[527]), .c ({signal_9392, signal_6124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5889 ( .a ({signal_20660, signal_20654}), .b ({signal_9228, signal_5972}), .clk (clk), .r (Fresh[528]), .c ({signal_9393, signal_6125}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5890 ( .a ({signal_20672, signal_20666}), .b ({signal_9227, signal_5971}), .clk (clk), .r (Fresh[529]), .c ({signal_9394, signal_6126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5891 ( .a ({signal_20684, signal_20678}), .b ({signal_9226, signal_5970}), .clk (clk), .r (Fresh[530]), .c ({signal_9395, signal_6127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5892 ( .a ({signal_20696, signal_20690}), .b ({signal_9225, signal_5969}), .clk (clk), .r (Fresh[531]), .c ({signal_9396, signal_6128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5893 ( .a ({signal_20708, signal_20702}), .b ({signal_9228, signal_5972}), .clk (clk), .r (Fresh[532]), .c ({signal_9397, signal_6129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5894 ( .a ({signal_20720, signal_20714}), .b ({signal_9227, signal_5971}), .clk (clk), .r (Fresh[533]), .c ({signal_9398, signal_6130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5895 ( .a ({signal_20732, signal_20726}), .b ({signal_9226, signal_5970}), .clk (clk), .r (Fresh[534]), .c ({signal_9399, signal_6131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5896 ( .a ({signal_20744, signal_20738}), .b ({signal_9225, signal_5969}), .clk (clk), .r (Fresh[535]), .c ({signal_9400, signal_6132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5926 ( .a ({signal_9231, signal_5839}), .b ({signal_9233, signal_5841}), .c ({signal_9494, signal_6162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5927 ( .a ({signal_9232, signal_5840}), .b ({signal_9235, signal_5843}), .c ({signal_9495, signal_6163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5928 ( .a ({signal_9230, signal_5838}), .b ({signal_9232, signal_5840}), .c ({signal_9496, signal_6164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5942 ( .a ({signal_9239, signal_5847}), .b ({signal_9241, signal_5849}), .c ({signal_9498, signal_6178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5943 ( .a ({signal_9240, signal_5848}), .b ({signal_9243, signal_5851}), .c ({signal_9499, signal_6179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5944 ( .a ({signal_9238, signal_5846}), .b ({signal_9240, signal_5848}), .c ({signal_9500, signal_6180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5958 ( .a ({signal_9247, signal_5855}), .b ({signal_9249, signal_5857}), .c ({signal_9502, signal_6194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5959 ( .a ({signal_9248, signal_5856}), .b ({signal_9251, signal_5859}), .c ({signal_9503, signal_6195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5960 ( .a ({signal_9246, signal_5854}), .b ({signal_9248, signal_5856}), .c ({signal_9504, signal_6196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5962 ( .a ({signal_9131, signal_5863}), .b ({signal_9133, signal_5865}), .c ({signal_9454, signal_6198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5963 ( .a ({signal_9132, signal_5864}), .b ({signal_9135, signal_5867}), .c ({signal_9455, signal_6199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5964 ( .a ({signal_9130, signal_5862}), .b ({signal_9132, signal_5864}), .c ({signal_9456, signal_6200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5966 ( .a ({signal_9139, signal_5871}), .b ({signal_9141, signal_5873}), .c ({signal_9458, signal_6202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5967 ( .a ({signal_9140, signal_5872}), .b ({signal_9143, signal_5875}), .c ({signal_9459, signal_6203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5968 ( .a ({signal_9138, signal_5870}), .b ({signal_9140, signal_5872}), .c ({signal_9460, signal_6204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5970 ( .a ({signal_9147, signal_5879}), .b ({signal_9149, signal_5881}), .c ({signal_9462, signal_6206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5971 ( .a ({signal_9148, signal_5880}), .b ({signal_9151, signal_5883}), .c ({signal_9463, signal_6207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5972 ( .a ({signal_9146, signal_5878}), .b ({signal_9148, signal_5880}), .c ({signal_9464, signal_6208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5974 ( .a ({signal_9155, signal_5887}), .b ({signal_9157, signal_5889}), .c ({signal_9466, signal_6210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5975 ( .a ({signal_9156, signal_5888}), .b ({signal_9159, signal_5891}), .c ({signal_9467, signal_6211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5976 ( .a ({signal_9154, signal_5886}), .b ({signal_9156, signal_5888}), .c ({signal_9468, signal_6212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5977 ( .a ({signal_20756, signal_20750}), .b ({signal_9404, signal_6136}), .clk (clk), .r (Fresh[536]), .c ({signal_9505, signal_6213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5978 ( .a ({signal_20768, signal_20762}), .b ({signal_9403, signal_6135}), .clk (clk), .r (Fresh[537]), .c ({signal_9506, signal_6214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5979 ( .a ({signal_20780, signal_20774}), .b ({signal_9402, signal_6134}), .clk (clk), .r (Fresh[538]), .c ({signal_9507, signal_6215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5980 ( .a ({signal_20792, signal_20786}), .b ({signal_9401, signal_6133}), .clk (clk), .r (Fresh[539]), .c ({signal_9508, signal_6216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5981 ( .a ({signal_20804, signal_20798}), .b ({signal_9404, signal_6136}), .clk (clk), .r (Fresh[540]), .c ({signal_9509, signal_6217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5982 ( .a ({signal_20816, signal_20810}), .b ({signal_9403, signal_6135}), .clk (clk), .r (Fresh[541]), .c ({signal_9510, signal_6218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5983 ( .a ({signal_20828, signal_20822}), .b ({signal_9402, signal_6134}), .clk (clk), .r (Fresh[542]), .c ({signal_9511, signal_6219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5984 ( .a ({signal_20840, signal_20834}), .b ({signal_9401, signal_6133}), .clk (clk), .r (Fresh[543]), .c ({signal_9512, signal_6220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5985 ( .a ({signal_20852, signal_20846}), .b ({signal_9408, signal_6140}), .clk (clk), .r (Fresh[544]), .c ({signal_9513, signal_6221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5986 ( .a ({signal_20864, signal_20858}), .b ({signal_9407, signal_6139}), .clk (clk), .r (Fresh[545]), .c ({signal_9514, signal_6222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5987 ( .a ({signal_20876, signal_20870}), .b ({signal_9406, signal_6138}), .clk (clk), .r (Fresh[546]), .c ({signal_9515, signal_6223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5988 ( .a ({signal_20888, signal_20882}), .b ({signal_9405, signal_6137}), .clk (clk), .r (Fresh[547]), .c ({signal_9516, signal_6224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5989 ( .a ({signal_20900, signal_20894}), .b ({signal_9408, signal_6140}), .clk (clk), .r (Fresh[548]), .c ({signal_9517, signal_6225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5990 ( .a ({signal_20912, signal_20906}), .b ({signal_9407, signal_6139}), .clk (clk), .r (Fresh[549]), .c ({signal_9518, signal_6226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5991 ( .a ({signal_20924, signal_20918}), .b ({signal_9406, signal_6138}), .clk (clk), .r (Fresh[550]), .c ({signal_9519, signal_6227}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5992 ( .a ({signal_20936, signal_20930}), .b ({signal_9405, signal_6137}), .clk (clk), .r (Fresh[551]), .c ({signal_9520, signal_6228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5993 ( .a ({signal_20948, signal_20942}), .b ({signal_9412, signal_6144}), .clk (clk), .r (Fresh[552]), .c ({signal_9521, signal_6229}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5994 ( .a ({signal_20960, signal_20954}), .b ({signal_9411, signal_6143}), .clk (clk), .r (Fresh[553]), .c ({signal_9522, signal_6230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5995 ( .a ({signal_20972, signal_20966}), .b ({signal_9410, signal_6142}), .clk (clk), .r (Fresh[554]), .c ({signal_9523, signal_6231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5996 ( .a ({signal_20984, signal_20978}), .b ({signal_9409, signal_6141}), .clk (clk), .r (Fresh[555]), .c ({signal_9524, signal_6232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5997 ( .a ({signal_20996, signal_20990}), .b ({signal_9412, signal_6144}), .clk (clk), .r (Fresh[556]), .c ({signal_9525, signal_6233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5998 ( .a ({signal_21008, signal_21002}), .b ({signal_9411, signal_6143}), .clk (clk), .r (Fresh[557]), .c ({signal_9526, signal_6234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_5999 ( .a ({signal_21020, signal_21014}), .b ({signal_9410, signal_6142}), .clk (clk), .r (Fresh[558]), .c ({signal_9527, signal_6235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6000 ( .a ({signal_21032, signal_21026}), .b ({signal_9409, signal_6141}), .clk (clk), .r (Fresh[559]), .c ({signal_9528, signal_6236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6001 ( .a ({signal_21044, signal_21038}), .b ({signal_9416, signal_6148}), .clk (clk), .r (Fresh[560]), .c ({signal_9529, signal_6237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6002 ( .a ({signal_21056, signal_21050}), .b ({signal_9415, signal_6147}), .clk (clk), .r (Fresh[561]), .c ({signal_9530, signal_6238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6003 ( .a ({signal_21068, signal_21062}), .b ({signal_9414, signal_6146}), .clk (clk), .r (Fresh[562]), .c ({signal_9531, signal_6239}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6004 ( .a ({signal_21080, signal_21074}), .b ({signal_9413, signal_6145}), .clk (clk), .r (Fresh[563]), .c ({signal_9532, signal_6240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6005 ( .a ({signal_21092, signal_21086}), .b ({signal_9416, signal_6148}), .clk (clk), .r (Fresh[564]), .c ({signal_9533, signal_6241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6006 ( .a ({signal_21104, signal_21098}), .b ({signal_9415, signal_6147}), .clk (clk), .r (Fresh[565]), .c ({signal_9534, signal_6242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6007 ( .a ({signal_21116, signal_21110}), .b ({signal_9414, signal_6146}), .clk (clk), .r (Fresh[566]), .c ({signal_9535, signal_6243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6008 ( .a ({signal_21128, signal_21122}), .b ({signal_9413, signal_6145}), .clk (clk), .r (Fresh[567]), .c ({signal_9536, signal_6244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6009 ( .a ({signal_21140, signal_21134}), .b ({signal_9420, signal_6152}), .clk (clk), .r (Fresh[568]), .c ({signal_9537, signal_6245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6010 ( .a ({signal_21152, signal_21146}), .b ({signal_9419, signal_6151}), .clk (clk), .r (Fresh[569]), .c ({signal_9538, signal_6246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6011 ( .a ({signal_21164, signal_21158}), .b ({signal_9418, signal_6150}), .clk (clk), .r (Fresh[570]), .c ({signal_9539, signal_6247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6012 ( .a ({signal_21176, signal_21170}), .b ({signal_9417, signal_6149}), .clk (clk), .r (Fresh[571]), .c ({signal_9540, signal_6248}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6013 ( .a ({signal_21188, signal_21182}), .b ({signal_9420, signal_6152}), .clk (clk), .r (Fresh[572]), .c ({signal_9541, signal_6249}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6014 ( .a ({signal_21200, signal_21194}), .b ({signal_9419, signal_6151}), .clk (clk), .r (Fresh[573]), .c ({signal_9542, signal_6250}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6015 ( .a ({signal_21212, signal_21206}), .b ({signal_9418, signal_6150}), .clk (clk), .r (Fresh[574]), .c ({signal_9543, signal_6251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6016 ( .a ({signal_21224, signal_21218}), .b ({signal_9417, signal_6149}), .clk (clk), .r (Fresh[575]), .c ({signal_9544, signal_6252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6017 ( .a ({signal_21236, signal_21230}), .b ({signal_9424, signal_6156}), .clk (clk), .r (Fresh[576]), .c ({signal_9545, signal_6253}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6018 ( .a ({signal_21248, signal_21242}), .b ({signal_9423, signal_6155}), .clk (clk), .r (Fresh[577]), .c ({signal_9546, signal_6254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6019 ( .a ({signal_21260, signal_21254}), .b ({signal_9422, signal_6154}), .clk (clk), .r (Fresh[578]), .c ({signal_9547, signal_6255}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6020 ( .a ({signal_21272, signal_21266}), .b ({signal_9421, signal_6153}), .clk (clk), .r (Fresh[579]), .c ({signal_9548, signal_6256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6021 ( .a ({signal_21284, signal_21278}), .b ({signal_9424, signal_6156}), .clk (clk), .r (Fresh[580]), .c ({signal_9549, signal_6257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6022 ( .a ({signal_21296, signal_21290}), .b ({signal_9423, signal_6155}), .clk (clk), .r (Fresh[581]), .c ({signal_9550, signal_6258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6023 ( .a ({signal_21308, signal_21302}), .b ({signal_9422, signal_6154}), .clk (clk), .r (Fresh[582]), .c ({signal_9551, signal_6259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6024 ( .a ({signal_21320, signal_21314}), .b ({signal_9421, signal_6153}), .clk (clk), .r (Fresh[583]), .c ({signal_9552, signal_6260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6025 ( .a ({signal_21332, signal_21326}), .b ({signal_9428, signal_6160}), .clk (clk), .r (Fresh[584]), .c ({signal_9553, signal_6261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6026 ( .a ({signal_21344, signal_21338}), .b ({signal_9427, signal_6159}), .clk (clk), .r (Fresh[585]), .c ({signal_9554, signal_6262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6027 ( .a ({signal_21356, signal_21350}), .b ({signal_9426, signal_6158}), .clk (clk), .r (Fresh[586]), .c ({signal_9555, signal_6263}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6028 ( .a ({signal_21368, signal_21362}), .b ({signal_9425, signal_6157}), .clk (clk), .r (Fresh[587]), .c ({signal_9556, signal_6264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6029 ( .a ({signal_21380, signal_21374}), .b ({signal_9428, signal_6160}), .clk (clk), .r (Fresh[588]), .c ({signal_9557, signal_6265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6030 ( .a ({signal_21392, signal_21386}), .b ({signal_9427, signal_6159}), .clk (clk), .r (Fresh[589]), .c ({signal_9558, signal_6266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6031 ( .a ({signal_21404, signal_21398}), .b ({signal_9426, signal_6158}), .clk (clk), .r (Fresh[590]), .c ({signal_9559, signal_6267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6032 ( .a ({signal_21416, signal_21410}), .b ({signal_9425, signal_6157}), .clk (clk), .r (Fresh[591]), .c ({signal_9560, signal_6268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6033 ( .a ({signal_21428, signal_21422}), .b ({signal_9493, signal_6161}), .clk (clk), .r (Fresh[592]), .c ({signal_9701, signal_6269}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6034 ( .a ({signal_21440, signal_21434}), .b ({signal_9493, signal_6161}), .clk (clk), .r (Fresh[593]), .c ({signal_9702, signal_6270}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6035 ( .a ({signal_21452, signal_21446}), .b ({signal_9432, signal_6168}), .clk (clk), .r (Fresh[594]), .c ({signal_9561, signal_6271}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6036 ( .a ({signal_21464, signal_21458}), .b ({signal_9431, signal_6167}), .clk (clk), .r (Fresh[595]), .c ({signal_9562, signal_6272}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6037 ( .a ({signal_21476, signal_21470}), .b ({signal_9430, signal_6166}), .clk (clk), .r (Fresh[596]), .c ({signal_9563, signal_6273}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6038 ( .a ({signal_21488, signal_21482}), .b ({signal_9429, signal_6165}), .clk (clk), .r (Fresh[597]), .c ({signal_9564, signal_6274}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6039 ( .a ({signal_21500, signal_21494}), .b ({signal_9432, signal_6168}), .clk (clk), .r (Fresh[598]), .c ({signal_9565, signal_6275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6040 ( .a ({signal_21512, signal_21506}), .b ({signal_9431, signal_6167}), .clk (clk), .r (Fresh[599]), .c ({signal_9566, signal_6276}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6041 ( .a ({signal_21524, signal_21518}), .b ({signal_9430, signal_6166}), .clk (clk), .r (Fresh[600]), .c ({signal_9567, signal_6277}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6042 ( .a ({signal_21536, signal_21530}), .b ({signal_9429, signal_6165}), .clk (clk), .r (Fresh[601]), .c ({signal_9568, signal_6278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6043 ( .a ({signal_21548, signal_21542}), .b ({signal_9436, signal_6172}), .clk (clk), .r (Fresh[602]), .c ({signal_9569, signal_6279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6044 ( .a ({signal_21560, signal_21554}), .b ({signal_9435, signal_6171}), .clk (clk), .r (Fresh[603]), .c ({signal_9570, signal_6280}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6045 ( .a ({signal_21572, signal_21566}), .b ({signal_9434, signal_6170}), .clk (clk), .r (Fresh[604]), .c ({signal_9571, signal_6281}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6046 ( .a ({signal_21584, signal_21578}), .b ({signal_9433, signal_6169}), .clk (clk), .r (Fresh[605]), .c ({signal_9572, signal_6282}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6047 ( .a ({signal_21596, signal_21590}), .b ({signal_9436, signal_6172}), .clk (clk), .r (Fresh[606]), .c ({signal_9573, signal_6283}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6048 ( .a ({signal_21608, signal_21602}), .b ({signal_9435, signal_6171}), .clk (clk), .r (Fresh[607]), .c ({signal_9574, signal_6284}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6049 ( .a ({signal_21620, signal_21614}), .b ({signal_9434, signal_6170}), .clk (clk), .r (Fresh[608]), .c ({signal_9575, signal_6285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6050 ( .a ({signal_21632, signal_21626}), .b ({signal_9433, signal_6169}), .clk (clk), .r (Fresh[609]), .c ({signal_9576, signal_6286}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6051 ( .a ({signal_21644, signal_21638}), .b ({signal_9440, signal_6176}), .clk (clk), .r (Fresh[610]), .c ({signal_9577, signal_6287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6052 ( .a ({signal_21656, signal_21650}), .b ({signal_9439, signal_6175}), .clk (clk), .r (Fresh[611]), .c ({signal_9578, signal_6288}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6053 ( .a ({signal_21668, signal_21662}), .b ({signal_9438, signal_6174}), .clk (clk), .r (Fresh[612]), .c ({signal_9579, signal_6289}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6054 ( .a ({signal_21680, signal_21674}), .b ({signal_9437, signal_6173}), .clk (clk), .r (Fresh[613]), .c ({signal_9580, signal_6290}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6055 ( .a ({signal_21692, signal_21686}), .b ({signal_9440, signal_6176}), .clk (clk), .r (Fresh[614]), .c ({signal_9581, signal_6291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6056 ( .a ({signal_21704, signal_21698}), .b ({signal_9439, signal_6175}), .clk (clk), .r (Fresh[615]), .c ({signal_9582, signal_6292}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6057 ( .a ({signal_21716, signal_21710}), .b ({signal_9438, signal_6174}), .clk (clk), .r (Fresh[616]), .c ({signal_9583, signal_6293}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6058 ( .a ({signal_21728, signal_21722}), .b ({signal_9437, signal_6173}), .clk (clk), .r (Fresh[617]), .c ({signal_9584, signal_6294}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6059 ( .a ({signal_21740, signal_21734}), .b ({signal_9497, signal_6177}), .clk (clk), .r (Fresh[618]), .c ({signal_9703, signal_6295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6060 ( .a ({signal_21752, signal_21746}), .b ({signal_9497, signal_6177}), .clk (clk), .r (Fresh[619]), .c ({signal_9704, signal_6296}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6061 ( .a ({signal_21764, signal_21758}), .b ({signal_9444, signal_6184}), .clk (clk), .r (Fresh[620]), .c ({signal_9585, signal_6297}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6062 ( .a ({signal_21776, signal_21770}), .b ({signal_9443, signal_6183}), .clk (clk), .r (Fresh[621]), .c ({signal_9586, signal_6298}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6063 ( .a ({signal_21788, signal_21782}), .b ({signal_9442, signal_6182}), .clk (clk), .r (Fresh[622]), .c ({signal_9587, signal_6299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6064 ( .a ({signal_21800, signal_21794}), .b ({signal_9441, signal_6181}), .clk (clk), .r (Fresh[623]), .c ({signal_9588, signal_6300}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6065 ( .a ({signal_21812, signal_21806}), .b ({signal_9444, signal_6184}), .clk (clk), .r (Fresh[624]), .c ({signal_9589, signal_6301}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6066 ( .a ({signal_21824, signal_21818}), .b ({signal_9443, signal_6183}), .clk (clk), .r (Fresh[625]), .c ({signal_9590, signal_6302}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6067 ( .a ({signal_21836, signal_21830}), .b ({signal_9442, signal_6182}), .clk (clk), .r (Fresh[626]), .c ({signal_9591, signal_6303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6068 ( .a ({signal_21848, signal_21842}), .b ({signal_9441, signal_6181}), .clk (clk), .r (Fresh[627]), .c ({signal_9592, signal_6304}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6069 ( .a ({signal_21860, signal_21854}), .b ({signal_9448, signal_6188}), .clk (clk), .r (Fresh[628]), .c ({signal_9593, signal_6305}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6070 ( .a ({signal_21872, signal_21866}), .b ({signal_9447, signal_6187}), .clk (clk), .r (Fresh[629]), .c ({signal_9594, signal_6306}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6071 ( .a ({signal_21884, signal_21878}), .b ({signal_9446, signal_6186}), .clk (clk), .r (Fresh[630]), .c ({signal_9595, signal_6307}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6072 ( .a ({signal_21896, signal_21890}), .b ({signal_9445, signal_6185}), .clk (clk), .r (Fresh[631]), .c ({signal_9596, signal_6308}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6073 ( .a ({signal_21908, signal_21902}), .b ({signal_9448, signal_6188}), .clk (clk), .r (Fresh[632]), .c ({signal_9597, signal_6309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6074 ( .a ({signal_21920, signal_21914}), .b ({signal_9447, signal_6187}), .clk (clk), .r (Fresh[633]), .c ({signal_9598, signal_6310}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6075 ( .a ({signal_21932, signal_21926}), .b ({signal_9446, signal_6186}), .clk (clk), .r (Fresh[634]), .c ({signal_9599, signal_6311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6076 ( .a ({signal_21944, signal_21938}), .b ({signal_9445, signal_6185}), .clk (clk), .r (Fresh[635]), .c ({signal_9600, signal_6312}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6077 ( .a ({signal_21956, signal_21950}), .b ({signal_9452, signal_6192}), .clk (clk), .r (Fresh[636]), .c ({signal_9601, signal_6313}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6078 ( .a ({signal_21968, signal_21962}), .b ({signal_9451, signal_6191}), .clk (clk), .r (Fresh[637]), .c ({signal_9602, signal_6314}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6079 ( .a ({signal_21980, signal_21974}), .b ({signal_9450, signal_6190}), .clk (clk), .r (Fresh[638]), .c ({signal_9603, signal_6315}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6080 ( .a ({signal_21992, signal_21986}), .b ({signal_9449, signal_6189}), .clk (clk), .r (Fresh[639]), .c ({signal_9604, signal_6316}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6081 ( .a ({signal_22004, signal_21998}), .b ({signal_9452, signal_6192}), .clk (clk), .r (Fresh[640]), .c ({signal_9605, signal_6317}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6082 ( .a ({signal_22016, signal_22010}), .b ({signal_9451, signal_6191}), .clk (clk), .r (Fresh[641]), .c ({signal_9606, signal_6318}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6083 ( .a ({signal_22028, signal_22022}), .b ({signal_9450, signal_6190}), .clk (clk), .r (Fresh[642]), .c ({signal_9607, signal_6319}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6084 ( .a ({signal_22040, signal_22034}), .b ({signal_9449, signal_6189}), .clk (clk), .r (Fresh[643]), .c ({signal_9608, signal_6320}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6085 ( .a ({signal_22052, signal_22046}), .b ({signal_9501, signal_6193}), .clk (clk), .r (Fresh[644]), .c ({signal_9705, signal_6321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6086 ( .a ({signal_22064, signal_22058}), .b ({signal_9501, signal_6193}), .clk (clk), .r (Fresh[645]), .c ({signal_9706, signal_6322}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6087 ( .a ({signal_22076, signal_22070}), .b ({signal_9453, signal_6197}), .clk (clk), .r (Fresh[646]), .c ({signal_9609, signal_6323}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6088 ( .a ({signal_22088, signal_22082}), .b ({signal_9453, signal_6197}), .clk (clk), .r (Fresh[647]), .c ({signal_9610, signal_6324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6089 ( .a ({signal_22100, signal_22094}), .b ({signal_9457, signal_6201}), .clk (clk), .r (Fresh[648]), .c ({signal_9611, signal_6325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6090 ( .a ({signal_22112, signal_22106}), .b ({signal_9457, signal_6201}), .clk (clk), .r (Fresh[649]), .c ({signal_9612, signal_6326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6091 ( .a ({signal_22124, signal_22118}), .b ({signal_9461, signal_6205}), .clk (clk), .r (Fresh[650]), .c ({signal_9613, signal_6327}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6092 ( .a ({signal_22136, signal_22130}), .b ({signal_9461, signal_6205}), .clk (clk), .r (Fresh[651]), .c ({signal_9614, signal_6328}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6093 ( .a ({signal_22148, signal_22142}), .b ({signal_9465, signal_6209}), .clk (clk), .r (Fresh[652]), .c ({signal_9615, signal_6329}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6094 ( .a ({signal_22160, signal_22154}), .b ({signal_9465, signal_6209}), .clk (clk), .r (Fresh[653]), .c ({signal_9616, signal_6330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6096 ( .a ({signal_9267, signal_5975}), .b ({signal_9269, signal_5977}), .c ({signal_9618, signal_6332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6097 ( .a ({signal_9268, signal_5976}), .b ({signal_9271, signal_5979}), .c ({signal_9619, signal_6333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6098 ( .a ({signal_9266, signal_5974}), .b ({signal_9268, signal_5976}), .c ({signal_9620, signal_6334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6100 ( .a ({signal_9275, signal_5983}), .b ({signal_9277, signal_5985}), .c ({signal_9622, signal_6336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6101 ( .a ({signal_9276, signal_5984}), .b ({signal_9279, signal_5987}), .c ({signal_9623, signal_6337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6102 ( .a ({signal_9274, signal_5982}), .b ({signal_9276, signal_5984}), .c ({signal_9624, signal_6338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6104 ( .a ({signal_9283, signal_5991}), .b ({signal_9285, signal_5993}), .c ({signal_9626, signal_6340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6105 ( .a ({signal_9284, signal_5992}), .b ({signal_9287, signal_5995}), .c ({signal_9627, signal_6341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6106 ( .a ({signal_9282, signal_5990}), .b ({signal_9284, signal_5992}), .c ({signal_9628, signal_6342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6108 ( .a ({signal_9291, signal_5999}), .b ({signal_9293, signal_6001}), .c ({signal_9630, signal_6344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6109 ( .a ({signal_9292, signal_6000}), .b ({signal_9295, signal_6003}), .c ({signal_9631, signal_6345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6110 ( .a ({signal_9290, signal_5998}), .b ({signal_9292, signal_6000}), .c ({signal_9632, signal_6346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6112 ( .a ({signal_9299, signal_6007}), .b ({signal_9301, signal_6009}), .c ({signal_9634, signal_6348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6113 ( .a ({signal_9300, signal_6008}), .b ({signal_9303, signal_6011}), .c ({signal_9635, signal_6349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6114 ( .a ({signal_9298, signal_6006}), .b ({signal_9300, signal_6008}), .c ({signal_9636, signal_6350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6116 ( .a ({signal_9307, signal_6015}), .b ({signal_9309, signal_6017}), .c ({signal_9638, signal_6352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6117 ( .a ({signal_9308, signal_6016}), .b ({signal_9311, signal_6019}), .c ({signal_9639, signal_6353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6118 ( .a ({signal_9306, signal_6014}), .b ({signal_9308, signal_6016}), .c ({signal_9640, signal_6354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6120 ( .a ({signal_9315, signal_6023}), .b ({signal_9317, signal_6025}), .c ({signal_9642, signal_6356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6121 ( .a ({signal_9316, signal_6024}), .b ({signal_9319, signal_6027}), .c ({signal_9643, signal_6357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6122 ( .a ({signal_9314, signal_6022}), .b ({signal_9316, signal_6024}), .c ({signal_9644, signal_6358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6123 ( .a ({signal_9230, signal_5838}), .b ({signal_9469, signal_6029}), .c ({signal_9707, signal_6359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6124 ( .a ({signal_9229, signal_5837}), .b ({signal_9473, signal_6033}), .c ({signal_9708, signal_6360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6125 ( .a ({signal_9472, signal_6032}), .b ({signal_9474, signal_6034}), .c ({signal_9709, signal_6361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6126 ( .a ({signal_9470, signal_6030}), .b ({signal_9475, signal_6035}), .c ({signal_9710, signal_6362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6127 ( .a ({signal_9471, signal_6031}), .b ({signal_9475, signal_6035}), .c ({signal_9711, signal_6363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6128 ( .a ({signal_9473, signal_6033}), .b ({signal_9494, signal_6162}), .c ({signal_9712, signal_6364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6129 ( .a ({signal_9234, signal_5842}), .b ({signal_9494, signal_6162}), .c ({signal_9713, signal_6365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6130 ( .a ({signal_9474, signal_6034}), .b ({signal_9495, signal_6163}), .c ({signal_9714, signal_6366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6132 ( .a ({signal_9323, signal_6039}), .b ({signal_9325, signal_6041}), .c ({signal_9646, signal_6368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6133 ( .a ({signal_9324, signal_6040}), .b ({signal_9327, signal_6043}), .c ({signal_9647, signal_6369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6134 ( .a ({signal_9322, signal_6038}), .b ({signal_9324, signal_6040}), .c ({signal_9648, signal_6370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6136 ( .a ({signal_9331, signal_6047}), .b ({signal_9333, signal_6049}), .c ({signal_9650, signal_6372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6137 ( .a ({signal_9332, signal_6048}), .b ({signal_9335, signal_6051}), .c ({signal_9651, signal_6373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6138 ( .a ({signal_9330, signal_6046}), .b ({signal_9332, signal_6048}), .c ({signal_9652, signal_6374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6140 ( .a ({signal_9339, signal_6055}), .b ({signal_9341, signal_6057}), .c ({signal_9654, signal_6376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6141 ( .a ({signal_9340, signal_6056}), .b ({signal_9343, signal_6059}), .c ({signal_9655, signal_6377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6142 ( .a ({signal_9338, signal_6054}), .b ({signal_9340, signal_6056}), .c ({signal_9656, signal_6378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6143 ( .a ({signal_9238, signal_5846}), .b ({signal_9477, signal_6061}), .c ({signal_9715, signal_6379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6144 ( .a ({signal_9237, signal_5845}), .b ({signal_9481, signal_6065}), .c ({signal_9716, signal_6380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6145 ( .a ({signal_9480, signal_6064}), .b ({signal_9482, signal_6066}), .c ({signal_9717, signal_6381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6146 ( .a ({signal_9478, signal_6062}), .b ({signal_9483, signal_6067}), .c ({signal_9718, signal_6382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6147 ( .a ({signal_9479, signal_6063}), .b ({signal_9483, signal_6067}), .c ({signal_9719, signal_6383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6148 ( .a ({signal_9481, signal_6065}), .b ({signal_9498, signal_6178}), .c ({signal_9720, signal_6384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6149 ( .a ({signal_9242, signal_5850}), .b ({signal_9498, signal_6178}), .c ({signal_9721, signal_6385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6150 ( .a ({signal_9482, signal_6066}), .b ({signal_9499, signal_6179}), .c ({signal_9722, signal_6386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6152 ( .a ({signal_9347, signal_6071}), .b ({signal_9349, signal_6073}), .c ({signal_9658, signal_6388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6153 ( .a ({signal_9348, signal_6072}), .b ({signal_9351, signal_6075}), .c ({signal_9659, signal_6389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6154 ( .a ({signal_9346, signal_6070}), .b ({signal_9348, signal_6072}), .c ({signal_9660, signal_6390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6156 ( .a ({signal_9355, signal_6079}), .b ({signal_9357, signal_6081}), .c ({signal_9662, signal_6392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6157 ( .a ({signal_9356, signal_6080}), .b ({signal_9359, signal_6083}), .c ({signal_9663, signal_6393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6158 ( .a ({signal_9354, signal_6078}), .b ({signal_9356, signal_6080}), .c ({signal_9664, signal_6394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6160 ( .a ({signal_9363, signal_6087}), .b ({signal_9365, signal_6089}), .c ({signal_9666, signal_6396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6161 ( .a ({signal_9364, signal_6088}), .b ({signal_9367, signal_6091}), .c ({signal_9667, signal_6397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6162 ( .a ({signal_9362, signal_6086}), .b ({signal_9364, signal_6088}), .c ({signal_9668, signal_6398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6163 ( .a ({signal_9246, signal_5854}), .b ({signal_9485, signal_6093}), .c ({signal_9723, signal_6399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6164 ( .a ({signal_9245, signal_5853}), .b ({signal_9489, signal_6097}), .c ({signal_9724, signal_6400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6165 ( .a ({signal_9488, signal_6096}), .b ({signal_9490, signal_6098}), .c ({signal_9725, signal_6401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6166 ( .a ({signal_9486, signal_6094}), .b ({signal_9491, signal_6099}), .c ({signal_9726, signal_6402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6167 ( .a ({signal_9487, signal_6095}), .b ({signal_9491, signal_6099}), .c ({signal_9727, signal_6403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6168 ( .a ({signal_9489, signal_6097}), .b ({signal_9502, signal_6194}), .c ({signal_9728, signal_6404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6169 ( .a ({signal_9250, signal_5858}), .b ({signal_9502, signal_6194}), .c ({signal_9729, signal_6405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6170 ( .a ({signal_9490, signal_6098}), .b ({signal_9503, signal_6195}), .c ({signal_9730, signal_6406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6171 ( .a ({signal_9130, signal_5862}), .b ({signal_9369, signal_6101}), .c ({signal_9669, signal_6407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6172 ( .a ({signal_9129, signal_5861}), .b ({signal_9373, signal_6105}), .c ({signal_9670, signal_6408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6173 ( .a ({signal_9372, signal_6104}), .b ({signal_9374, signal_6106}), .c ({signal_9671, signal_6409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6174 ( .a ({signal_9370, signal_6102}), .b ({signal_9375, signal_6107}), .c ({signal_9672, signal_6410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6175 ( .a ({signal_9371, signal_6103}), .b ({signal_9375, signal_6107}), .c ({signal_9673, signal_6411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6176 ( .a ({signal_9373, signal_6105}), .b ({signal_9454, signal_6198}), .c ({signal_9674, signal_6412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6177 ( .a ({signal_9134, signal_5866}), .b ({signal_9454, signal_6198}), .c ({signal_9675, signal_6413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6178 ( .a ({signal_9374, signal_6106}), .b ({signal_9455, signal_6199}), .c ({signal_9676, signal_6414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6179 ( .a ({signal_9138, signal_5870}), .b ({signal_9377, signal_6109}), .c ({signal_9677, signal_6415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6180 ( .a ({signal_9137, signal_5869}), .b ({signal_9381, signal_6113}), .c ({signal_9678, signal_6416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6181 ( .a ({signal_9380, signal_6112}), .b ({signal_9382, signal_6114}), .c ({signal_9679, signal_6417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6182 ( .a ({signal_9378, signal_6110}), .b ({signal_9383, signal_6115}), .c ({signal_9680, signal_6418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6183 ( .a ({signal_9379, signal_6111}), .b ({signal_9383, signal_6115}), .c ({signal_9681, signal_6419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6184 ( .a ({signal_9381, signal_6113}), .b ({signal_9458, signal_6202}), .c ({signal_9682, signal_6420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6185 ( .a ({signal_9142, signal_5874}), .b ({signal_9458, signal_6202}), .c ({signal_9683, signal_6421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6186 ( .a ({signal_9382, signal_6114}), .b ({signal_9459, signal_6203}), .c ({signal_9684, signal_6422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6187 ( .a ({signal_9146, signal_5878}), .b ({signal_9385, signal_6117}), .c ({signal_9685, signal_6423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6188 ( .a ({signal_9145, signal_5877}), .b ({signal_9389, signal_6121}), .c ({signal_9686, signal_6424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6189 ( .a ({signal_9388, signal_6120}), .b ({signal_9390, signal_6122}), .c ({signal_9687, signal_6425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6190 ( .a ({signal_9386, signal_6118}), .b ({signal_9391, signal_6123}), .c ({signal_9688, signal_6426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6191 ( .a ({signal_9387, signal_6119}), .b ({signal_9391, signal_6123}), .c ({signal_9689, signal_6427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6192 ( .a ({signal_9389, signal_6121}), .b ({signal_9462, signal_6206}), .c ({signal_9690, signal_6428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6193 ( .a ({signal_9150, signal_5882}), .b ({signal_9462, signal_6206}), .c ({signal_9691, signal_6429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6194 ( .a ({signal_9390, signal_6122}), .b ({signal_9463, signal_6207}), .c ({signal_9692, signal_6430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6195 ( .a ({signal_9154, signal_5886}), .b ({signal_9393, signal_6125}), .c ({signal_9693, signal_6431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6196 ( .a ({signal_9153, signal_5885}), .b ({signal_9397, signal_6129}), .c ({signal_9694, signal_6432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6197 ( .a ({signal_9396, signal_6128}), .b ({signal_9398, signal_6130}), .c ({signal_9695, signal_6433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6198 ( .a ({signal_9394, signal_6126}), .b ({signal_9399, signal_6131}), .c ({signal_9696, signal_6434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6199 ( .a ({signal_9395, signal_6127}), .b ({signal_9399, signal_6131}), .c ({signal_9697, signal_6435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6200 ( .a ({signal_9397, signal_6129}), .b ({signal_9466, signal_6210}), .c ({signal_9698, signal_6436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6201 ( .a ({signal_9158, signal_5890}), .b ({signal_9466, signal_6210}), .c ({signal_9699, signal_6437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6202 ( .a ({signal_9398, signal_6130}), .b ({signal_9467, signal_6211}), .c ({signal_9700, signal_6438}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6203 ( .a ({signal_22172, signal_22166}), .b ({signal_9617, signal_6331}), .clk (clk), .r (Fresh[654]), .c ({signal_9731, signal_6439}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6204 ( .a ({signal_22184, signal_22178}), .b ({signal_9617, signal_6331}), .clk (clk), .r (Fresh[655]), .c ({signal_9732, signal_6440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6205 ( .a ({signal_22196, signal_22190}), .b ({signal_9621, signal_6335}), .clk (clk), .r (Fresh[656]), .c ({signal_9733, signal_6441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6206 ( .a ({signal_22208, signal_22202}), .b ({signal_9621, signal_6335}), .clk (clk), .r (Fresh[657]), .c ({signal_9734, signal_6442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6207 ( .a ({signal_22220, signal_22214}), .b ({signal_9625, signal_6339}), .clk (clk), .r (Fresh[658]), .c ({signal_9735, signal_6443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6208 ( .a ({signal_22232, signal_22226}), .b ({signal_9625, signal_6339}), .clk (clk), .r (Fresh[659]), .c ({signal_9736, signal_6444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6209 ( .a ({signal_22244, signal_22238}), .b ({signal_9629, signal_6343}), .clk (clk), .r (Fresh[660]), .c ({signal_9737, signal_6445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6210 ( .a ({signal_22256, signal_22250}), .b ({signal_9629, signal_6343}), .clk (clk), .r (Fresh[661]), .c ({signal_9738, signal_6446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6211 ( .a ({signal_22268, signal_22262}), .b ({signal_9633, signal_6347}), .clk (clk), .r (Fresh[662]), .c ({signal_9739, signal_6447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6212 ( .a ({signal_22280, signal_22274}), .b ({signal_9633, signal_6347}), .clk (clk), .r (Fresh[663]), .c ({signal_9740, signal_6448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6213 ( .a ({signal_22292, signal_22286}), .b ({signal_9637, signal_6351}), .clk (clk), .r (Fresh[664]), .c ({signal_9741, signal_6449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6214 ( .a ({signal_22304, signal_22298}), .b ({signal_9637, signal_6351}), .clk (clk), .r (Fresh[665]), .c ({signal_9742, signal_6450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6215 ( .a ({signal_22316, signal_22310}), .b ({signal_9641, signal_6355}), .clk (clk), .r (Fresh[666]), .c ({signal_9743, signal_6451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6216 ( .a ({signal_22328, signal_22322}), .b ({signal_9641, signal_6355}), .clk (clk), .r (Fresh[667]), .c ({signal_9744, signal_6452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6217 ( .a ({signal_22340, signal_22334}), .b ({signal_9645, signal_6367}), .clk (clk), .r (Fresh[668]), .c ({signal_9745, signal_6453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6218 ( .a ({signal_22352, signal_22346}), .b ({signal_9645, signal_6367}), .clk (clk), .r (Fresh[669]), .c ({signal_9746, signal_6454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6219 ( .a ({signal_22364, signal_22358}), .b ({signal_9649, signal_6371}), .clk (clk), .r (Fresh[670]), .c ({signal_9747, signal_6455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6220 ( .a ({signal_22376, signal_22370}), .b ({signal_9649, signal_6371}), .clk (clk), .r (Fresh[671]), .c ({signal_9748, signal_6456}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6221 ( .a ({signal_22388, signal_22382}), .b ({signal_9653, signal_6375}), .clk (clk), .r (Fresh[672]), .c ({signal_9749, signal_6457}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6222 ( .a ({signal_22400, signal_22394}), .b ({signal_9653, signal_6375}), .clk (clk), .r (Fresh[673]), .c ({signal_9750, signal_6458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6223 ( .a ({signal_22412, signal_22406}), .b ({signal_9657, signal_6387}), .clk (clk), .r (Fresh[674]), .c ({signal_9751, signal_6459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6224 ( .a ({signal_22424, signal_22418}), .b ({signal_9657, signal_6387}), .clk (clk), .r (Fresh[675]), .c ({signal_9752, signal_6460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6225 ( .a ({signal_22436, signal_22430}), .b ({signal_9661, signal_6391}), .clk (clk), .r (Fresh[676]), .c ({signal_9753, signal_6461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6226 ( .a ({signal_22448, signal_22442}), .b ({signal_9661, signal_6391}), .clk (clk), .r (Fresh[677]), .c ({signal_9754, signal_6462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6227 ( .a ({signal_22460, signal_22454}), .b ({signal_9665, signal_6395}), .clk (clk), .r (Fresh[678]), .c ({signal_9755, signal_6463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_6228 ( .a ({signal_22472, signal_22466}), .b ({signal_9665, signal_6395}), .clk (clk), .r (Fresh[679]), .c ({signal_9756, signal_6464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6229 ( .a ({signal_9266, signal_5974}), .b ({signal_9505, signal_6213}), .c ({signal_9757, signal_6465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6230 ( .a ({signal_9265, signal_5973}), .b ({signal_9509, signal_6217}), .c ({signal_9758, signal_6466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6231 ( .a ({signal_9508, signal_6216}), .b ({signal_9510, signal_6218}), .c ({signal_9759, signal_6467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6232 ( .a ({signal_9506, signal_6214}), .b ({signal_9511, signal_6219}), .c ({signal_9760, signal_6468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6233 ( .a ({signal_9507, signal_6215}), .b ({signal_9511, signal_6219}), .c ({signal_9761, signal_6469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6234 ( .a ({signal_9509, signal_6217}), .b ({signal_9618, signal_6332}), .c ({signal_9762, signal_6470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6235 ( .a ({signal_9270, signal_5978}), .b ({signal_9618, signal_6332}), .c ({signal_9763, signal_6471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6236 ( .a ({signal_9510, signal_6218}), .b ({signal_9619, signal_6333}), .c ({signal_9764, signal_6472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6237 ( .a ({signal_9274, signal_5982}), .b ({signal_9513, signal_6221}), .c ({signal_9765, signal_6473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6238 ( .a ({signal_9273, signal_5981}), .b ({signal_9517, signal_6225}), .c ({signal_9766, signal_6474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6239 ( .a ({signal_9516, signal_6224}), .b ({signal_9518, signal_6226}), .c ({signal_9767, signal_6475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6240 ( .a ({signal_9514, signal_6222}), .b ({signal_9519, signal_6227}), .c ({signal_9768, signal_6476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6241 ( .a ({signal_9515, signal_6223}), .b ({signal_9519, signal_6227}), .c ({signal_9769, signal_6477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6242 ( .a ({signal_9517, signal_6225}), .b ({signal_9622, signal_6336}), .c ({signal_9770, signal_6478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6243 ( .a ({signal_9278, signal_5986}), .b ({signal_9622, signal_6336}), .c ({signal_9771, signal_6479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6244 ( .a ({signal_9518, signal_6226}), .b ({signal_9623, signal_6337}), .c ({signal_9772, signal_6480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6245 ( .a ({signal_9282, signal_5990}), .b ({signal_9521, signal_6229}), .c ({signal_9773, signal_6481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6246 ( .a ({signal_9281, signal_5989}), .b ({signal_9525, signal_6233}), .c ({signal_9774, signal_6482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6247 ( .a ({signal_9524, signal_6232}), .b ({signal_9526, signal_6234}), .c ({signal_9775, signal_6483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6248 ( .a ({signal_9522, signal_6230}), .b ({signal_9527, signal_6235}), .c ({signal_9776, signal_6484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6249 ( .a ({signal_9523, signal_6231}), .b ({signal_9527, signal_6235}), .c ({signal_9777, signal_6485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6250 ( .a ({signal_9525, signal_6233}), .b ({signal_9626, signal_6340}), .c ({signal_9778, signal_6486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6251 ( .a ({signal_9286, signal_5994}), .b ({signal_9626, signal_6340}), .c ({signal_9779, signal_6487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6252 ( .a ({signal_9526, signal_6234}), .b ({signal_9627, signal_6341}), .c ({signal_9780, signal_6488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6253 ( .a ({signal_9290, signal_5998}), .b ({signal_9529, signal_6237}), .c ({signal_9781, signal_6489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6254 ( .a ({signal_9289, signal_5997}), .b ({signal_9533, signal_6241}), .c ({signal_9782, signal_6490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6255 ( .a ({signal_9532, signal_6240}), .b ({signal_9534, signal_6242}), .c ({signal_9783, signal_6491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6256 ( .a ({signal_9530, signal_6238}), .b ({signal_9535, signal_6243}), .c ({signal_9784, signal_6492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6257 ( .a ({signal_9531, signal_6239}), .b ({signal_9535, signal_6243}), .c ({signal_9785, signal_6493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6258 ( .a ({signal_9533, signal_6241}), .b ({signal_9630, signal_6344}), .c ({signal_9786, signal_6494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6259 ( .a ({signal_9294, signal_6002}), .b ({signal_9630, signal_6344}), .c ({signal_9787, signal_6495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6260 ( .a ({signal_9534, signal_6242}), .b ({signal_9631, signal_6345}), .c ({signal_9788, signal_6496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6261 ( .a ({signal_9298, signal_6006}), .b ({signal_9537, signal_6245}), .c ({signal_9789, signal_6497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6262 ( .a ({signal_9297, signal_6005}), .b ({signal_9541, signal_6249}), .c ({signal_9790, signal_6498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6263 ( .a ({signal_9540, signal_6248}), .b ({signal_9542, signal_6250}), .c ({signal_9791, signal_6499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6264 ( .a ({signal_9538, signal_6246}), .b ({signal_9543, signal_6251}), .c ({signal_9792, signal_6500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6265 ( .a ({signal_9539, signal_6247}), .b ({signal_9543, signal_6251}), .c ({signal_9793, signal_6501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6266 ( .a ({signal_9541, signal_6249}), .b ({signal_9634, signal_6348}), .c ({signal_9794, signal_6502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6267 ( .a ({signal_9302, signal_6010}), .b ({signal_9634, signal_6348}), .c ({signal_9795, signal_6503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6268 ( .a ({signal_9542, signal_6250}), .b ({signal_9635, signal_6349}), .c ({signal_9796, signal_6504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6269 ( .a ({signal_9306, signal_6014}), .b ({signal_9545, signal_6253}), .c ({signal_9797, signal_6505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6270 ( .a ({signal_9305, signal_6013}), .b ({signal_9549, signal_6257}), .c ({signal_9798, signal_6506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6271 ( .a ({signal_9548, signal_6256}), .b ({signal_9550, signal_6258}), .c ({signal_9799, signal_6507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6272 ( .a ({signal_9546, signal_6254}), .b ({signal_9551, signal_6259}), .c ({signal_9800, signal_6508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6273 ( .a ({signal_9547, signal_6255}), .b ({signal_9551, signal_6259}), .c ({signal_9801, signal_6509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6274 ( .a ({signal_9549, signal_6257}), .b ({signal_9638, signal_6352}), .c ({signal_9802, signal_6510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6275 ( .a ({signal_9310, signal_6018}), .b ({signal_9638, signal_6352}), .c ({signal_9803, signal_6511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6276 ( .a ({signal_9550, signal_6258}), .b ({signal_9639, signal_6353}), .c ({signal_9804, signal_6512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6277 ( .a ({signal_9314, signal_6022}), .b ({signal_9553, signal_6261}), .c ({signal_9805, signal_6513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6278 ( .a ({signal_9313, signal_6021}), .b ({signal_9557, signal_6265}), .c ({signal_9806, signal_6514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6279 ( .a ({signal_9556, signal_6264}), .b ({signal_9558, signal_6266}), .c ({signal_9807, signal_6515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6280 ( .a ({signal_9554, signal_6262}), .b ({signal_9559, signal_6267}), .c ({signal_9808, signal_6516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6281 ( .a ({signal_9555, signal_6263}), .b ({signal_9559, signal_6267}), .c ({signal_9809, signal_6517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6282 ( .a ({signal_9557, signal_6265}), .b ({signal_9642, signal_6356}), .c ({signal_9810, signal_6518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6283 ( .a ({signal_9318, signal_6026}), .b ({signal_9642, signal_6356}), .c ({signal_9811, signal_6519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6284 ( .a ({signal_9558, signal_6266}), .b ({signal_9643, signal_6357}), .c ({signal_9812, signal_6520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6285 ( .a ({signal_9475, signal_6035}), .b ({signal_9702, signal_6270}), .c ({signal_9897, signal_6521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6286 ( .a ({signal_9702, signal_6270}), .b ({signal_9710, signal_6362}), .c ({signal_9898, signal_6522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6287 ( .a ({signal_9469, signal_6029}), .b ({signal_9708, signal_6360}), .c ({signal_9899, signal_6523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6288 ( .a ({signal_9471, signal_6031}), .b ({signal_9701, signal_6269}), .c ({signal_9900, signal_6524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6289 ( .a ({signal_9701, signal_6269}), .b ({signal_9709, signal_6361}), .c ({signal_9901, signal_6525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6290 ( .a ({signal_9236, signal_5844}), .b ({signal_9707, signal_6359}), .c ({signal_9902, signal_6526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6291 ( .a ({signal_9476, signal_6036}), .b ({signal_9709, signal_6361}), .c ({signal_9903, signal_6527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6292 ( .a ({signal_9496, signal_6164}), .b ({signal_9708, signal_6360}), .c ({signal_9904, signal_6528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6293 ( .a ({signal_9707, signal_6359}), .b ({signal_9714, signal_6366}), .c ({signal_9905, signal_6529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6294 ( .a ({signal_9322, signal_6038}), .b ({signal_9561, signal_6271}), .c ({signal_9813, signal_6530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6295 ( .a ({signal_9321, signal_6037}), .b ({signal_9565, signal_6275}), .c ({signal_9814, signal_6531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6296 ( .a ({signal_9564, signal_6274}), .b ({signal_9566, signal_6276}), .c ({signal_9815, signal_6532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6297 ( .a ({signal_9562, signal_6272}), .b ({signal_9567, signal_6277}), .c ({signal_9816, signal_6533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6298 ( .a ({signal_9563, signal_6273}), .b ({signal_9567, signal_6277}), .c ({signal_9817, signal_6534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6299 ( .a ({signal_9565, signal_6275}), .b ({signal_9646, signal_6368}), .c ({signal_9818, signal_6535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6300 ( .a ({signal_9326, signal_6042}), .b ({signal_9646, signal_6368}), .c ({signal_9819, signal_6536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6301 ( .a ({signal_9566, signal_6276}), .b ({signal_9647, signal_6369}), .c ({signal_9820, signal_6537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6302 ( .a ({signal_9330, signal_6046}), .b ({signal_9569, signal_6279}), .c ({signal_9821, signal_6538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6303 ( .a ({signal_9329, signal_6045}), .b ({signal_9573, signal_6283}), .c ({signal_9822, signal_6539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6304 ( .a ({signal_9572, signal_6282}), .b ({signal_9574, signal_6284}), .c ({signal_9823, signal_6540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6305 ( .a ({signal_9570, signal_6280}), .b ({signal_9575, signal_6285}), .c ({signal_9824, signal_6541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6306 ( .a ({signal_9571, signal_6281}), .b ({signal_9575, signal_6285}), .c ({signal_9825, signal_6542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6307 ( .a ({signal_9573, signal_6283}), .b ({signal_9650, signal_6372}), .c ({signal_9826, signal_6543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6308 ( .a ({signal_9334, signal_6050}), .b ({signal_9650, signal_6372}), .c ({signal_9827, signal_6544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6309 ( .a ({signal_9574, signal_6284}), .b ({signal_9651, signal_6373}), .c ({signal_9828, signal_6545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6310 ( .a ({signal_9338, signal_6054}), .b ({signal_9577, signal_6287}), .c ({signal_9829, signal_6546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6311 ( .a ({signal_9337, signal_6053}), .b ({signal_9581, signal_6291}), .c ({signal_9830, signal_6547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6312 ( .a ({signal_9580, signal_6290}), .b ({signal_9582, signal_6292}), .c ({signal_9831, signal_6548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6313 ( .a ({signal_9578, signal_6288}), .b ({signal_9583, signal_6293}), .c ({signal_9832, signal_6549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6314 ( .a ({signal_9579, signal_6289}), .b ({signal_9583, signal_6293}), .c ({signal_9833, signal_6550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6315 ( .a ({signal_9581, signal_6291}), .b ({signal_9654, signal_6376}), .c ({signal_9834, signal_6551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6316 ( .a ({signal_9342, signal_6058}), .b ({signal_9654, signal_6376}), .c ({signal_9835, signal_6552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6317 ( .a ({signal_9582, signal_6292}), .b ({signal_9655, signal_6377}), .c ({signal_9836, signal_6553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6318 ( .a ({signal_9483, signal_6067}), .b ({signal_9704, signal_6296}), .c ({signal_9906, signal_6554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6319 ( .a ({signal_9704, signal_6296}), .b ({signal_9718, signal_6382}), .c ({signal_9907, signal_6555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6320 ( .a ({signal_9477, signal_6061}), .b ({signal_9716, signal_6380}), .c ({signal_9908, signal_6556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6321 ( .a ({signal_9479, signal_6063}), .b ({signal_9703, signal_6295}), .c ({signal_9909, signal_6557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6322 ( .a ({signal_9703, signal_6295}), .b ({signal_9717, signal_6381}), .c ({signal_9910, signal_6558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6323 ( .a ({signal_9244, signal_5852}), .b ({signal_9715, signal_6379}), .c ({signal_9911, signal_6559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6324 ( .a ({signal_9484, signal_6068}), .b ({signal_9717, signal_6381}), .c ({signal_9912, signal_6560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6325 ( .a ({signal_9500, signal_6180}), .b ({signal_9716, signal_6380}), .c ({signal_9913, signal_6561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6326 ( .a ({signal_9715, signal_6379}), .b ({signal_9722, signal_6386}), .c ({signal_9914, signal_6562}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6327 ( .a ({signal_9346, signal_6070}), .b ({signal_9585, signal_6297}), .c ({signal_9837, signal_6563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6328 ( .a ({signal_9345, signal_6069}), .b ({signal_9589, signal_6301}), .c ({signal_9838, signal_6564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6329 ( .a ({signal_9588, signal_6300}), .b ({signal_9590, signal_6302}), .c ({signal_9839, signal_6565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6330 ( .a ({signal_9586, signal_6298}), .b ({signal_9591, signal_6303}), .c ({signal_9840, signal_6566}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6331 ( .a ({signal_9587, signal_6299}), .b ({signal_9591, signal_6303}), .c ({signal_9841, signal_6567}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6332 ( .a ({signal_9589, signal_6301}), .b ({signal_9658, signal_6388}), .c ({signal_9842, signal_6568}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6333 ( .a ({signal_9350, signal_6074}), .b ({signal_9658, signal_6388}), .c ({signal_9843, signal_6569}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6334 ( .a ({signal_9590, signal_6302}), .b ({signal_9659, signal_6389}), .c ({signal_9844, signal_6570}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6335 ( .a ({signal_9354, signal_6078}), .b ({signal_9593, signal_6305}), .c ({signal_9845, signal_6571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6336 ( .a ({signal_9353, signal_6077}), .b ({signal_9597, signal_6309}), .c ({signal_9846, signal_6572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6337 ( .a ({signal_9596, signal_6308}), .b ({signal_9598, signal_6310}), .c ({signal_9847, signal_6573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6338 ( .a ({signal_9594, signal_6306}), .b ({signal_9599, signal_6311}), .c ({signal_9848, signal_6574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6339 ( .a ({signal_9595, signal_6307}), .b ({signal_9599, signal_6311}), .c ({signal_9849, signal_6575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6340 ( .a ({signal_9597, signal_6309}), .b ({signal_9662, signal_6392}), .c ({signal_9850, signal_6576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6341 ( .a ({signal_9358, signal_6082}), .b ({signal_9662, signal_6392}), .c ({signal_9851, signal_6577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6342 ( .a ({signal_9598, signal_6310}), .b ({signal_9663, signal_6393}), .c ({signal_9852, signal_6578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6343 ( .a ({signal_9362, signal_6086}), .b ({signal_9601, signal_6313}), .c ({signal_9853, signal_6579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6344 ( .a ({signal_9361, signal_6085}), .b ({signal_9605, signal_6317}), .c ({signal_9854, signal_6580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6345 ( .a ({signal_9604, signal_6316}), .b ({signal_9606, signal_6318}), .c ({signal_9855, signal_6581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6346 ( .a ({signal_9602, signal_6314}), .b ({signal_9607, signal_6319}), .c ({signal_9856, signal_6582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6347 ( .a ({signal_9603, signal_6315}), .b ({signal_9607, signal_6319}), .c ({signal_9857, signal_6583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6348 ( .a ({signal_9605, signal_6317}), .b ({signal_9666, signal_6396}), .c ({signal_9858, signal_6584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6349 ( .a ({signal_9366, signal_6090}), .b ({signal_9666, signal_6396}), .c ({signal_9859, signal_6585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6350 ( .a ({signal_9606, signal_6318}), .b ({signal_9667, signal_6397}), .c ({signal_9860, signal_6586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6351 ( .a ({signal_9491, signal_6099}), .b ({signal_9706, signal_6322}), .c ({signal_9915, signal_6587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6352 ( .a ({signal_9706, signal_6322}), .b ({signal_9726, signal_6402}), .c ({signal_9916, signal_6588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6353 ( .a ({signal_9485, signal_6093}), .b ({signal_9724, signal_6400}), .c ({signal_9917, signal_6589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6354 ( .a ({signal_9487, signal_6095}), .b ({signal_9705, signal_6321}), .c ({signal_9918, signal_6590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6355 ( .a ({signal_9705, signal_6321}), .b ({signal_9725, signal_6401}), .c ({signal_9919, signal_6591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6356 ( .a ({signal_9252, signal_5860}), .b ({signal_9723, signal_6399}), .c ({signal_9920, signal_6592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6357 ( .a ({signal_9492, signal_6100}), .b ({signal_9725, signal_6401}), .c ({signal_9921, signal_6593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6358 ( .a ({signal_9504, signal_6196}), .b ({signal_9724, signal_6400}), .c ({signal_9922, signal_6594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6359 ( .a ({signal_9723, signal_6399}), .b ({signal_9730, signal_6406}), .c ({signal_9923, signal_6595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6360 ( .a ({signal_9375, signal_6107}), .b ({signal_9610, signal_6324}), .c ({signal_9861, signal_6596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6361 ( .a ({signal_9610, signal_6324}), .b ({signal_9672, signal_6410}), .c ({signal_9862, signal_6597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6362 ( .a ({signal_9369, signal_6101}), .b ({signal_9670, signal_6408}), .c ({signal_9863, signal_6598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6363 ( .a ({signal_9371, signal_6103}), .b ({signal_9609, signal_6323}), .c ({signal_9864, signal_6599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6364 ( .a ({signal_9609, signal_6323}), .b ({signal_9671, signal_6409}), .c ({signal_9865, signal_6600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6365 ( .a ({signal_9136, signal_5868}), .b ({signal_9669, signal_6407}), .c ({signal_9866, signal_6601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6366 ( .a ({signal_9376, signal_6108}), .b ({signal_9671, signal_6409}), .c ({signal_9867, signal_6602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6367 ( .a ({signal_9456, signal_6200}), .b ({signal_9670, signal_6408}), .c ({signal_9868, signal_6603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6368 ( .a ({signal_9669, signal_6407}), .b ({signal_9676, signal_6414}), .c ({signal_9869, signal_6604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6369 ( .a ({signal_9383, signal_6115}), .b ({signal_9612, signal_6326}), .c ({signal_9870, signal_6605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6370 ( .a ({signal_9612, signal_6326}), .b ({signal_9680, signal_6418}), .c ({signal_9871, signal_6606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6371 ( .a ({signal_9377, signal_6109}), .b ({signal_9678, signal_6416}), .c ({signal_9872, signal_6607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6372 ( .a ({signal_9379, signal_6111}), .b ({signal_9611, signal_6325}), .c ({signal_9873, signal_6608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6373 ( .a ({signal_9611, signal_6325}), .b ({signal_9679, signal_6417}), .c ({signal_9874, signal_6609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6374 ( .a ({signal_9144, signal_5876}), .b ({signal_9677, signal_6415}), .c ({signal_9875, signal_6610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6375 ( .a ({signal_9384, signal_6116}), .b ({signal_9679, signal_6417}), .c ({signal_9876, signal_6611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6376 ( .a ({signal_9460, signal_6204}), .b ({signal_9678, signal_6416}), .c ({signal_9877, signal_6612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6377 ( .a ({signal_9677, signal_6415}), .b ({signal_9684, signal_6422}), .c ({signal_9878, signal_6613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6378 ( .a ({signal_9391, signal_6123}), .b ({signal_9614, signal_6328}), .c ({signal_9879, signal_6614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6379 ( .a ({signal_9614, signal_6328}), .b ({signal_9688, signal_6426}), .c ({signal_9880, signal_6615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6380 ( .a ({signal_9385, signal_6117}), .b ({signal_9686, signal_6424}), .c ({signal_9881, signal_6616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6381 ( .a ({signal_9387, signal_6119}), .b ({signal_9613, signal_6327}), .c ({signal_9882, signal_6617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6382 ( .a ({signal_9613, signal_6327}), .b ({signal_9687, signal_6425}), .c ({signal_9883, signal_6618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6383 ( .a ({signal_9152, signal_5884}), .b ({signal_9685, signal_6423}), .c ({signal_9884, signal_6619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6384 ( .a ({signal_9392, signal_6124}), .b ({signal_9687, signal_6425}), .c ({signal_9885, signal_6620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6385 ( .a ({signal_9464, signal_6208}), .b ({signal_9686, signal_6424}), .c ({signal_9886, signal_6621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6386 ( .a ({signal_9685, signal_6423}), .b ({signal_9692, signal_6430}), .c ({signal_9887, signal_6622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6387 ( .a ({signal_9399, signal_6131}), .b ({signal_9616, signal_6330}), .c ({signal_9888, signal_6623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6388 ( .a ({signal_9616, signal_6330}), .b ({signal_9696, signal_6434}), .c ({signal_9889, signal_6624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6389 ( .a ({signal_9393, signal_6125}), .b ({signal_9694, signal_6432}), .c ({signal_9890, signal_6625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6390 ( .a ({signal_9395, signal_6127}), .b ({signal_9615, signal_6329}), .c ({signal_9891, signal_6626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6391 ( .a ({signal_9615, signal_6329}), .b ({signal_9695, signal_6433}), .c ({signal_9892, signal_6627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6392 ( .a ({signal_9160, signal_5892}), .b ({signal_9693, signal_6431}), .c ({signal_9893, signal_6628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6393 ( .a ({signal_9400, signal_6132}), .b ({signal_9695, signal_6433}), .c ({signal_9894, signal_6629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6394 ( .a ({signal_9468, signal_6212}), .b ({signal_9694, signal_6432}), .c ({signal_9895, signal_6630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6395 ( .a ({signal_9693, signal_6431}), .b ({signal_9700, signal_6438}), .c ({signal_9896, signal_6631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6396 ( .a ({signal_9511, signal_6219}), .b ({signal_9732, signal_6440}), .c ({signal_9924, signal_6632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6397 ( .a ({signal_9732, signal_6440}), .b ({signal_9760, signal_6468}), .c ({signal_9925, signal_6633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6398 ( .a ({signal_9505, signal_6213}), .b ({signal_9758, signal_6466}), .c ({signal_9926, signal_6634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6399 ( .a ({signal_9507, signal_6215}), .b ({signal_9731, signal_6439}), .c ({signal_9927, signal_6635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6400 ( .a ({signal_9731, signal_6439}), .b ({signal_9759, signal_6467}), .c ({signal_9928, signal_6636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6401 ( .a ({signal_9272, signal_5980}), .b ({signal_9757, signal_6465}), .c ({signal_9929, signal_6637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6402 ( .a ({signal_9512, signal_6220}), .b ({signal_9759, signal_6467}), .c ({signal_9930, signal_6638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6403 ( .a ({signal_9620, signal_6334}), .b ({signal_9758, signal_6466}), .c ({signal_9931, signal_6639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6404 ( .a ({signal_9757, signal_6465}), .b ({signal_9764, signal_6472}), .c ({signal_9932, signal_6640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6405 ( .a ({signal_9519, signal_6227}), .b ({signal_9734, signal_6442}), .c ({signal_9933, signal_6641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6406 ( .a ({signal_9734, signal_6442}), .b ({signal_9768, signal_6476}), .c ({signal_9934, signal_6642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6407 ( .a ({signal_9513, signal_6221}), .b ({signal_9766, signal_6474}), .c ({signal_9935, signal_6643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6408 ( .a ({signal_9515, signal_6223}), .b ({signal_9733, signal_6441}), .c ({signal_9936, signal_6644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6409 ( .a ({signal_9733, signal_6441}), .b ({signal_9767, signal_6475}), .c ({signal_9937, signal_6645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6410 ( .a ({signal_9280, signal_5988}), .b ({signal_9765, signal_6473}), .c ({signal_9938, signal_6646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6411 ( .a ({signal_9520, signal_6228}), .b ({signal_9767, signal_6475}), .c ({signal_9939, signal_6647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6412 ( .a ({signal_9624, signal_6338}), .b ({signal_9766, signal_6474}), .c ({signal_9940, signal_6648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6413 ( .a ({signal_9765, signal_6473}), .b ({signal_9772, signal_6480}), .c ({signal_9941, signal_6649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6414 ( .a ({signal_9527, signal_6235}), .b ({signal_9736, signal_6444}), .c ({signal_9942, signal_6650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6415 ( .a ({signal_9736, signal_6444}), .b ({signal_9776, signal_6484}), .c ({signal_9943, signal_6651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6416 ( .a ({signal_9521, signal_6229}), .b ({signal_9774, signal_6482}), .c ({signal_9944, signal_6652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6417 ( .a ({signal_9523, signal_6231}), .b ({signal_9735, signal_6443}), .c ({signal_9945, signal_6653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6418 ( .a ({signal_9735, signal_6443}), .b ({signal_9775, signal_6483}), .c ({signal_9946, signal_6654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6419 ( .a ({signal_9288, signal_5996}), .b ({signal_9773, signal_6481}), .c ({signal_9947, signal_6655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6420 ( .a ({signal_9528, signal_6236}), .b ({signal_9775, signal_6483}), .c ({signal_9948, signal_6656}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6421 ( .a ({signal_9628, signal_6342}), .b ({signal_9774, signal_6482}), .c ({signal_9949, signal_6657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6422 ( .a ({signal_9773, signal_6481}), .b ({signal_9780, signal_6488}), .c ({signal_9950, signal_6658}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6423 ( .a ({signal_9535, signal_6243}), .b ({signal_9738, signal_6446}), .c ({signal_9951, signal_6659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6424 ( .a ({signal_9738, signal_6446}), .b ({signal_9784, signal_6492}), .c ({signal_9952, signal_6660}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6425 ( .a ({signal_9529, signal_6237}), .b ({signal_9782, signal_6490}), .c ({signal_9953, signal_6661}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6426 ( .a ({signal_9531, signal_6239}), .b ({signal_9737, signal_6445}), .c ({signal_9954, signal_6662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6427 ( .a ({signal_9737, signal_6445}), .b ({signal_9783, signal_6491}), .c ({signal_9955, signal_6663}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6428 ( .a ({signal_9296, signal_6004}), .b ({signal_9781, signal_6489}), .c ({signal_9956, signal_6664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6429 ( .a ({signal_9536, signal_6244}), .b ({signal_9783, signal_6491}), .c ({signal_9957, signal_6665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6430 ( .a ({signal_9632, signal_6346}), .b ({signal_9782, signal_6490}), .c ({signal_9958, signal_6666}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6431 ( .a ({signal_9781, signal_6489}), .b ({signal_9788, signal_6496}), .c ({signal_9959, signal_6667}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6432 ( .a ({signal_9543, signal_6251}), .b ({signal_9740, signal_6448}), .c ({signal_9960, signal_6668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6433 ( .a ({signal_9740, signal_6448}), .b ({signal_9792, signal_6500}), .c ({signal_9961, signal_6669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6434 ( .a ({signal_9537, signal_6245}), .b ({signal_9790, signal_6498}), .c ({signal_9962, signal_6670}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6435 ( .a ({signal_9539, signal_6247}), .b ({signal_9739, signal_6447}), .c ({signal_9963, signal_6671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6436 ( .a ({signal_9739, signal_6447}), .b ({signal_9791, signal_6499}), .c ({signal_9964, signal_6672}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6437 ( .a ({signal_9304, signal_6012}), .b ({signal_9789, signal_6497}), .c ({signal_9965, signal_6673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6438 ( .a ({signal_9544, signal_6252}), .b ({signal_9791, signal_6499}), .c ({signal_9966, signal_6674}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6439 ( .a ({signal_9636, signal_6350}), .b ({signal_9790, signal_6498}), .c ({signal_9967, signal_6675}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6440 ( .a ({signal_9789, signal_6497}), .b ({signal_9796, signal_6504}), .c ({signal_9968, signal_6676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6441 ( .a ({signal_9551, signal_6259}), .b ({signal_9742, signal_6450}), .c ({signal_9969, signal_6677}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6442 ( .a ({signal_9742, signal_6450}), .b ({signal_9800, signal_6508}), .c ({signal_9970, signal_6678}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6443 ( .a ({signal_9545, signal_6253}), .b ({signal_9798, signal_6506}), .c ({signal_9971, signal_6679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6444 ( .a ({signal_9547, signal_6255}), .b ({signal_9741, signal_6449}), .c ({signal_9972, signal_6680}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6445 ( .a ({signal_9741, signal_6449}), .b ({signal_9799, signal_6507}), .c ({signal_9973, signal_6681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6446 ( .a ({signal_9312, signal_6020}), .b ({signal_9797, signal_6505}), .c ({signal_9974, signal_6682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6447 ( .a ({signal_9552, signal_6260}), .b ({signal_9799, signal_6507}), .c ({signal_9975, signal_6683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6448 ( .a ({signal_9640, signal_6354}), .b ({signal_9798, signal_6506}), .c ({signal_9976, signal_6684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6449 ( .a ({signal_9797, signal_6505}), .b ({signal_9804, signal_6512}), .c ({signal_9977, signal_6685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6450 ( .a ({signal_9559, signal_6267}), .b ({signal_9744, signal_6452}), .c ({signal_9978, signal_6686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6451 ( .a ({signal_9744, signal_6452}), .b ({signal_9808, signal_6516}), .c ({signal_9979, signal_6687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6452 ( .a ({signal_9553, signal_6261}), .b ({signal_9806, signal_6514}), .c ({signal_9980, signal_6688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6453 ( .a ({signal_9555, signal_6263}), .b ({signal_9743, signal_6451}), .c ({signal_9981, signal_6689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6454 ( .a ({signal_9743, signal_6451}), .b ({signal_9807, signal_6515}), .c ({signal_9982, signal_6690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6455 ( .a ({signal_9320, signal_6028}), .b ({signal_9805, signal_6513}), .c ({signal_9983, signal_6691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6456 ( .a ({signal_9560, signal_6268}), .b ({signal_9807, signal_6515}), .c ({signal_9984, signal_6692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6457 ( .a ({signal_9644, signal_6358}), .b ({signal_9806, signal_6514}), .c ({signal_9985, signal_6693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6458 ( .a ({signal_9805, signal_6513}), .b ({signal_9812, signal_6520}), .c ({signal_9986, signal_6694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6459 ( .a ({signal_9231, signal_5839}), .b ({signal_9897, signal_6521}), .c ({signal_10085, signal_6695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6460 ( .a ({signal_9233, signal_5841}), .b ({signal_9897, signal_6521}), .c ({signal_10086, signal_6696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6461 ( .a ({signal_9494, signal_6162}), .b ({signal_9897, signal_6521}), .c ({signal_10087, signal_6697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6462 ( .a ({signal_9494, signal_6162}), .b ({signal_9899, signal_6523}), .c ({signal_10088, signal_6698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6463 ( .a ({signal_9712, signal_6364}), .b ({signal_9900, signal_6524}), .c ({signal_10089, signal_6699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6464 ( .a ({signal_9898, signal_6522}), .b ({signal_9901, signal_6525}), .c ({signal_10090, signal_6700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6465 ( .a ({signal_9899, signal_6523}), .b ({signal_9900, signal_6524}), .c ({signal_10091, signal_6701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6466 ( .a ({signal_9495, signal_6163}), .b ({signal_9901, signal_6525}), .c ({signal_10092, signal_6702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6467 ( .a ({signal_9711, signal_6363}), .b ({signal_9902, signal_6526}), .c ({signal_10093, signal_6703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6468 ( .a ({signal_9713, signal_6365}), .b ({signal_9902, signal_6526}), .c ({signal_10094, signal_6704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6469 ( .a ({signal_9898, signal_6522}), .b ({signal_9905, signal_6529}), .c ({signal_10095, signal_6705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6470 ( .a ({signal_9567, signal_6277}), .b ({signal_9746, signal_6454}), .c ({signal_9987, signal_6706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6471 ( .a ({signal_9746, signal_6454}), .b ({signal_9816, signal_6533}), .c ({signal_9988, signal_6707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6472 ( .a ({signal_9561, signal_6271}), .b ({signal_9814, signal_6531}), .c ({signal_9989, signal_6708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6473 ( .a ({signal_9563, signal_6273}), .b ({signal_9745, signal_6453}), .c ({signal_9990, signal_6709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6474 ( .a ({signal_9745, signal_6453}), .b ({signal_9815, signal_6532}), .c ({signal_9991, signal_6710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6475 ( .a ({signal_9328, signal_6044}), .b ({signal_9813, signal_6530}), .c ({signal_9992, signal_6711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6476 ( .a ({signal_9568, signal_6278}), .b ({signal_9815, signal_6532}), .c ({signal_9993, signal_6712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6477 ( .a ({signal_9648, signal_6370}), .b ({signal_9814, signal_6531}), .c ({signal_9994, signal_6713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6478 ( .a ({signal_9813, signal_6530}), .b ({signal_9820, signal_6537}), .c ({signal_9995, signal_6714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6479 ( .a ({signal_9575, signal_6285}), .b ({signal_9748, signal_6456}), .c ({signal_9996, signal_6715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6480 ( .a ({signal_9748, signal_6456}), .b ({signal_9824, signal_6541}), .c ({signal_9997, signal_6716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6481 ( .a ({signal_9569, signal_6279}), .b ({signal_9822, signal_6539}), .c ({signal_9998, signal_6717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6482 ( .a ({signal_9571, signal_6281}), .b ({signal_9747, signal_6455}), .c ({signal_9999, signal_6718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6483 ( .a ({signal_9747, signal_6455}), .b ({signal_9823, signal_6540}), .c ({signal_10000, signal_6719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6484 ( .a ({signal_9336, signal_6052}), .b ({signal_9821, signal_6538}), .c ({signal_10001, signal_6720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6485 ( .a ({signal_9576, signal_6286}), .b ({signal_9823, signal_6540}), .c ({signal_10002, signal_6721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6486 ( .a ({signal_9652, signal_6374}), .b ({signal_9822, signal_6539}), .c ({signal_10003, signal_6722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6487 ( .a ({signal_9821, signal_6538}), .b ({signal_9828, signal_6545}), .c ({signal_10004, signal_6723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6488 ( .a ({signal_9583, signal_6293}), .b ({signal_9750, signal_6458}), .c ({signal_10005, signal_6724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6489 ( .a ({signal_9750, signal_6458}), .b ({signal_9832, signal_6549}), .c ({signal_10006, signal_6725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6490 ( .a ({signal_9577, signal_6287}), .b ({signal_9830, signal_6547}), .c ({signal_10007, signal_6726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6491 ( .a ({signal_9579, signal_6289}), .b ({signal_9749, signal_6457}), .c ({signal_10008, signal_6727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6492 ( .a ({signal_9749, signal_6457}), .b ({signal_9831, signal_6548}), .c ({signal_10009, signal_6728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6493 ( .a ({signal_9344, signal_6060}), .b ({signal_9829, signal_6546}), .c ({signal_10010, signal_6729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6494 ( .a ({signal_9584, signal_6294}), .b ({signal_9831, signal_6548}), .c ({signal_10011, signal_6730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6495 ( .a ({signal_9656, signal_6378}), .b ({signal_9830, signal_6547}), .c ({signal_10012, signal_6731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6496 ( .a ({signal_9829, signal_6546}), .b ({signal_9836, signal_6553}), .c ({signal_10013, signal_6732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6497 ( .a ({signal_9239, signal_5847}), .b ({signal_9906, signal_6554}), .c ({signal_10096, signal_6733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6498 ( .a ({signal_9241, signal_5849}), .b ({signal_9906, signal_6554}), .c ({signal_10097, signal_6734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6499 ( .a ({signal_9498, signal_6178}), .b ({signal_9906, signal_6554}), .c ({signal_10098, signal_6735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6500 ( .a ({signal_9498, signal_6178}), .b ({signal_9908, signal_6556}), .c ({signal_10099, signal_6736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6501 ( .a ({signal_9720, signal_6384}), .b ({signal_9909, signal_6557}), .c ({signal_10100, signal_6737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6502 ( .a ({signal_9907, signal_6555}), .b ({signal_9910, signal_6558}), .c ({signal_10101, signal_6738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6503 ( .a ({signal_9908, signal_6556}), .b ({signal_9909, signal_6557}), .c ({signal_10102, signal_6739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6504 ( .a ({signal_9499, signal_6179}), .b ({signal_9910, signal_6558}), .c ({signal_10103, signal_6740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6505 ( .a ({signal_9719, signal_6383}), .b ({signal_9911, signal_6559}), .c ({signal_10104, signal_6741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6506 ( .a ({signal_9721, signal_6385}), .b ({signal_9911, signal_6559}), .c ({signal_10105, signal_6742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6507 ( .a ({signal_9907, signal_6555}), .b ({signal_9914, signal_6562}), .c ({signal_10106, signal_6743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6508 ( .a ({signal_9591, signal_6303}), .b ({signal_9752, signal_6460}), .c ({signal_10014, signal_6744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6509 ( .a ({signal_9752, signal_6460}), .b ({signal_9840, signal_6566}), .c ({signal_10015, signal_6745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6510 ( .a ({signal_9585, signal_6297}), .b ({signal_9838, signal_6564}), .c ({signal_10016, signal_6746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6511 ( .a ({signal_9587, signal_6299}), .b ({signal_9751, signal_6459}), .c ({signal_10017, signal_6747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6512 ( .a ({signal_9751, signal_6459}), .b ({signal_9839, signal_6565}), .c ({signal_10018, signal_6748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6513 ( .a ({signal_9352, signal_6076}), .b ({signal_9837, signal_6563}), .c ({signal_10019, signal_6749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6514 ( .a ({signal_9592, signal_6304}), .b ({signal_9839, signal_6565}), .c ({signal_10020, signal_6750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6515 ( .a ({signal_9660, signal_6390}), .b ({signal_9838, signal_6564}), .c ({signal_10021, signal_6751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6516 ( .a ({signal_9837, signal_6563}), .b ({signal_9844, signal_6570}), .c ({signal_10022, signal_6752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6517 ( .a ({signal_9599, signal_6311}), .b ({signal_9754, signal_6462}), .c ({signal_10023, signal_6753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6518 ( .a ({signal_9754, signal_6462}), .b ({signal_9848, signal_6574}), .c ({signal_10024, signal_6754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6519 ( .a ({signal_9593, signal_6305}), .b ({signal_9846, signal_6572}), .c ({signal_10025, signal_6755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6520 ( .a ({signal_9595, signal_6307}), .b ({signal_9753, signal_6461}), .c ({signal_10026, signal_6756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6521 ( .a ({signal_9753, signal_6461}), .b ({signal_9847, signal_6573}), .c ({signal_10027, signal_6757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6522 ( .a ({signal_9360, signal_6084}), .b ({signal_9845, signal_6571}), .c ({signal_10028, signal_6758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6523 ( .a ({signal_9600, signal_6312}), .b ({signal_9847, signal_6573}), .c ({signal_10029, signal_6759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6524 ( .a ({signal_9664, signal_6394}), .b ({signal_9846, signal_6572}), .c ({signal_10030, signal_6760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6525 ( .a ({signal_9845, signal_6571}), .b ({signal_9852, signal_6578}), .c ({signal_10031, signal_6761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6526 ( .a ({signal_9607, signal_6319}), .b ({signal_9756, signal_6464}), .c ({signal_10032, signal_6762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6527 ( .a ({signal_9756, signal_6464}), .b ({signal_9856, signal_6582}), .c ({signal_10033, signal_6763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6528 ( .a ({signal_9601, signal_6313}), .b ({signal_9854, signal_6580}), .c ({signal_10034, signal_6764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6529 ( .a ({signal_9603, signal_6315}), .b ({signal_9755, signal_6463}), .c ({signal_10035, signal_6765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6530 ( .a ({signal_9755, signal_6463}), .b ({signal_9855, signal_6581}), .c ({signal_10036, signal_6766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6531 ( .a ({signal_9368, signal_6092}), .b ({signal_9853, signal_6579}), .c ({signal_10037, signal_6767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6532 ( .a ({signal_9608, signal_6320}), .b ({signal_9855, signal_6581}), .c ({signal_10038, signal_6768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6533 ( .a ({signal_9668, signal_6398}), .b ({signal_9854, signal_6580}), .c ({signal_10039, signal_6769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6534 ( .a ({signal_9853, signal_6579}), .b ({signal_9860, signal_6586}), .c ({signal_10040, signal_6770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6535 ( .a ({signal_9247, signal_5855}), .b ({signal_9915, signal_6587}), .c ({signal_10107, signal_6771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6536 ( .a ({signal_9249, signal_5857}), .b ({signal_9915, signal_6587}), .c ({signal_10108, signal_6772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6537 ( .a ({signal_9502, signal_6194}), .b ({signal_9915, signal_6587}), .c ({signal_10109, signal_6773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6538 ( .a ({signal_9502, signal_6194}), .b ({signal_9917, signal_6589}), .c ({signal_10110, signal_6774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6539 ( .a ({signal_9728, signal_6404}), .b ({signal_9918, signal_6590}), .c ({signal_10111, signal_6775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6540 ( .a ({signal_9916, signal_6588}), .b ({signal_9919, signal_6591}), .c ({signal_10112, signal_6776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6541 ( .a ({signal_9917, signal_6589}), .b ({signal_9918, signal_6590}), .c ({signal_10113, signal_6777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6542 ( .a ({signal_9503, signal_6195}), .b ({signal_9919, signal_6591}), .c ({signal_10114, signal_6778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6543 ( .a ({signal_9727, signal_6403}), .b ({signal_9920, signal_6592}), .c ({signal_10115, signal_6779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6544 ( .a ({signal_9729, signal_6405}), .b ({signal_9920, signal_6592}), .c ({signal_10116, signal_6780}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6545 ( .a ({signal_9916, signal_6588}), .b ({signal_9923, signal_6595}), .c ({signal_10117, signal_6781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6546 ( .a ({signal_9131, signal_5863}), .b ({signal_9861, signal_6596}), .c ({signal_10041, signal_6782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6547 ( .a ({signal_9133, signal_5865}), .b ({signal_9861, signal_6596}), .c ({signal_10042, signal_6783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6548 ( .a ({signal_9454, signal_6198}), .b ({signal_9861, signal_6596}), .c ({signal_10043, signal_6784}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6549 ( .a ({signal_9454, signal_6198}), .b ({signal_9863, signal_6598}), .c ({signal_10044, signal_6785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6550 ( .a ({signal_9674, signal_6412}), .b ({signal_9864, signal_6599}), .c ({signal_10045, signal_6786}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6551 ( .a ({signal_9862, signal_6597}), .b ({signal_9865, signal_6600}), .c ({signal_10046, signal_6787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6552 ( .a ({signal_9863, signal_6598}), .b ({signal_9864, signal_6599}), .c ({signal_10047, signal_6788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6553 ( .a ({signal_9455, signal_6199}), .b ({signal_9865, signal_6600}), .c ({signal_10048, signal_6789}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6554 ( .a ({signal_9673, signal_6411}), .b ({signal_9866, signal_6601}), .c ({signal_10049, signal_6790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6555 ( .a ({signal_9675, signal_6413}), .b ({signal_9866, signal_6601}), .c ({signal_10050, signal_6791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6556 ( .a ({signal_9862, signal_6597}), .b ({signal_9869, signal_6604}), .c ({signal_10051, signal_6792}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6557 ( .a ({signal_9139, signal_5871}), .b ({signal_9870, signal_6605}), .c ({signal_10052, signal_6793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6558 ( .a ({signal_9141, signal_5873}), .b ({signal_9870, signal_6605}), .c ({signal_10053, signal_6794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6559 ( .a ({signal_9458, signal_6202}), .b ({signal_9870, signal_6605}), .c ({signal_10054, signal_6795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6560 ( .a ({signal_9458, signal_6202}), .b ({signal_9872, signal_6607}), .c ({signal_10055, signal_6796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6561 ( .a ({signal_9682, signal_6420}), .b ({signal_9873, signal_6608}), .c ({signal_10056, signal_6797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6562 ( .a ({signal_9871, signal_6606}), .b ({signal_9874, signal_6609}), .c ({signal_10057, signal_6798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6563 ( .a ({signal_9872, signal_6607}), .b ({signal_9873, signal_6608}), .c ({signal_10058, signal_6799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6564 ( .a ({signal_9459, signal_6203}), .b ({signal_9874, signal_6609}), .c ({signal_10059, signal_6800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6565 ( .a ({signal_9681, signal_6419}), .b ({signal_9875, signal_6610}), .c ({signal_10060, signal_6801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6566 ( .a ({signal_9683, signal_6421}), .b ({signal_9875, signal_6610}), .c ({signal_10061, signal_6802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6567 ( .a ({signal_9871, signal_6606}), .b ({signal_9878, signal_6613}), .c ({signal_10062, signal_6803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6568 ( .a ({signal_9147, signal_5879}), .b ({signal_9879, signal_6614}), .c ({signal_10063, signal_6804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6569 ( .a ({signal_9149, signal_5881}), .b ({signal_9879, signal_6614}), .c ({signal_10064, signal_6805}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6570 ( .a ({signal_9462, signal_6206}), .b ({signal_9879, signal_6614}), .c ({signal_10065, signal_6806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6571 ( .a ({signal_9462, signal_6206}), .b ({signal_9881, signal_6616}), .c ({signal_10066, signal_6807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6572 ( .a ({signal_9690, signal_6428}), .b ({signal_9882, signal_6617}), .c ({signal_10067, signal_6808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6573 ( .a ({signal_9880, signal_6615}), .b ({signal_9883, signal_6618}), .c ({signal_10068, signal_6809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6574 ( .a ({signal_9881, signal_6616}), .b ({signal_9882, signal_6617}), .c ({signal_10069, signal_6810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6575 ( .a ({signal_9463, signal_6207}), .b ({signal_9883, signal_6618}), .c ({signal_10070, signal_6811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6576 ( .a ({signal_9689, signal_6427}), .b ({signal_9884, signal_6619}), .c ({signal_10071, signal_6812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6577 ( .a ({signal_9691, signal_6429}), .b ({signal_9884, signal_6619}), .c ({signal_10072, signal_6813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6578 ( .a ({signal_9880, signal_6615}), .b ({signal_9887, signal_6622}), .c ({signal_10073, signal_6814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6579 ( .a ({signal_9155, signal_5887}), .b ({signal_9888, signal_6623}), .c ({signal_10074, signal_6815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6580 ( .a ({signal_9157, signal_5889}), .b ({signal_9888, signal_6623}), .c ({signal_10075, signal_6816}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6581 ( .a ({signal_9466, signal_6210}), .b ({signal_9888, signal_6623}), .c ({signal_10076, signal_6817}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6582 ( .a ({signal_9466, signal_6210}), .b ({signal_9890, signal_6625}), .c ({signal_10077, signal_6818}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6583 ( .a ({signal_9698, signal_6436}), .b ({signal_9891, signal_6626}), .c ({signal_10078, signal_6819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6584 ( .a ({signal_9889, signal_6624}), .b ({signal_9892, signal_6627}), .c ({signal_10079, signal_6820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6585 ( .a ({signal_9890, signal_6625}), .b ({signal_9891, signal_6626}), .c ({signal_10080, signal_6821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6586 ( .a ({signal_9467, signal_6211}), .b ({signal_9892, signal_6627}), .c ({signal_10081, signal_6822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6587 ( .a ({signal_9697, signal_6435}), .b ({signal_9893, signal_6628}), .c ({signal_10082, signal_6823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6588 ( .a ({signal_9699, signal_6437}), .b ({signal_9893, signal_6628}), .c ({signal_10083, signal_6824}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6589 ( .a ({signal_9889, signal_6624}), .b ({signal_9896, signal_6631}), .c ({signal_10084, signal_6825}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6590 ( .a ({signal_10095, signal_6705}), .b ({signal_10298, signal_3938}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6591 ( .a ({signal_10106, signal_6743}), .b ({signal_10299, signal_3906}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6592 ( .a ({signal_10117, signal_6781}), .b ({signal_10300, signal_3874}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6593 ( .a ({signal_10051, signal_6792}), .b ({signal_10118, signal_3109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6594 ( .a ({signal_9267, signal_5975}), .b ({signal_9924, signal_6632}), .c ({signal_10119, signal_6826}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6595 ( .a ({signal_9269, signal_5977}), .b ({signal_9924, signal_6632}), .c ({signal_10120, signal_6827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6596 ( .a ({signal_9618, signal_6332}), .b ({signal_9924, signal_6632}), .c ({signal_10121, signal_6828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6597 ( .a ({signal_9618, signal_6332}), .b ({signal_9926, signal_6634}), .c ({signal_10122, signal_6829}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6598 ( .a ({signal_9762, signal_6470}), .b ({signal_9927, signal_6635}), .c ({signal_10123, signal_6830}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6599 ( .a ({signal_9925, signal_6633}), .b ({signal_9928, signal_6636}), .c ({signal_10124, signal_6831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6600 ( .a ({signal_9926, signal_6634}), .b ({signal_9927, signal_6635}), .c ({signal_10125, signal_6832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6601 ( .a ({signal_9619, signal_6333}), .b ({signal_9928, signal_6636}), .c ({signal_10126, signal_6833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6602 ( .a ({signal_9761, signal_6469}), .b ({signal_9929, signal_6637}), .c ({signal_10127, signal_6834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6603 ( .a ({signal_9763, signal_6471}), .b ({signal_9929, signal_6637}), .c ({signal_10128, signal_6835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6604 ( .a ({signal_9925, signal_6633}), .b ({signal_9932, signal_6640}), .c ({signal_10129, signal_6836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6605 ( .a ({signal_9275, signal_5983}), .b ({signal_9933, signal_6641}), .c ({signal_10130, signal_6837}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6606 ( .a ({signal_9277, signal_5985}), .b ({signal_9933, signal_6641}), .c ({signal_10131, signal_6838}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6607 ( .a ({signal_9622, signal_6336}), .b ({signal_9933, signal_6641}), .c ({signal_10132, signal_6839}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6608 ( .a ({signal_9622, signal_6336}), .b ({signal_9935, signal_6643}), .c ({signal_10133, signal_6840}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6609 ( .a ({signal_9770, signal_6478}), .b ({signal_9936, signal_6644}), .c ({signal_10134, signal_6841}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6610 ( .a ({signal_9934, signal_6642}), .b ({signal_9937, signal_6645}), .c ({signal_10135, signal_6842}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6611 ( .a ({signal_9935, signal_6643}), .b ({signal_9936, signal_6644}), .c ({signal_10136, signal_6843}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6612 ( .a ({signal_9623, signal_6337}), .b ({signal_9937, signal_6645}), .c ({signal_10137, signal_6844}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6613 ( .a ({signal_9769, signal_6477}), .b ({signal_9938, signal_6646}), .c ({signal_10138, signal_6845}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6614 ( .a ({signal_9771, signal_6479}), .b ({signal_9938, signal_6646}), .c ({signal_10139, signal_6846}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6615 ( .a ({signal_9934, signal_6642}), .b ({signal_9941, signal_6649}), .c ({signal_10140, signal_6847}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6616 ( .a ({signal_9283, signal_5991}), .b ({signal_9942, signal_6650}), .c ({signal_10141, signal_6848}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6617 ( .a ({signal_9285, signal_5993}), .b ({signal_9942, signal_6650}), .c ({signal_10142, signal_6849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6618 ( .a ({signal_9626, signal_6340}), .b ({signal_9942, signal_6650}), .c ({signal_10143, signal_6850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6619 ( .a ({signal_9626, signal_6340}), .b ({signal_9944, signal_6652}), .c ({signal_10144, signal_6851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6620 ( .a ({signal_9778, signal_6486}), .b ({signal_9945, signal_6653}), .c ({signal_10145, signal_6852}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6621 ( .a ({signal_9943, signal_6651}), .b ({signal_9946, signal_6654}), .c ({signal_10146, signal_6853}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6622 ( .a ({signal_9944, signal_6652}), .b ({signal_9945, signal_6653}), .c ({signal_10147, signal_6854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6623 ( .a ({signal_9627, signal_6341}), .b ({signal_9946, signal_6654}), .c ({signal_10148, signal_6855}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6624 ( .a ({signal_9777, signal_6485}), .b ({signal_9947, signal_6655}), .c ({signal_10149, signal_6856}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6625 ( .a ({signal_9779, signal_6487}), .b ({signal_9947, signal_6655}), .c ({signal_10150, signal_6857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6626 ( .a ({signal_9943, signal_6651}), .b ({signal_9950, signal_6658}), .c ({signal_10151, signal_6858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6627 ( .a ({signal_9291, signal_5999}), .b ({signal_9951, signal_6659}), .c ({signal_10152, signal_6859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6628 ( .a ({signal_9293, signal_6001}), .b ({signal_9951, signal_6659}), .c ({signal_10153, signal_6860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6629 ( .a ({signal_9630, signal_6344}), .b ({signal_9951, signal_6659}), .c ({signal_10154, signal_6861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6630 ( .a ({signal_9630, signal_6344}), .b ({signal_9953, signal_6661}), .c ({signal_10155, signal_6862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6631 ( .a ({signal_9786, signal_6494}), .b ({signal_9954, signal_6662}), .c ({signal_10156, signal_6863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6632 ( .a ({signal_9952, signal_6660}), .b ({signal_9955, signal_6663}), .c ({signal_10157, signal_6864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6633 ( .a ({signal_9953, signal_6661}), .b ({signal_9954, signal_6662}), .c ({signal_10158, signal_6865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6634 ( .a ({signal_9631, signal_6345}), .b ({signal_9955, signal_6663}), .c ({signal_10159, signal_6866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6635 ( .a ({signal_9785, signal_6493}), .b ({signal_9956, signal_6664}), .c ({signal_10160, signal_6867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6636 ( .a ({signal_9787, signal_6495}), .b ({signal_9956, signal_6664}), .c ({signal_10161, signal_6868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6637 ( .a ({signal_9952, signal_6660}), .b ({signal_9959, signal_6667}), .c ({signal_10162, signal_6869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6638 ( .a ({signal_9299, signal_6007}), .b ({signal_9960, signal_6668}), .c ({signal_10163, signal_6870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6639 ( .a ({signal_9301, signal_6009}), .b ({signal_9960, signal_6668}), .c ({signal_10164, signal_6871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6640 ( .a ({signal_9634, signal_6348}), .b ({signal_9960, signal_6668}), .c ({signal_10165, signal_6872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6641 ( .a ({signal_9634, signal_6348}), .b ({signal_9962, signal_6670}), .c ({signal_10166, signal_6873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6642 ( .a ({signal_9794, signal_6502}), .b ({signal_9963, signal_6671}), .c ({signal_10167, signal_6874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6643 ( .a ({signal_9961, signal_6669}), .b ({signal_9964, signal_6672}), .c ({signal_10168, signal_6875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6644 ( .a ({signal_9962, signal_6670}), .b ({signal_9963, signal_6671}), .c ({signal_10169, signal_6876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6645 ( .a ({signal_9635, signal_6349}), .b ({signal_9964, signal_6672}), .c ({signal_10170, signal_6877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6646 ( .a ({signal_9793, signal_6501}), .b ({signal_9965, signal_6673}), .c ({signal_10171, signal_6878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6647 ( .a ({signal_9795, signal_6503}), .b ({signal_9965, signal_6673}), .c ({signal_10172, signal_6879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6648 ( .a ({signal_9961, signal_6669}), .b ({signal_9968, signal_6676}), .c ({signal_10173, signal_6880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6649 ( .a ({signal_9307, signal_6015}), .b ({signal_9969, signal_6677}), .c ({signal_10174, signal_6881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6650 ( .a ({signal_9309, signal_6017}), .b ({signal_9969, signal_6677}), .c ({signal_10175, signal_6882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6651 ( .a ({signal_9638, signal_6352}), .b ({signal_9969, signal_6677}), .c ({signal_10176, signal_6883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6652 ( .a ({signal_9638, signal_6352}), .b ({signal_9971, signal_6679}), .c ({signal_10177, signal_6884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6653 ( .a ({signal_9802, signal_6510}), .b ({signal_9972, signal_6680}), .c ({signal_10178, signal_6885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6654 ( .a ({signal_9970, signal_6678}), .b ({signal_9973, signal_6681}), .c ({signal_10179, signal_6886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6655 ( .a ({signal_9971, signal_6679}), .b ({signal_9972, signal_6680}), .c ({signal_10180, signal_6887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6656 ( .a ({signal_9639, signal_6353}), .b ({signal_9973, signal_6681}), .c ({signal_10181, signal_6888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6657 ( .a ({signal_9801, signal_6509}), .b ({signal_9974, signal_6682}), .c ({signal_10182, signal_6889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6658 ( .a ({signal_9803, signal_6511}), .b ({signal_9974, signal_6682}), .c ({signal_10183, signal_6890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6659 ( .a ({signal_9970, signal_6678}), .b ({signal_9977, signal_6685}), .c ({signal_10184, signal_6891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6660 ( .a ({signal_9315, signal_6023}), .b ({signal_9978, signal_6686}), .c ({signal_10185, signal_6892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6661 ( .a ({signal_9317, signal_6025}), .b ({signal_9978, signal_6686}), .c ({signal_10186, signal_6893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6662 ( .a ({signal_9642, signal_6356}), .b ({signal_9978, signal_6686}), .c ({signal_10187, signal_6894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6663 ( .a ({signal_9642, signal_6356}), .b ({signal_9980, signal_6688}), .c ({signal_10188, signal_6895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6664 ( .a ({signal_9810, signal_6518}), .b ({signal_9981, signal_6689}), .c ({signal_10189, signal_6896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6665 ( .a ({signal_9979, signal_6687}), .b ({signal_9982, signal_6690}), .c ({signal_10190, signal_6897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6666 ( .a ({signal_9980, signal_6688}), .b ({signal_9981, signal_6689}), .c ({signal_10191, signal_6898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6667 ( .a ({signal_9643, signal_6357}), .b ({signal_9982, signal_6690}), .c ({signal_10192, signal_6899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6668 ( .a ({signal_9809, signal_6517}), .b ({signal_9983, signal_6691}), .c ({signal_10193, signal_6900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6669 ( .a ({signal_9811, signal_6519}), .b ({signal_9983, signal_6691}), .c ({signal_10194, signal_6901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6670 ( .a ({signal_9979, signal_6687}), .b ({signal_9986, signal_6694}), .c ({signal_10195, signal_6902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6671 ( .a ({signal_9898, signal_6522}), .b ({signal_10089, signal_6699}), .c ({signal_10301, signal_4460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6672 ( .a ({signal_10086, signal_6696}), .b ({signal_10091, signal_6701}), .c ({signal_10302, signal_6903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6673 ( .a ({signal_9903, signal_6527}), .b ({signal_10093, signal_6703}), .c ({signal_10303, signal_6904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6674 ( .a ({signal_9898, signal_6522}), .b ({signal_10088, signal_6698}), .c ({signal_10304, signal_4455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6675 ( .a ({signal_9904, signal_6528}), .b ({signal_10087, signal_6697}), .c ({signal_10305, signal_3935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6676 ( .a ({signal_10090, signal_6700}), .b ({signal_10094, signal_6704}), .c ({signal_10306, signal_3936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6677 ( .a ({signal_10085, signal_6695}), .b ({signal_10092, signal_6702}), .c ({signal_10307, signal_6905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6678 ( .a ({signal_9323, signal_6039}), .b ({signal_9987, signal_6706}), .c ({signal_10196, signal_6906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6679 ( .a ({signal_9325, signal_6041}), .b ({signal_9987, signal_6706}), .c ({signal_10197, signal_6907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6680 ( .a ({signal_9646, signal_6368}), .b ({signal_9987, signal_6706}), .c ({signal_10198, signal_6908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6681 ( .a ({signal_9646, signal_6368}), .b ({signal_9989, signal_6708}), .c ({signal_10199, signal_6909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6682 ( .a ({signal_9818, signal_6535}), .b ({signal_9990, signal_6709}), .c ({signal_10200, signal_6910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6683 ( .a ({signal_9988, signal_6707}), .b ({signal_9991, signal_6710}), .c ({signal_10201, signal_6911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6684 ( .a ({signal_9989, signal_6708}), .b ({signal_9990, signal_6709}), .c ({signal_10202, signal_6912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6685 ( .a ({signal_9647, signal_6369}), .b ({signal_9991, signal_6710}), .c ({signal_10203, signal_6913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6686 ( .a ({signal_9817, signal_6534}), .b ({signal_9992, signal_6711}), .c ({signal_10204, signal_6914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6687 ( .a ({signal_9819, signal_6536}), .b ({signal_9992, signal_6711}), .c ({signal_10205, signal_6915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6688 ( .a ({signal_9988, signal_6707}), .b ({signal_9995, signal_6714}), .c ({signal_10206, signal_6916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6689 ( .a ({signal_9331, signal_6047}), .b ({signal_9996, signal_6715}), .c ({signal_10207, signal_6917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6690 ( .a ({signal_9333, signal_6049}), .b ({signal_9996, signal_6715}), .c ({signal_10208, signal_6918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6691 ( .a ({signal_9650, signal_6372}), .b ({signal_9996, signal_6715}), .c ({signal_10209, signal_6919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6692 ( .a ({signal_9650, signal_6372}), .b ({signal_9998, signal_6717}), .c ({signal_10210, signal_6920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6693 ( .a ({signal_9826, signal_6543}), .b ({signal_9999, signal_6718}), .c ({signal_10211, signal_6921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6694 ( .a ({signal_9997, signal_6716}), .b ({signal_10000, signal_6719}), .c ({signal_10212, signal_6922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6695 ( .a ({signal_9998, signal_6717}), .b ({signal_9999, signal_6718}), .c ({signal_10213, signal_6923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6696 ( .a ({signal_9651, signal_6373}), .b ({signal_10000, signal_6719}), .c ({signal_10214, signal_6924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6697 ( .a ({signal_9825, signal_6542}), .b ({signal_10001, signal_6720}), .c ({signal_10215, signal_6925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6698 ( .a ({signal_9827, signal_6544}), .b ({signal_10001, signal_6720}), .c ({signal_10216, signal_6926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6699 ( .a ({signal_9997, signal_6716}), .b ({signal_10004, signal_6723}), .c ({signal_10217, signal_6927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6700 ( .a ({signal_9339, signal_6055}), .b ({signal_10005, signal_6724}), .c ({signal_10218, signal_6928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6701 ( .a ({signal_9341, signal_6057}), .b ({signal_10005, signal_6724}), .c ({signal_10219, signal_6929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6702 ( .a ({signal_9654, signal_6376}), .b ({signal_10005, signal_6724}), .c ({signal_10220, signal_6930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6703 ( .a ({signal_9654, signal_6376}), .b ({signal_10007, signal_6726}), .c ({signal_10221, signal_6931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6704 ( .a ({signal_9834, signal_6551}), .b ({signal_10008, signal_6727}), .c ({signal_10222, signal_6932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6705 ( .a ({signal_10006, signal_6725}), .b ({signal_10009, signal_6728}), .c ({signal_10223, signal_6933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6706 ( .a ({signal_10007, signal_6726}), .b ({signal_10008, signal_6727}), .c ({signal_10224, signal_6934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6707 ( .a ({signal_9655, signal_6377}), .b ({signal_10009, signal_6728}), .c ({signal_10225, signal_6935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6708 ( .a ({signal_9833, signal_6550}), .b ({signal_10010, signal_6729}), .c ({signal_10226, signal_6936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6709 ( .a ({signal_9835, signal_6552}), .b ({signal_10010, signal_6729}), .c ({signal_10227, signal_6937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6710 ( .a ({signal_10006, signal_6725}), .b ({signal_10013, signal_6732}), .c ({signal_10228, signal_6938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6711 ( .a ({signal_9907, signal_6555}), .b ({signal_10100, signal_6737}), .c ({signal_10308, signal_4428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6712 ( .a ({signal_10097, signal_6734}), .b ({signal_10102, signal_6739}), .c ({signal_10309, signal_6939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6713 ( .a ({signal_9912, signal_6560}), .b ({signal_10104, signal_6741}), .c ({signal_10310, signal_6940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6714 ( .a ({signal_9907, signal_6555}), .b ({signal_10099, signal_6736}), .c ({signal_10311, signal_4423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6715 ( .a ({signal_9913, signal_6561}), .b ({signal_10098, signal_6735}), .c ({signal_10312, signal_3903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6716 ( .a ({signal_10101, signal_6738}), .b ({signal_10105, signal_6742}), .c ({signal_10313, signal_3904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6717 ( .a ({signal_10096, signal_6733}), .b ({signal_10103, signal_6740}), .c ({signal_10314, signal_6941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6718 ( .a ({signal_9347, signal_6071}), .b ({signal_10014, signal_6744}), .c ({signal_10229, signal_6942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6719 ( .a ({signal_9349, signal_6073}), .b ({signal_10014, signal_6744}), .c ({signal_10230, signal_6943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6720 ( .a ({signal_9658, signal_6388}), .b ({signal_10014, signal_6744}), .c ({signal_10231, signal_6944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6721 ( .a ({signal_9658, signal_6388}), .b ({signal_10016, signal_6746}), .c ({signal_10232, signal_6945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6722 ( .a ({signal_9842, signal_6568}), .b ({signal_10017, signal_6747}), .c ({signal_10233, signal_6946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6723 ( .a ({signal_10015, signal_6745}), .b ({signal_10018, signal_6748}), .c ({signal_10234, signal_6947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6724 ( .a ({signal_10016, signal_6746}), .b ({signal_10017, signal_6747}), .c ({signal_10235, signal_6948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6725 ( .a ({signal_9659, signal_6389}), .b ({signal_10018, signal_6748}), .c ({signal_10236, signal_6949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6726 ( .a ({signal_9841, signal_6567}), .b ({signal_10019, signal_6749}), .c ({signal_10237, signal_6950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6727 ( .a ({signal_9843, signal_6569}), .b ({signal_10019, signal_6749}), .c ({signal_10238, signal_6951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6728 ( .a ({signal_10015, signal_6745}), .b ({signal_10022, signal_6752}), .c ({signal_10239, signal_6952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6729 ( .a ({signal_9355, signal_6079}), .b ({signal_10023, signal_6753}), .c ({signal_10240, signal_6953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6730 ( .a ({signal_9357, signal_6081}), .b ({signal_10023, signal_6753}), .c ({signal_10241, signal_6954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6731 ( .a ({signal_9662, signal_6392}), .b ({signal_10023, signal_6753}), .c ({signal_10242, signal_6955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6732 ( .a ({signal_9662, signal_6392}), .b ({signal_10025, signal_6755}), .c ({signal_10243, signal_6956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6733 ( .a ({signal_9850, signal_6576}), .b ({signal_10026, signal_6756}), .c ({signal_10244, signal_6957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6734 ( .a ({signal_10024, signal_6754}), .b ({signal_10027, signal_6757}), .c ({signal_10245, signal_6958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6735 ( .a ({signal_10025, signal_6755}), .b ({signal_10026, signal_6756}), .c ({signal_10246, signal_6959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6736 ( .a ({signal_9663, signal_6393}), .b ({signal_10027, signal_6757}), .c ({signal_10247, signal_6960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6737 ( .a ({signal_9849, signal_6575}), .b ({signal_10028, signal_6758}), .c ({signal_10248, signal_6961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6738 ( .a ({signal_9851, signal_6577}), .b ({signal_10028, signal_6758}), .c ({signal_10249, signal_6962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6739 ( .a ({signal_10024, signal_6754}), .b ({signal_10031, signal_6761}), .c ({signal_10250, signal_6963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6740 ( .a ({signal_9363, signal_6087}), .b ({signal_10032, signal_6762}), .c ({signal_10251, signal_6964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6741 ( .a ({signal_9365, signal_6089}), .b ({signal_10032, signal_6762}), .c ({signal_10252, signal_6965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6742 ( .a ({signal_9666, signal_6396}), .b ({signal_10032, signal_6762}), .c ({signal_10253, signal_6966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6743 ( .a ({signal_9666, signal_6396}), .b ({signal_10034, signal_6764}), .c ({signal_10254, signal_6967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6744 ( .a ({signal_9858, signal_6584}), .b ({signal_10035, signal_6765}), .c ({signal_10255, signal_6968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6745 ( .a ({signal_10033, signal_6763}), .b ({signal_10036, signal_6766}), .c ({signal_10256, signal_6969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6746 ( .a ({signal_10034, signal_6764}), .b ({signal_10035, signal_6765}), .c ({signal_10257, signal_6970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6747 ( .a ({signal_9667, signal_6397}), .b ({signal_10036, signal_6766}), .c ({signal_10258, signal_6971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6748 ( .a ({signal_9857, signal_6583}), .b ({signal_10037, signal_6767}), .c ({signal_10259, signal_6972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6749 ( .a ({signal_9859, signal_6585}), .b ({signal_10037, signal_6767}), .c ({signal_10260, signal_6973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6750 ( .a ({signal_10033, signal_6763}), .b ({signal_10040, signal_6770}), .c ({signal_10261, signal_6974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6751 ( .a ({signal_9916, signal_6588}), .b ({signal_10111, signal_6775}), .c ({signal_10315, signal_4396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6752 ( .a ({signal_10108, signal_6772}), .b ({signal_10113, signal_6777}), .c ({signal_10316, signal_6975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6753 ( .a ({signal_9921, signal_6593}), .b ({signal_10115, signal_6779}), .c ({signal_10317, signal_6976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6754 ( .a ({signal_9916, signal_6588}), .b ({signal_10110, signal_6774}), .c ({signal_10318, signal_4391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6755 ( .a ({signal_9922, signal_6594}), .b ({signal_10109, signal_6773}), .c ({signal_10319, signal_3871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6756 ( .a ({signal_10112, signal_6776}), .b ({signal_10116, signal_6780}), .c ({signal_10320, signal_3872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6757 ( .a ({signal_10107, signal_6771}), .b ({signal_10114, signal_6778}), .c ({signal_10321, signal_6977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6758 ( .a ({signal_22488, signal_22480}), .b ({signal_10062, signal_6803}), .c ({signal_10262, signal_6978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6759 ( .a ({signal_22504, signal_22496}), .b ({signal_10073, signal_6814}), .c ({signal_10263, signal_6979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6760 ( .a ({signal_22520, signal_22512}), .b ({signal_10084, signal_6825}), .c ({signal_10264, signal_6980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6761 ( .a ({signal_9862, signal_6597}), .b ({signal_10045, signal_6786}), .c ({signal_10265, signal_3116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6762 ( .a ({signal_10042, signal_6783}), .b ({signal_10047, signal_6788}), .c ({signal_10266, signal_6981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6763 ( .a ({signal_9867, signal_6602}), .b ({signal_10049, signal_6790}), .c ({signal_10267, signal_6982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6764 ( .a ({signal_9862, signal_6597}), .b ({signal_10044, signal_6785}), .c ({signal_10268, signal_3113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6765 ( .a ({signal_9868, signal_6603}), .b ({signal_10043, signal_6784}), .c ({signal_10269, signal_3112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6766 ( .a ({signal_10046, signal_6787}), .b ({signal_10050, signal_6791}), .c ({signal_10270, signal_3111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6767 ( .a ({signal_10041, signal_6782}), .b ({signal_10048, signal_6789}), .c ({signal_10271, signal_6983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6768 ( .a ({signal_9871, signal_6606}), .b ({signal_10056, signal_6797}), .c ({signal_10272, signal_6984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6769 ( .a ({signal_10053, signal_6794}), .b ({signal_10058, signal_6799}), .c ({signal_10273, signal_6985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6770 ( .a ({signal_9876, signal_6611}), .b ({signal_10060, signal_6801}), .c ({signal_10274, signal_6986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6771 ( .a ({signal_9871, signal_6606}), .b ({signal_10055, signal_6796}), .c ({signal_10275, signal_6987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6772 ( .a ({signal_9877, signal_6612}), .b ({signal_10054, signal_6795}), .c ({signal_10276, signal_6988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6773 ( .a ({signal_10057, signal_6798}), .b ({signal_10061, signal_6802}), .c ({signal_10277, signal_6989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6774 ( .a ({signal_10052, signal_6793}), .b ({signal_10059, signal_6800}), .c ({signal_10278, signal_6990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6775 ( .a ({signal_9880, signal_6615}), .b ({signal_10067, signal_6808}), .c ({signal_10279, signal_6991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6776 ( .a ({signal_10064, signal_6805}), .b ({signal_10069, signal_6810}), .c ({signal_10280, signal_6992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6777 ( .a ({signal_9885, signal_6620}), .b ({signal_10071, signal_6812}), .c ({signal_10281, signal_6993}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6778 ( .a ({signal_9880, signal_6615}), .b ({signal_10066, signal_6807}), .c ({signal_10282, signal_6994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6779 ( .a ({signal_9886, signal_6621}), .b ({signal_10065, signal_6806}), .c ({signal_10283, signal_6995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6780 ( .a ({signal_10068, signal_6809}), .b ({signal_10072, signal_6813}), .c ({signal_10284, signal_6996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6781 ( .a ({signal_10063, signal_6804}), .b ({signal_10070, signal_6811}), .c ({signal_10285, signal_6997}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6782 ( .a ({signal_9889, signal_6624}), .b ({signal_10078, signal_6819}), .c ({signal_10286, signal_6998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6783 ( .a ({signal_10075, signal_6816}), .b ({signal_10080, signal_6821}), .c ({signal_10287, signal_6999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6784 ( .a ({signal_9894, signal_6629}), .b ({signal_10082, signal_6823}), .c ({signal_10288, signal_7000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6785 ( .a ({signal_9889, signal_6624}), .b ({signal_10077, signal_6818}), .c ({signal_10289, signal_7001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6786 ( .a ({signal_9895, signal_6630}), .b ({signal_10076, signal_6817}), .c ({signal_10290, signal_7002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6787 ( .a ({signal_10079, signal_6820}), .b ({signal_10083, signal_6824}), .c ({signal_10291, signal_7003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6788 ( .a ({signal_10074, signal_6815}), .b ({signal_10081, signal_6822}), .c ({signal_10292, signal_7004}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6789 ( .a ({signal_10129, signal_6836}), .b ({signal_10322, signal_3898}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6790 ( .a ({signal_10140, signal_6847}), .b ({signal_10323, signal_3922}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6791 ( .a ({signal_10151, signal_6858}), .b ({signal_10324, signal_3946}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6792 ( .a ({signal_10162, signal_6869}), .b ({signal_10325, signal_3970}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6793 ( .a ({signal_10173, signal_6880}), .b ({signal_10326, signal_3994}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6794 ( .a ({signal_10184, signal_6891}), .b ({signal_10327, signal_3890}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6795 ( .a ({signal_10195, signal_6902}), .b ({signal_10328, signal_3914}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6796 ( .a ({signal_10302, signal_6903}), .b ({signal_10494, signal_4453}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6797 ( .a ({signal_10303, signal_6904}), .b ({signal_10495, signal_4454}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6798 ( .a ({signal_10307, signal_6905}), .b ({signal_10496, signal_4458}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6799 ( .a ({signal_10206, signal_6916}), .b ({signal_10329, signal_3962}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6800 ( .a ({signal_10217, signal_6927}), .b ({signal_10330, signal_3986}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6801 ( .a ({signal_10228, signal_6938}), .b ({signal_10331, signal_3882}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6802 ( .a ({signal_10309, signal_6939}), .b ({signal_10497, signal_4421}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6803 ( .a ({signal_10310, signal_6940}), .b ({signal_10498, signal_4422}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6804 ( .a ({signal_10314, signal_6941}), .b ({signal_10499, signal_4426}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6805 ( .a ({signal_10239, signal_6952}), .b ({signal_10332, signal_3930}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6806 ( .a ({signal_10250, signal_6963}), .b ({signal_10333, signal_3954}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6807 ( .a ({signal_10261, signal_6974}), .b ({signal_10334, signal_3978}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6808 ( .a ({signal_10316, signal_6975}), .b ({signal_10500, signal_4389}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6809 ( .a ({signal_10317, signal_6976}), .b ({signal_10501, signal_4390}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6810 ( .a ({signal_10321, signal_6977}), .b ({signal_10502, signal_4394}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6811 ( .a ({signal_10262, signal_6978}), .b ({signal_10335, signal_4138}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6812 ( .a ({signal_10263, signal_6979}), .b ({signal_10336, signal_4146}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6813 ( .a ({signal_10264, signal_6980}), .b ({signal_10337, signal_4154}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6814 ( .a ({signal_10266, signal_6981}), .b ({signal_10338, signal_3115}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6815 ( .a ({signal_10267, signal_6982}), .b ({signal_10339, signal_3114}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6816 ( .a ({signal_10271, signal_6983}), .b ({signal_10340, signal_3110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6817 ( .a ({signal_9925, signal_6633}), .b ({signal_10123, signal_6830}), .c ({signal_10341, signal_4420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6818 ( .a ({signal_10120, signal_6827}), .b ({signal_10125, signal_6832}), .c ({signal_10342, signal_7005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6819 ( .a ({signal_9930, signal_6638}), .b ({signal_10127, signal_6834}), .c ({signal_10343, signal_7006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6820 ( .a ({signal_9925, signal_6633}), .b ({signal_10122, signal_6829}), .c ({signal_10344, signal_4415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6821 ( .a ({signal_9931, signal_6639}), .b ({signal_10121, signal_6828}), .c ({signal_10345, signal_3895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6822 ( .a ({signal_10124, signal_6831}), .b ({signal_10128, signal_6835}), .c ({signal_10346, signal_3896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6823 ( .a ({signal_10119, signal_6826}), .b ({signal_10126, signal_6833}), .c ({signal_10347, signal_7007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6824 ( .a ({signal_9934, signal_6642}), .b ({signal_10134, signal_6841}), .c ({signal_10348, signal_4444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6825 ( .a ({signal_10131, signal_6838}), .b ({signal_10136, signal_6843}), .c ({signal_10349, signal_7008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6826 ( .a ({signal_9939, signal_6647}), .b ({signal_10138, signal_6845}), .c ({signal_10350, signal_7009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6827 ( .a ({signal_9934, signal_6642}), .b ({signal_10133, signal_6840}), .c ({signal_10351, signal_4439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6828 ( .a ({signal_9940, signal_6648}), .b ({signal_10132, signal_6839}), .c ({signal_10352, signal_3919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6829 ( .a ({signal_10135, signal_6842}), .b ({signal_10139, signal_6846}), .c ({signal_10353, signal_3920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6830 ( .a ({signal_10130, signal_6837}), .b ({signal_10137, signal_6844}), .c ({signal_10354, signal_7010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6831 ( .a ({signal_9943, signal_6651}), .b ({signal_10145, signal_6852}), .c ({signal_10355, signal_4468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6832 ( .a ({signal_10142, signal_6849}), .b ({signal_10147, signal_6854}), .c ({signal_10356, signal_7011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6833 ( .a ({signal_9948, signal_6656}), .b ({signal_10149, signal_6856}), .c ({signal_10357, signal_7012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6834 ( .a ({signal_9943, signal_6651}), .b ({signal_10144, signal_6851}), .c ({signal_10358, signal_4463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6835 ( .a ({signal_9949, signal_6657}), .b ({signal_10143, signal_6850}), .c ({signal_10359, signal_3943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6836 ( .a ({signal_10146, signal_6853}), .b ({signal_10150, signal_6857}), .c ({signal_10360, signal_3944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6837 ( .a ({signal_10141, signal_6848}), .b ({signal_10148, signal_6855}), .c ({signal_10361, signal_7013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6838 ( .a ({signal_9952, signal_6660}), .b ({signal_10156, signal_6863}), .c ({signal_10362, signal_4492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6839 ( .a ({signal_10153, signal_6860}), .b ({signal_10158, signal_6865}), .c ({signal_10363, signal_7014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6840 ( .a ({signal_9957, signal_6665}), .b ({signal_10160, signal_6867}), .c ({signal_10364, signal_7015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6841 ( .a ({signal_9952, signal_6660}), .b ({signal_10155, signal_6862}), .c ({signal_10365, signal_4487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6842 ( .a ({signal_9958, signal_6666}), .b ({signal_10154, signal_6861}), .c ({signal_10366, signal_3967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6843 ( .a ({signal_10157, signal_6864}), .b ({signal_10161, signal_6868}), .c ({signal_10367, signal_3968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6844 ( .a ({signal_10152, signal_6859}), .b ({signal_10159, signal_6866}), .c ({signal_10368, signal_7016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6845 ( .a ({signal_9961, signal_6669}), .b ({signal_10167, signal_6874}), .c ({signal_10369, signal_4516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6846 ( .a ({signal_10164, signal_6871}), .b ({signal_10169, signal_6876}), .c ({signal_10370, signal_7017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6847 ( .a ({signal_9966, signal_6674}), .b ({signal_10171, signal_6878}), .c ({signal_10371, signal_7018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6848 ( .a ({signal_9961, signal_6669}), .b ({signal_10166, signal_6873}), .c ({signal_10372, signal_4511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6849 ( .a ({signal_9967, signal_6675}), .b ({signal_10165, signal_6872}), .c ({signal_10373, signal_3991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6850 ( .a ({signal_10168, signal_6875}), .b ({signal_10172, signal_6879}), .c ({signal_10374, signal_3992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6851 ( .a ({signal_10163, signal_6870}), .b ({signal_10170, signal_6877}), .c ({signal_10375, signal_7019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6852 ( .a ({signal_9970, signal_6678}), .b ({signal_10178, signal_6885}), .c ({signal_10376, signal_4412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6853 ( .a ({signal_10175, signal_6882}), .b ({signal_10180, signal_6887}), .c ({signal_10377, signal_7020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6854 ( .a ({signal_9975, signal_6683}), .b ({signal_10182, signal_6889}), .c ({signal_10378, signal_7021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6855 ( .a ({signal_9970, signal_6678}), .b ({signal_10177, signal_6884}), .c ({signal_10379, signal_4407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6856 ( .a ({signal_9976, signal_6684}), .b ({signal_10176, signal_6883}), .c ({signal_10380, signal_3887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6857 ( .a ({signal_10179, signal_6886}), .b ({signal_10183, signal_6890}), .c ({signal_10381, signal_3888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6858 ( .a ({signal_10174, signal_6881}), .b ({signal_10181, signal_6888}), .c ({signal_10382, signal_7022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6859 ( .a ({signal_9979, signal_6687}), .b ({signal_10189, signal_6896}), .c ({signal_10383, signal_4436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6860 ( .a ({signal_10186, signal_6893}), .b ({signal_10191, signal_6898}), .c ({signal_10384, signal_7023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6861 ( .a ({signal_9984, signal_6692}), .b ({signal_10193, signal_6900}), .c ({signal_10385, signal_7024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6862 ( .a ({signal_9979, signal_6687}), .b ({signal_10188, signal_6895}), .c ({signal_10386, signal_4431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6863 ( .a ({signal_9985, signal_6693}), .b ({signal_10187, signal_6894}), .c ({signal_10387, signal_3911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6864 ( .a ({signal_10190, signal_6897}), .b ({signal_10194, signal_6901}), .c ({signal_10388, signal_3912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6865 ( .a ({signal_10185, signal_6892}), .b ({signal_10192, signal_6899}), .c ({signal_10389, signal_7025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6866 ( .a ({signal_9988, signal_6707}), .b ({signal_10200, signal_6910}), .c ({signal_10390, signal_4484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6867 ( .a ({signal_10197, signal_6907}), .b ({signal_10202, signal_6912}), .c ({signal_10391, signal_7026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6868 ( .a ({signal_9993, signal_6712}), .b ({signal_10204, signal_6914}), .c ({signal_10392, signal_7027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6869 ( .a ({signal_9988, signal_6707}), .b ({signal_10199, signal_6909}), .c ({signal_10393, signal_4479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6870 ( .a ({signal_9994, signal_6713}), .b ({signal_10198, signal_6908}), .c ({signal_10394, signal_3959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6871 ( .a ({signal_10201, signal_6911}), .b ({signal_10205, signal_6915}), .c ({signal_10395, signal_3960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6872 ( .a ({signal_10196, signal_6906}), .b ({signal_10203, signal_6913}), .c ({signal_10396, signal_7028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6873 ( .a ({signal_9997, signal_6716}), .b ({signal_10211, signal_6921}), .c ({signal_10397, signal_4508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6874 ( .a ({signal_10208, signal_6918}), .b ({signal_10213, signal_6923}), .c ({signal_10398, signal_7029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6875 ( .a ({signal_10002, signal_6721}), .b ({signal_10215, signal_6925}), .c ({signal_10399, signal_7030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6876 ( .a ({signal_9997, signal_6716}), .b ({signal_10210, signal_6920}), .c ({signal_10400, signal_4503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6877 ( .a ({signal_10003, signal_6722}), .b ({signal_10209, signal_6919}), .c ({signal_10401, signal_3983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6878 ( .a ({signal_10212, signal_6922}), .b ({signal_10216, signal_6926}), .c ({signal_10402, signal_3984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6879 ( .a ({signal_10207, signal_6917}), .b ({signal_10214, signal_6924}), .c ({signal_10403, signal_7031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6880 ( .a ({signal_10006, signal_6725}), .b ({signal_10222, signal_6932}), .c ({signal_10404, signal_4404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6881 ( .a ({signal_10219, signal_6929}), .b ({signal_10224, signal_6934}), .c ({signal_10405, signal_7032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6882 ( .a ({signal_10011, signal_6730}), .b ({signal_10226, signal_6936}), .c ({signal_10406, signal_7033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6883 ( .a ({signal_10006, signal_6725}), .b ({signal_10221, signal_6931}), .c ({signal_10407, signal_4399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6884 ( .a ({signal_10012, signal_6731}), .b ({signal_10220, signal_6930}), .c ({signal_10408, signal_3879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6885 ( .a ({signal_10223, signal_6933}), .b ({signal_10227, signal_6937}), .c ({signal_10409, signal_3880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6886 ( .a ({signal_10218, signal_6928}), .b ({signal_10225, signal_6935}), .c ({signal_10410, signal_7034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6887 ( .a ({signal_10015, signal_6745}), .b ({signal_10233, signal_6946}), .c ({signal_10411, signal_4452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6888 ( .a ({signal_10230, signal_6943}), .b ({signal_10235, signal_6948}), .c ({signal_10412, signal_7035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6889 ( .a ({signal_10020, signal_6750}), .b ({signal_10237, signal_6950}), .c ({signal_10413, signal_7036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6890 ( .a ({signal_10015, signal_6745}), .b ({signal_10232, signal_6945}), .c ({signal_10414, signal_4447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6891 ( .a ({signal_10021, signal_6751}), .b ({signal_10231, signal_6944}), .c ({signal_10415, signal_3927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6892 ( .a ({signal_10234, signal_6947}), .b ({signal_10238, signal_6951}), .c ({signal_10416, signal_3928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6893 ( .a ({signal_10229, signal_6942}), .b ({signal_10236, signal_6949}), .c ({signal_10417, signal_7037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6894 ( .a ({signal_10024, signal_6754}), .b ({signal_10244, signal_6957}), .c ({signal_10418, signal_4476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6895 ( .a ({signal_10241, signal_6954}), .b ({signal_10246, signal_6959}), .c ({signal_10419, signal_7038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6896 ( .a ({signal_10029, signal_6759}), .b ({signal_10248, signal_6961}), .c ({signal_10420, signal_7039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6897 ( .a ({signal_10024, signal_6754}), .b ({signal_10243, signal_6956}), .c ({signal_10421, signal_4471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6898 ( .a ({signal_10030, signal_6760}), .b ({signal_10242, signal_6955}), .c ({signal_10422, signal_3951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6899 ( .a ({signal_10245, signal_6958}), .b ({signal_10249, signal_6962}), .c ({signal_10423, signal_3952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6900 ( .a ({signal_10240, signal_6953}), .b ({signal_10247, signal_6960}), .c ({signal_10424, signal_7040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6901 ( .a ({signal_10033, signal_6763}), .b ({signal_10255, signal_6968}), .c ({signal_10425, signal_4500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6902 ( .a ({signal_10252, signal_6965}), .b ({signal_10257, signal_6970}), .c ({signal_10426, signal_7041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6903 ( .a ({signal_10038, signal_6768}), .b ({signal_10259, signal_6972}), .c ({signal_10427, signal_7042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6904 ( .a ({signal_10033, signal_6763}), .b ({signal_10254, signal_6967}), .c ({signal_10428, signal_4495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6905 ( .a ({signal_10039, signal_6769}), .b ({signal_10253, signal_6966}), .c ({signal_10429, signal_3975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6906 ( .a ({signal_10256, signal_6969}), .b ({signal_10260, signal_6973}), .c ({signal_10430, signal_3976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6907 ( .a ({signal_10251, signal_6964}), .b ({signal_10258, signal_6971}), .c ({signal_10431, signal_7043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6908 ( .a ({signal_10228, signal_6938}), .b ({signal_10315, signal_4396}), .c ({signal_10503, signal_7044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6909 ( .a ({signal_10315, signal_4396}), .b ({signal_10319, signal_3871}), .c ({signal_10504, signal_7045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6910 ( .a ({signal_10315, signal_4396}), .b ({signal_10320, signal_3872}), .c ({signal_10505, signal_7046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6911 ( .a ({signal_10117, signal_6781}), .b ({signal_10315, signal_4396}), .c ({signal_10506, signal_7047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6912 ( .a ({signal_10195, signal_6902}), .b ({signal_10308, signal_4428}), .c ({signal_10507, signal_7048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6913 ( .a ({signal_10308, signal_4428}), .b ({signal_10312, signal_3903}), .c ({signal_10508, signal_7049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6914 ( .a ({signal_10308, signal_4428}), .b ({signal_10313, signal_3904}), .c ({signal_10509, signal_7050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6915 ( .a ({signal_10106, signal_6743}), .b ({signal_10308, signal_4428}), .c ({signal_10510, signal_7051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6916 ( .a ({signal_10151, signal_6858}), .b ({signal_10301, signal_4460}), .c ({signal_10511, signal_7052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6917 ( .a ({signal_10301, signal_4460}), .b ({signal_10305, signal_3935}), .c ({signal_10512, signal_7053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6918 ( .a ({signal_10301, signal_4460}), .b ({signal_10306, signal_3936}), .c ({signal_10513, signal_7054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6919 ( .a ({signal_10095, signal_6705}), .b ({signal_10301, signal_4460}), .c ({signal_10514, signal_7055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6920 ( .a ({signal_22536, signal_22528}), .b ({signal_10263, signal_6979}), .c ({signal_10432, signal_7056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6921 ( .a ({signal_22552, signal_22544}), .b ({signal_10290, signal_7002}), .c ({signal_10433, signal_4151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6922 ( .a ({signal_22568, signal_22560}), .b ({signal_10291, signal_7003}), .c ({signal_10434, signal_4152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6923 ( .a ({signal_22584, signal_22576}), .b ({signal_10292, signal_7004}), .c ({signal_10435, signal_7057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6924 ( .a ({signal_22600, signal_22592}), .b ({signal_10262, signal_6978}), .c ({signal_10436, signal_7058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6925 ( .a ({signal_22616, signal_22608}), .b ({signal_10272, signal_6984}), .c ({signal_10437, signal_4131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6926 ( .a ({signal_22632, signal_22624}), .b ({signal_10273, signal_6985}), .c ({signal_10438, signal_7059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6927 ( .a ({signal_22648, signal_22640}), .b ({signal_10274, signal_6986}), .c ({signal_10439, signal_7060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6928 ( .a ({signal_22664, signal_22656}), .b ({signal_10275, signal_6987}), .c ({signal_10440, signal_4134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6929 ( .a ({signal_22680, signal_22672}), .b ({signal_10276, signal_6988}), .c ({signal_10441, signal_4135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6930 ( .a ({signal_22696, signal_22688}), .b ({signal_10277, signal_6989}), .c ({signal_10442, signal_4136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6931 ( .a ({signal_22712, signal_22704}), .b ({signal_10278, signal_6990}), .c ({signal_10443, signal_7061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6932 ( .a ({signal_22728, signal_22720}), .b ({signal_10279, signal_6991}), .c ({signal_10444, signal_4139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6933 ( .a ({signal_22744, signal_22736}), .b ({signal_10280, signal_6992}), .c ({signal_10445, signal_7062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6934 ( .a ({signal_22760, signal_22752}), .b ({signal_10281, signal_6993}), .c ({signal_10446, signal_7063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6935 ( .a ({signal_22776, signal_22768}), .b ({signal_10282, signal_6994}), .c ({signal_10447, signal_4142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6936 ( .a ({signal_22792, signal_22784}), .b ({signal_10283, signal_6995}), .c ({signal_10448, signal_4143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6937 ( .a ({signal_22808, signal_22800}), .b ({signal_10284, signal_6996}), .c ({signal_10449, signal_4144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6938 ( .a ({signal_22824, signal_22816}), .b ({signal_10285, signal_6997}), .c ({signal_10450, signal_7064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6939 ( .a ({signal_22840, signal_22832}), .b ({signal_10286, signal_6998}), .c ({signal_10451, signal_4147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6940 ( .a ({signal_22856, signal_22848}), .b ({signal_10287, signal_6999}), .c ({signal_10452, signal_7065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6941 ( .a ({signal_22872, signal_22864}), .b ({signal_10288, signal_7000}), .c ({signal_10453, signal_7066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6942 ( .a ({signal_22888, signal_22880}), .b ({signal_10289, signal_7001}), .c ({signal_10454, signal_4150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6943 ( .a ({signal_22904, signal_22896}), .b ({signal_10264, signal_6980}), .c ({signal_10455, signal_7067}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6944 ( .a ({signal_10342, signal_7005}), .b ({signal_10515, signal_4413}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6945 ( .a ({signal_10343, signal_7006}), .b ({signal_10516, signal_4414}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6946 ( .a ({signal_10347, signal_7007}), .b ({signal_10517, signal_4418}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6947 ( .a ({signal_10349, signal_7008}), .b ({signal_10518, signal_4437}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6948 ( .a ({signal_10350, signal_7009}), .b ({signal_10519, signal_4438}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6949 ( .a ({signal_10354, signal_7010}), .b ({signal_10520, signal_4442}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6950 ( .a ({signal_10356, signal_7011}), .b ({signal_10521, signal_4461}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6951 ( .a ({signal_10357, signal_7012}), .b ({signal_10522, signal_4462}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6952 ( .a ({signal_10361, signal_7013}), .b ({signal_10523, signal_4466}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6953 ( .a ({signal_10363, signal_7014}), .b ({signal_10524, signal_4485}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6954 ( .a ({signal_10364, signal_7015}), .b ({signal_10525, signal_4486}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6955 ( .a ({signal_10368, signal_7016}), .b ({signal_10526, signal_4490}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6956 ( .a ({signal_10370, signal_7017}), .b ({signal_10527, signal_4509}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6957 ( .a ({signal_10371, signal_7018}), .b ({signal_10528, signal_4510}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6958 ( .a ({signal_10375, signal_7019}), .b ({signal_10529, signal_4514}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6959 ( .a ({signal_10377, signal_7020}), .b ({signal_10530, signal_4405}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6960 ( .a ({signal_10378, signal_7021}), .b ({signal_10531, signal_4406}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6961 ( .a ({signal_10382, signal_7022}), .b ({signal_10532, signal_4410}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6962 ( .a ({signal_10384, signal_7023}), .b ({signal_10533, signal_4429}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6963 ( .a ({signal_10385, signal_7024}), .b ({signal_10534, signal_4430}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6964 ( .a ({signal_10389, signal_7025}), .b ({signal_10535, signal_4434}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6965 ( .a ({signal_10391, signal_7026}), .b ({signal_10536, signal_4477}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6966 ( .a ({signal_10392, signal_7027}), .b ({signal_10537, signal_4478}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6967 ( .a ({signal_10396, signal_7028}), .b ({signal_10538, signal_4482}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6968 ( .a ({signal_10398, signal_7029}), .b ({signal_10539, signal_4501}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6969 ( .a ({signal_10399, signal_7030}), .b ({signal_10540, signal_4502}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6970 ( .a ({signal_10403, signal_7031}), .b ({signal_10541, signal_4506}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6971 ( .a ({signal_10405, signal_7032}), .b ({signal_10542, signal_4397}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6972 ( .a ({signal_10406, signal_7033}), .b ({signal_10543, signal_4398}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6973 ( .a ({signal_10410, signal_7034}), .b ({signal_10544, signal_4402}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6974 ( .a ({signal_10412, signal_7035}), .b ({signal_10545, signal_4445}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6975 ( .a ({signal_10413, signal_7036}), .b ({signal_10546, signal_4446}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6976 ( .a ({signal_10417, signal_7037}), .b ({signal_10547, signal_4450}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6977 ( .a ({signal_10419, signal_7038}), .b ({signal_10548, signal_4469}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6978 ( .a ({signal_10420, signal_7039}), .b ({signal_10549, signal_4470}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6979 ( .a ({signal_10424, signal_7040}), .b ({signal_10550, signal_4474}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6980 ( .a ({signal_10426, signal_7041}), .b ({signal_10551, signal_4493}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6981 ( .a ({signal_10427, signal_7042}), .b ({signal_10552, signal_4494}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6982 ( .a ({signal_10431, signal_7043}), .b ({signal_10553, signal_4498}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6983 ( .a ({signal_10432, signal_7056}), .b ({signal_10554, signal_4178}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6984 ( .a ({signal_10435, signal_7057}), .b ({signal_10555, signal_4153}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6985 ( .a ({signal_10436, signal_7058}), .b ({signal_10556, signal_4170}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6986 ( .a ({signal_10438, signal_7059}), .b ({signal_10557, signal_4132}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6987 ( .a ({signal_10439, signal_7060}), .b ({signal_10558, signal_4133}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6988 ( .a ({signal_10443, signal_7061}), .b ({signal_10559, signal_4137}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6989 ( .a ({signal_10445, signal_7062}), .b ({signal_10560, signal_4140}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6990 ( .a ({signal_10446, signal_7063}), .b ({signal_10561, signal_4141}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6991 ( .a ({signal_10450, signal_7064}), .b ({signal_10562, signal_4145}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6992 ( .a ({signal_10452, signal_7065}), .b ({signal_10563, signal_4148}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6993 ( .a ({signal_10453, signal_7066}), .b ({signal_10564, signal_4149}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_6994 ( .a ({signal_10455, signal_7067}), .b ({signal_10565, signal_4186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6995 ( .a ({signal_10316, signal_6975}), .b ({signal_10404, signal_4404}), .c ({signal_10566, signal_7068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6996 ( .a ({signal_10317, signal_6976}), .b ({signal_10405, signal_7032}), .c ({signal_10567, signal_7069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6997 ( .a ({signal_10318, signal_4391}), .b ({signal_10406, signal_7033}), .c ({signal_10568, signal_7070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6998 ( .a ({signal_10407, signal_4399}), .b ({signal_10504, signal_7045}), .c ({signal_10772, signal_7071}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6999 ( .a ({signal_10408, signal_3879}), .b ({signal_10505, signal_7046}), .c ({signal_10773, signal_7072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7000 ( .a ({signal_10321, signal_6977}), .b ({signal_10409, signal_3880}), .c ({signal_10569, signal_7073}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7001 ( .a ({signal_10129, signal_6836}), .b ({signal_10503, signal_7044}), .c ({signal_10774, signal_7074}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7002 ( .a ({signal_10376, signal_4412}), .b ({signal_10405, signal_7032}), .c ({signal_10570, signal_7075}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7003 ( .a ({signal_10377, signal_7020}), .b ({signal_10406, signal_7033}), .c ({signal_10571, signal_7076}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7004 ( .a ({signal_10378, signal_7021}), .b ({signal_10407, signal_4399}), .c ({signal_10572, signal_7077}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7005 ( .a ({signal_10410, signal_7034}), .b ({signal_10506, signal_7047}), .c ({signal_10775, signal_7078}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7006 ( .a ({signal_10381, signal_3888}), .b ({signal_10410, signal_7034}), .c ({signal_10573, signal_7079}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7007 ( .a ({signal_10184, signal_6891}), .b ({signal_10404, signal_4404}), .c ({signal_10574, signal_7080}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7008 ( .a ({signal_10129, signal_6836}), .b ({signal_10376, signal_4412}), .c ({signal_10575, signal_7081}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7009 ( .a ({signal_10341, signal_4420}), .b ({signal_10377, signal_7020}), .c ({signal_10576, signal_7082}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7010 ( .a ({signal_10315, signal_4396}), .b ({signal_10342, signal_7005}), .c ({signal_10577, signal_7083}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7011 ( .a ({signal_10342, signal_7005}), .b ({signal_10378, signal_7021}), .c ({signal_10578, signal_7084}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7012 ( .a ({signal_10316, signal_6975}), .b ({signal_10343, signal_7006}), .c ({signal_10579, signal_7085}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7013 ( .a ({signal_10343, signal_7006}), .b ({signal_10379, signal_4407}), .c ({signal_10580, signal_7086}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7014 ( .a ({signal_10317, signal_6976}), .b ({signal_10344, signal_4415}), .c ({signal_10581, signal_7087}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7015 ( .a ({signal_10346, signal_3896}), .b ({signal_10382, signal_7022}), .c ({signal_10582, signal_7088}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7016 ( .a ({signal_10320, signal_3872}), .b ({signal_10347, signal_7007}), .c ({signal_10583, signal_7089}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7017 ( .a ({signal_10117, signal_6781}), .b ({signal_10341, signal_4420}), .c ({signal_10584, signal_7090}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7018 ( .a ({signal_10404, signal_4404}), .b ({signal_10408, signal_3879}), .c ({signal_10585, signal_7091}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7019 ( .a ({signal_10404, signal_4404}), .b ({signal_10409, signal_3880}), .c ({signal_10586, signal_7092}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7020 ( .a ({signal_10228, signal_6938}), .b ({signal_10404, signal_4404}), .c ({signal_10587, signal_7093}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7021 ( .a ({signal_10376, signal_4412}), .b ({signal_10380, signal_3887}), .c ({signal_10588, signal_7094}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7022 ( .a ({signal_10376, signal_4412}), .b ({signal_10381, signal_3888}), .c ({signal_10589, signal_7095}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7023 ( .a ({signal_10184, signal_6891}), .b ({signal_10376, signal_4412}), .c ({signal_10590, signal_7096}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7024 ( .a ({signal_10341, signal_4420}), .b ({signal_10345, signal_3895}), .c ({signal_10591, signal_7097}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7025 ( .a ({signal_10341, signal_4420}), .b ({signal_10346, signal_3896}), .c ({signal_10592, signal_7098}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7026 ( .a ({signal_10129, signal_6836}), .b ({signal_10341, signal_4420}), .c ({signal_10593, signal_7099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7027 ( .a ({signal_10309, signal_6939}), .b ({signal_10383, signal_4436}), .c ({signal_10594, signal_7100}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7028 ( .a ({signal_10310, signal_6940}), .b ({signal_10384, signal_7023}), .c ({signal_10595, signal_7101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7029 ( .a ({signal_10311, signal_4423}), .b ({signal_10385, signal_7024}), .c ({signal_10596, signal_7102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7030 ( .a ({signal_10386, signal_4431}), .b ({signal_10508, signal_7049}), .c ({signal_10776, signal_7103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7031 ( .a ({signal_10387, signal_3911}), .b ({signal_10509, signal_7050}), .c ({signal_10777, signal_7104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7032 ( .a ({signal_10314, signal_6941}), .b ({signal_10388, signal_3912}), .c ({signal_10597, signal_7105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7033 ( .a ({signal_10239, signal_6952}), .b ({signal_10507, signal_7048}), .c ({signal_10778, signal_7106}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7034 ( .a ({signal_10348, signal_4444}), .b ({signal_10384, signal_7023}), .c ({signal_10598, signal_7107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7035 ( .a ({signal_10349, signal_7008}), .b ({signal_10385, signal_7024}), .c ({signal_10599, signal_7108}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7036 ( .a ({signal_10350, signal_7009}), .b ({signal_10386, signal_4431}), .c ({signal_10600, signal_7109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7037 ( .a ({signal_10389, signal_7025}), .b ({signal_10510, signal_7051}), .c ({signal_10779, signal_7110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7038 ( .a ({signal_10353, signal_3920}), .b ({signal_10389, signal_7025}), .c ({signal_10601, signal_7111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7039 ( .a ({signal_10140, signal_6847}), .b ({signal_10383, signal_4436}), .c ({signal_10602, signal_7112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7040 ( .a ({signal_10239, signal_6952}), .b ({signal_10348, signal_4444}), .c ({signal_10603, signal_7113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7041 ( .a ({signal_10349, signal_7008}), .b ({signal_10411, signal_4452}), .c ({signal_10604, signal_7114}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7042 ( .a ({signal_10308, signal_4428}), .b ({signal_10412, signal_7035}), .c ({signal_10605, signal_7115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7043 ( .a ({signal_10350, signal_7009}), .b ({signal_10412, signal_7035}), .c ({signal_10606, signal_7116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7044 ( .a ({signal_10309, signal_6939}), .b ({signal_10413, signal_7036}), .c ({signal_10607, signal_7117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7045 ( .a ({signal_10351, signal_4439}), .b ({signal_10413, signal_7036}), .c ({signal_10608, signal_7118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7046 ( .a ({signal_10310, signal_6940}), .b ({signal_10414, signal_4447}), .c ({signal_10609, signal_7119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7047 ( .a ({signal_10354, signal_7010}), .b ({signal_10416, signal_3928}), .c ({signal_10610, signal_7120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7048 ( .a ({signal_10313, signal_3904}), .b ({signal_10417, signal_7037}), .c ({signal_10611, signal_7121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7049 ( .a ({signal_10106, signal_6743}), .b ({signal_10411, signal_4452}), .c ({signal_10612, signal_7122}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7050 ( .a ({signal_10383, signal_4436}), .b ({signal_10387, signal_3911}), .c ({signal_10613, signal_7123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7051 ( .a ({signal_10383, signal_4436}), .b ({signal_10388, signal_3912}), .c ({signal_10614, signal_7124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7052 ( .a ({signal_10195, signal_6902}), .b ({signal_10383, signal_4436}), .c ({signal_10615, signal_7125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7053 ( .a ({signal_10348, signal_4444}), .b ({signal_10352, signal_3919}), .c ({signal_10616, signal_7126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7054 ( .a ({signal_10348, signal_4444}), .b ({signal_10353, signal_3920}), .c ({signal_10617, signal_7127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7055 ( .a ({signal_10140, signal_6847}), .b ({signal_10348, signal_4444}), .c ({signal_10618, signal_7128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7056 ( .a ({signal_10411, signal_4452}), .b ({signal_10415, signal_3927}), .c ({signal_10619, signal_7129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7057 ( .a ({signal_10411, signal_4452}), .b ({signal_10416, signal_3928}), .c ({signal_10620, signal_7130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7058 ( .a ({signal_10239, signal_6952}), .b ({signal_10411, signal_4452}), .c ({signal_10621, signal_7131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7059 ( .a ({signal_10302, signal_6903}), .b ({signal_10355, signal_4468}), .c ({signal_10622, signal_7132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7060 ( .a ({signal_10303, signal_6904}), .b ({signal_10356, signal_7011}), .c ({signal_10623, signal_7133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7061 ( .a ({signal_10304, signal_4455}), .b ({signal_10357, signal_7012}), .c ({signal_10624, signal_7134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7062 ( .a ({signal_10358, signal_4463}), .b ({signal_10512, signal_7053}), .c ({signal_10780, signal_7135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7063 ( .a ({signal_10359, signal_3943}), .b ({signal_10513, signal_7054}), .c ({signal_10781, signal_7136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7064 ( .a ({signal_10307, signal_6905}), .b ({signal_10360, signal_3944}), .c ({signal_10625, signal_7137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7065 ( .a ({signal_10206, signal_6916}), .b ({signal_10511, signal_7052}), .c ({signal_10782, signal_7138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7066 ( .a ({signal_10356, signal_7011}), .b ({signal_10418, signal_4476}), .c ({signal_10626, signal_7139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7067 ( .a ({signal_10357, signal_7012}), .b ({signal_10419, signal_7038}), .c ({signal_10627, signal_7140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7068 ( .a ({signal_10358, signal_4463}), .b ({signal_10420, signal_7039}), .c ({signal_10628, signal_7141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7069 ( .a ({signal_10361, signal_7013}), .b ({signal_10514, signal_7055}), .c ({signal_10783, signal_7142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7070 ( .a ({signal_10361, signal_7013}), .b ({signal_10423, signal_3952}), .c ({signal_10629, signal_7143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7071 ( .a ({signal_10250, signal_6963}), .b ({signal_10355, signal_4468}), .c ({signal_10630, signal_7144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7072 ( .a ({signal_10206, signal_6916}), .b ({signal_10418, signal_4476}), .c ({signal_10631, signal_7145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7073 ( .a ({signal_10390, signal_4484}), .b ({signal_10419, signal_7038}), .c ({signal_10632, signal_7146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7074 ( .a ({signal_10301, signal_4460}), .b ({signal_10391, signal_7026}), .c ({signal_10633, signal_7147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7075 ( .a ({signal_10391, signal_7026}), .b ({signal_10420, signal_7039}), .c ({signal_10634, signal_7148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7076 ( .a ({signal_10302, signal_6903}), .b ({signal_10392, signal_7027}), .c ({signal_10635, signal_7149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7077 ( .a ({signal_10392, signal_7027}), .b ({signal_10421, signal_4471}), .c ({signal_10636, signal_7150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7078 ( .a ({signal_10303, signal_6904}), .b ({signal_10393, signal_4479}), .c ({signal_10637, signal_7151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7079 ( .a ({signal_10395, signal_3960}), .b ({signal_10424, signal_7040}), .c ({signal_10638, signal_7152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7080 ( .a ({signal_10306, signal_3936}), .b ({signal_10396, signal_7028}), .c ({signal_10639, signal_7153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7081 ( .a ({signal_10095, signal_6705}), .b ({signal_10390, signal_4484}), .c ({signal_10640, signal_7154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7082 ( .a ({signal_10355, signal_4468}), .b ({signal_10359, signal_3943}), .c ({signal_10641, signal_7155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7083 ( .a ({signal_10355, signal_4468}), .b ({signal_10360, signal_3944}), .c ({signal_10642, signal_7156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7084 ( .a ({signal_10151, signal_6858}), .b ({signal_10355, signal_4468}), .c ({signal_10643, signal_7157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7085 ( .a ({signal_10418, signal_4476}), .b ({signal_10422, signal_3951}), .c ({signal_10644, signal_7158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7086 ( .a ({signal_10418, signal_4476}), .b ({signal_10423, signal_3952}), .c ({signal_10645, signal_7159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7087 ( .a ({signal_10250, signal_6963}), .b ({signal_10418, signal_4476}), .c ({signal_10646, signal_7160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7088 ( .a ({signal_10390, signal_4484}), .b ({signal_10394, signal_3959}), .c ({signal_10647, signal_7161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7089 ( .a ({signal_10390, signal_4484}), .b ({signal_10395, signal_3960}), .c ({signal_10648, signal_7162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7090 ( .a ({signal_10206, signal_6916}), .b ({signal_10390, signal_4484}), .c ({signal_10649, signal_7163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7091 ( .a ({signal_10363, signal_7014}), .b ({signal_10425, signal_4500}), .c ({signal_10650, signal_7164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7092 ( .a ({signal_10364, signal_7015}), .b ({signal_10426, signal_7041}), .c ({signal_10651, signal_7165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7093 ( .a ({signal_10365, signal_4487}), .b ({signal_10427, signal_7042}), .c ({signal_10652, signal_7166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7094 ( .a ({signal_10368, signal_7016}), .b ({signal_10430, signal_3976}), .c ({signal_10653, signal_7167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7095 ( .a ({signal_10397, signal_4508}), .b ({signal_10426, signal_7041}), .c ({signal_10654, signal_7168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7096 ( .a ({signal_10398, signal_7029}), .b ({signal_10427, signal_7042}), .c ({signal_10655, signal_7169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7097 ( .a ({signal_10399, signal_7030}), .b ({signal_10428, signal_4495}), .c ({signal_10656, signal_7170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7098 ( .a ({signal_10402, signal_3984}), .b ({signal_10431, signal_7043}), .c ({signal_10657, signal_7171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7099 ( .a ({signal_10217, signal_6927}), .b ({signal_10425, signal_4500}), .c ({signal_10658, signal_7172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7100 ( .a ({signal_10173, signal_6880}), .b ({signal_10397, signal_4508}), .c ({signal_10659, signal_7173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7101 ( .a ({signal_10369, signal_4516}), .b ({signal_10398, signal_7029}), .c ({signal_10660, signal_7174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7102 ( .a ({signal_10362, signal_4492}), .b ({signal_10370, signal_7017}), .c ({signal_10661, signal_7175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7103 ( .a ({signal_10370, signal_7017}), .b ({signal_10399, signal_7030}), .c ({signal_10662, signal_7176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7104 ( .a ({signal_10363, signal_7014}), .b ({signal_10371, signal_7018}), .c ({signal_10663, signal_7177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7105 ( .a ({signal_10371, signal_7018}), .b ({signal_10400, signal_4503}), .c ({signal_10664, signal_7178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7106 ( .a ({signal_10364, signal_7015}), .b ({signal_10372, signal_4511}), .c ({signal_10665, signal_7179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7107 ( .a ({signal_10374, signal_3992}), .b ({signal_10403, signal_7031}), .c ({signal_10666, signal_7180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7108 ( .a ({signal_10367, signal_3968}), .b ({signal_10375, signal_7019}), .c ({signal_10667, signal_7181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7109 ( .a ({signal_10261, signal_6974}), .b ({signal_10362, signal_4492}), .c ({signal_10668, signal_7182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7110 ( .a ({signal_10162, signal_6869}), .b ({signal_10369, signal_4516}), .c ({signal_10669, signal_7183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7111 ( .a ({signal_10362, signal_4492}), .b ({signal_10366, signal_3967}), .c ({signal_10670, signal_7184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7112 ( .a ({signal_10362, signal_4492}), .b ({signal_10367, signal_3968}), .c ({signal_10671, signal_7185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7113 ( .a ({signal_10162, signal_6869}), .b ({signal_10362, signal_4492}), .c ({signal_10672, signal_7186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7114 ( .a ({signal_10425, signal_4500}), .b ({signal_10429, signal_3975}), .c ({signal_10673, signal_7187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7115 ( .a ({signal_10425, signal_4500}), .b ({signal_10430, signal_3976}), .c ({signal_10674, signal_7188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7116 ( .a ({signal_10261, signal_6974}), .b ({signal_10425, signal_4500}), .c ({signal_10675, signal_7189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7117 ( .a ({signal_10397, signal_4508}), .b ({signal_10401, signal_3983}), .c ({signal_10676, signal_7190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7118 ( .a ({signal_10397, signal_4508}), .b ({signal_10402, signal_3984}), .c ({signal_10677, signal_7191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7119 ( .a ({signal_10217, signal_6927}), .b ({signal_10397, signal_4508}), .c ({signal_10678, signal_7192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7120 ( .a ({signal_10369, signal_4516}), .b ({signal_10373, signal_3991}), .c ({signal_10679, signal_7193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7121 ( .a ({signal_10369, signal_4516}), .b ({signal_10374, signal_3992}), .c ({signal_10680, signal_7194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7122 ( .a ({signal_10173, signal_6880}), .b ({signal_10369, signal_4516}), .c ({signal_10681, signal_7195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7123 ( .a ({signal_22920, signal_22912}), .b ({signal_10450, signal_7064}), .c ({signal_10682, signal_7196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7124 ( .a ({signal_22936, signal_22928}), .b ({signal_10432, signal_7056}), .c ({signal_10683, signal_7197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7125 ( .a ({signal_22952, signal_22944}), .b ({signal_10451, signal_4147}), .c ({signal_10684, signal_4179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7126 ( .a ({signal_22968, signal_22960}), .b ({signal_10452, signal_7065}), .c ({signal_10685, signal_7198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7127 ( .a ({signal_22984, signal_22976}), .b ({signal_10453, signal_7066}), .c ({signal_10686, signal_7199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7128 ( .a ({signal_23000, signal_22992}), .b ({signal_10454, signal_4150}), .c ({signal_10687, signal_4182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7129 ( .a ({signal_23016, signal_23008}), .b ({signal_10433, signal_4151}), .c ({signal_10688, signal_4183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7130 ( .a ({signal_23032, signal_23024}), .b ({signal_10434, signal_4152}), .c ({signal_10689, signal_4184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7131 ( .a ({signal_23048, signal_23040}), .b ({signal_10437, signal_4131}), .c ({signal_10690, signal_4163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7132 ( .a ({signal_23064, signal_23056}), .b ({signal_10438, signal_7059}), .c ({signal_10691, signal_7200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7133 ( .a ({signal_23080, signal_23072}), .b ({signal_10439, signal_7060}), .c ({signal_10692, signal_7201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7134 ( .a ({signal_23096, signal_23088}), .b ({signal_10440, signal_4134}), .c ({signal_10693, signal_4166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7135 ( .a ({signal_23112, signal_23104}), .b ({signal_10435, signal_7057}), .c ({signal_10694, signal_7202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7136 ( .a ({signal_23128, signal_23120}), .b ({signal_10441, signal_4135}), .c ({signal_10695, signal_4167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7137 ( .a ({signal_23144, signal_23136}), .b ({signal_10442, signal_4136}), .c ({signal_10696, signal_4168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7138 ( .a ({signal_23160, signal_23152}), .b ({signal_10443, signal_7061}), .c ({signal_10697, signal_7203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7139 ( .a ({signal_23176, signal_23168}), .b ({signal_10436, signal_7058}), .c ({signal_10698, signal_7204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7140 ( .a ({signal_23192, signal_23184}), .b ({signal_10444, signal_4139}), .c ({signal_10699, signal_4171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7141 ( .a ({signal_23208, signal_23200}), .b ({signal_10445, signal_7062}), .c ({signal_10700, signal_7205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7142 ( .a ({signal_23224, signal_23216}), .b ({signal_10446, signal_7063}), .c ({signal_10701, signal_7206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7143 ( .a ({signal_23240, signal_23232}), .b ({signal_10447, signal_4142}), .c ({signal_10702, signal_4174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7144 ( .a ({signal_23256, signal_23248}), .b ({signal_10448, signal_4143}), .c ({signal_10703, signal_4175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7145 ( .a ({signal_23272, signal_23264}), .b ({signal_10449, signal_4144}), .c ({signal_10704, signal_4176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7146 ( .a ({signal_23288, signal_23280}), .b ({signal_10455, signal_7067}), .c ({signal_10705, signal_7207}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7147 ( .a ({signal_10682, signal_7196}), .b ({signal_10784, signal_4177}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7148 ( .a ({signal_10683, signal_7197}), .b ({signal_10785, signal_4210}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7149 ( .a ({signal_10685, signal_7198}), .b ({signal_10786, signal_4180}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7150 ( .a ({signal_10686, signal_7199}), .b ({signal_10787, signal_4181}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7151 ( .a ({signal_10691, signal_7200}), .b ({signal_10788, signal_4164}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7152 ( .a ({signal_10692, signal_7201}), .b ({signal_10789, signal_4165}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7153 ( .a ({signal_10694, signal_7202}), .b ({signal_10790, signal_4185}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7154 ( .a ({signal_10697, signal_7203}), .b ({signal_10791, signal_4169}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7155 ( .a ({signal_10698, signal_7204}), .b ({signal_10792, signal_4202}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7156 ( .a ({signal_10700, signal_7205}), .b ({signal_10793, signal_4172}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7157 ( .a ({signal_10701, signal_7206}), .b ({signal_10794, signal_4173}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7158 ( .a ({signal_10705, signal_7207}), .b ({signal_10795, signal_4218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7159 ( .a ({signal_10228, signal_6938}), .b ({signal_10584, signal_7090}), .c ({signal_10796, signal_7208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7160 ( .a ({signal_10376, signal_4412}), .b ({signal_10577, signal_7083}), .c ({signal_10797, signal_7209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7161 ( .a ({signal_10377, signal_7020}), .b ({signal_10579, signal_7085}), .c ({signal_10798, signal_7210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7162 ( .a ({signal_10378, signal_7021}), .b ({signal_10581, signal_7087}), .c ({signal_10799, signal_7211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7163 ( .a ({signal_10341, signal_4420}), .b ({signal_10570, signal_7075}), .c ({signal_10800, signal_7212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7164 ( .a ({signal_10342, signal_7005}), .b ({signal_10571, signal_7076}), .c ({signal_10801, signal_7213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7165 ( .a ({signal_10381, signal_3888}), .b ({signal_10583, signal_7089}), .c ({signal_10802, signal_7214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7166 ( .a ({signal_10343, signal_7006}), .b ({signal_10572, signal_7077}), .c ({signal_10803, signal_7215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7167 ( .a ({signal_10346, signal_3896}), .b ({signal_10573, signal_7079}), .c ({signal_10804, signal_7216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7168 ( .a ({signal_10774, signal_7074}), .b ({signal_10574, signal_7080}), .c ({signal_11008, signal_7217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7169 ( .a ({signal_10315, signal_4396}), .b ({signal_10576, signal_7082}), .c ({signal_10805, signal_7218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7170 ( .a ({signal_10316, signal_6975}), .b ({signal_10578, signal_7084}), .c ({signal_10806, signal_7219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7171 ( .a ({signal_10317, signal_6976}), .b ({signal_10580, signal_7086}), .c ({signal_10807, signal_7220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7172 ( .a ({signal_10379, signal_4407}), .b ({signal_10585, signal_7091}), .c ({signal_10808, signal_7221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7173 ( .a ({signal_10321, signal_6977}), .b ({signal_10593, signal_7099}), .c ({signal_10809, signal_7222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7174 ( .a ({signal_10380, signal_3887}), .b ({signal_10586, signal_7092}), .c ({signal_10810, signal_7223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7175 ( .a ({signal_10320, signal_3872}), .b ({signal_10582, signal_7088}), .c ({signal_10811, signal_7224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7176 ( .a ({signal_10382, signal_7022}), .b ({signal_10587, signal_7093}), .c ({signal_10812, signal_7225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7177 ( .a ({signal_10347, signal_7007}), .b ({signal_10590, signal_7096}), .c ({signal_10813, signal_7226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7178 ( .a ({signal_10117, signal_6781}), .b ({signal_10575, signal_7081}), .c ({signal_10814, signal_7227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7179 ( .a ({signal_10404, signal_4404}), .b ({signal_10577, signal_7083}), .c ({signal_10815, signal_7228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7180 ( .a ({signal_10405, signal_7032}), .b ({signal_10579, signal_7085}), .c ({signal_10816, signal_7229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7181 ( .a ({signal_10406, signal_7033}), .b ({signal_10581, signal_7087}), .c ({signal_10817, signal_7230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7182 ( .a ({signal_10344, signal_4415}), .b ({signal_10588, signal_7094}), .c ({signal_10818, signal_7231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7183 ( .a ({signal_10318, signal_4391}), .b ({signal_10591, signal_7097}), .c ({signal_10819, signal_7232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7184 ( .a ({signal_10345, signal_3895}), .b ({signal_10589, signal_7095}), .c ({signal_10820, signal_7233}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7185 ( .a ({signal_10319, signal_3871}), .b ({signal_10592, signal_7098}), .c ({signal_10821, signal_7234}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7186 ( .a ({signal_10409, signal_3880}), .b ({signal_10583, signal_7089}), .c ({signal_10822, signal_7235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7187 ( .a ({signal_10503, signal_7044}), .b ({signal_10584, signal_7090}), .c ({signal_10823, signal_7236}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7188 ( .a ({signal_10195, signal_6902}), .b ({signal_10612, signal_7122}), .c ({signal_10824, signal_7237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7189 ( .a ({signal_10348, signal_4444}), .b ({signal_10605, signal_7115}), .c ({signal_10825, signal_7238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7190 ( .a ({signal_10349, signal_7008}), .b ({signal_10607, signal_7117}), .c ({signal_10826, signal_7239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7191 ( .a ({signal_10350, signal_7009}), .b ({signal_10609, signal_7119}), .c ({signal_10827, signal_7240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7192 ( .a ({signal_10411, signal_4452}), .b ({signal_10598, signal_7107}), .c ({signal_10828, signal_7241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7193 ( .a ({signal_10412, signal_7035}), .b ({signal_10599, signal_7108}), .c ({signal_10829, signal_7242}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7194 ( .a ({signal_10353, signal_3920}), .b ({signal_10611, signal_7121}), .c ({signal_10830, signal_7243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7195 ( .a ({signal_10413, signal_7036}), .b ({signal_10600, signal_7109}), .c ({signal_10831, signal_7244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7196 ( .a ({signal_10416, signal_3928}), .b ({signal_10601, signal_7111}), .c ({signal_10832, signal_7245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7197 ( .a ({signal_10778, signal_7106}), .b ({signal_10602, signal_7112}), .c ({signal_11009, signal_7246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7198 ( .a ({signal_10308, signal_4428}), .b ({signal_10604, signal_7114}), .c ({signal_10833, signal_7247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7199 ( .a ({signal_10309, signal_6939}), .b ({signal_10606, signal_7116}), .c ({signal_10834, signal_7248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7200 ( .a ({signal_10310, signal_6940}), .b ({signal_10608, signal_7118}), .c ({signal_10835, signal_7249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7201 ( .a ({signal_10351, signal_4439}), .b ({signal_10613, signal_7123}), .c ({signal_10836, signal_7250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7202 ( .a ({signal_10314, signal_6941}), .b ({signal_10621, signal_7131}), .c ({signal_10837, signal_7251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7203 ( .a ({signal_10352, signal_3919}), .b ({signal_10614, signal_7124}), .c ({signal_10838, signal_7252}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7204 ( .a ({signal_10313, signal_3904}), .b ({signal_10610, signal_7120}), .c ({signal_10839, signal_7253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7205 ( .a ({signal_10354, signal_7010}), .b ({signal_10615, signal_7125}), .c ({signal_10840, signal_7254}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7206 ( .a ({signal_10417, signal_7037}), .b ({signal_10618, signal_7128}), .c ({signal_10841, signal_7255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7207 ( .a ({signal_10106, signal_6743}), .b ({signal_10603, signal_7113}), .c ({signal_10842, signal_7256}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7208 ( .a ({signal_10383, signal_4436}), .b ({signal_10605, signal_7115}), .c ({signal_10843, signal_7257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7209 ( .a ({signal_10384, signal_7023}), .b ({signal_10607, signal_7117}), .c ({signal_10844, signal_7258}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7210 ( .a ({signal_10385, signal_7024}), .b ({signal_10609, signal_7119}), .c ({signal_10845, signal_7259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7211 ( .a ({signal_10414, signal_4447}), .b ({signal_10616, signal_7126}), .c ({signal_10846, signal_7260}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7212 ( .a ({signal_10311, signal_4423}), .b ({signal_10619, signal_7129}), .c ({signal_10847, signal_7261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7213 ( .a ({signal_10415, signal_3927}), .b ({signal_10617, signal_7127}), .c ({signal_10848, signal_7262}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7214 ( .a ({signal_10312, signal_3903}), .b ({signal_10620, signal_7130}), .c ({signal_10849, signal_7263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7215 ( .a ({signal_10388, signal_3912}), .b ({signal_10611, signal_7121}), .c ({signal_10850, signal_7264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7216 ( .a ({signal_10507, signal_7048}), .b ({signal_10612, signal_7122}), .c ({signal_10851, signal_7265}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7217 ( .a ({signal_10151, signal_6858}), .b ({signal_10640, signal_7154}), .c ({signal_10852, signal_7266}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7218 ( .a ({signal_10418, signal_4476}), .b ({signal_10633, signal_7147}), .c ({signal_10853, signal_7267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7219 ( .a ({signal_10419, signal_7038}), .b ({signal_10635, signal_7149}), .c ({signal_10854, signal_7268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7220 ( .a ({signal_10420, signal_7039}), .b ({signal_10637, signal_7151}), .c ({signal_10855, signal_7269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7221 ( .a ({signal_10390, signal_4484}), .b ({signal_10626, signal_7139}), .c ({signal_10856, signal_7270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7222 ( .a ({signal_10391, signal_7026}), .b ({signal_10627, signal_7140}), .c ({signal_10857, signal_7271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7223 ( .a ({signal_10423, signal_3952}), .b ({signal_10639, signal_7153}), .c ({signal_10858, signal_7272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7224 ( .a ({signal_10392, signal_7027}), .b ({signal_10628, signal_7141}), .c ({signal_10859, signal_7273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7225 ( .a ({signal_10395, signal_3960}), .b ({signal_10629, signal_7143}), .c ({signal_10860, signal_7274}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7226 ( .a ({signal_10782, signal_7138}), .b ({signal_10630, signal_7144}), .c ({signal_11010, signal_7275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7227 ( .a ({signal_10301, signal_4460}), .b ({signal_10632, signal_7146}), .c ({signal_10861, signal_7276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7228 ( .a ({signal_10302, signal_6903}), .b ({signal_10634, signal_7148}), .c ({signal_10862, signal_7277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7229 ( .a ({signal_10303, signal_6904}), .b ({signal_10636, signal_7150}), .c ({signal_10863, signal_7278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7230 ( .a ({signal_10421, signal_4471}), .b ({signal_10641, signal_7155}), .c ({signal_10864, signal_7279}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7231 ( .a ({signal_10307, signal_6905}), .b ({signal_10649, signal_7163}), .c ({signal_10865, signal_7280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7232 ( .a ({signal_10422, signal_3951}), .b ({signal_10642, signal_7156}), .c ({signal_10866, signal_7281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7233 ( .a ({signal_10306, signal_3936}), .b ({signal_10638, signal_7152}), .c ({signal_10867, signal_7282}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7234 ( .a ({signal_10424, signal_7040}), .b ({signal_10643, signal_7157}), .c ({signal_10868, signal_7283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7235 ( .a ({signal_10396, signal_7028}), .b ({signal_10646, signal_7160}), .c ({signal_10869, signal_7284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7236 ( .a ({signal_10095, signal_6705}), .b ({signal_10631, signal_7145}), .c ({signal_10870, signal_7285}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7237 ( .a ({signal_10355, signal_4468}), .b ({signal_10633, signal_7147}), .c ({signal_10871, signal_7286}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7238 ( .a ({signal_10356, signal_7011}), .b ({signal_10635, signal_7149}), .c ({signal_10872, signal_7287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7239 ( .a ({signal_10357, signal_7012}), .b ({signal_10637, signal_7151}), .c ({signal_10873, signal_7288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7240 ( .a ({signal_10393, signal_4479}), .b ({signal_10644, signal_7158}), .c ({signal_10874, signal_7289}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7241 ( .a ({signal_10304, signal_4455}), .b ({signal_10647, signal_7161}), .c ({signal_10875, signal_7290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7242 ( .a ({signal_10394, signal_3959}), .b ({signal_10645, signal_7159}), .c ({signal_10876, signal_7291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7243 ( .a ({signal_10305, signal_3935}), .b ({signal_10648, signal_7162}), .c ({signal_10877, signal_7292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7244 ( .a ({signal_10360, signal_3944}), .b ({signal_10639, signal_7153}), .c ({signal_10878, signal_7293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7245 ( .a ({signal_10511, signal_7052}), .b ({signal_10640, signal_7154}), .c ({signal_10879, signal_7294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7246 ( .a ({signal_10261, signal_6974}), .b ({signal_10669, signal_7183}), .c ({signal_10880, signal_7295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7247 ( .a ({signal_10397, signal_4508}), .b ({signal_10661, signal_7175}), .c ({signal_10881, signal_7296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7248 ( .a ({signal_10398, signal_7029}), .b ({signal_10663, signal_7177}), .c ({signal_10882, signal_7297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7249 ( .a ({signal_10399, signal_7030}), .b ({signal_10665, signal_7179}), .c ({signal_10883, signal_7298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7250 ( .a ({signal_10369, signal_4516}), .b ({signal_10654, signal_7168}), .c ({signal_10884, signal_7299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7251 ( .a ({signal_10370, signal_7017}), .b ({signal_10655, signal_7169}), .c ({signal_10885, signal_7300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7252 ( .a ({signal_10402, signal_3984}), .b ({signal_10667, signal_7181}), .c ({signal_10886, signal_7301}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7253 ( .a ({signal_10371, signal_7018}), .b ({signal_10656, signal_7170}), .c ({signal_10887, signal_7302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7254 ( .a ({signal_10428, signal_4495}), .b ({signal_10670, signal_7184}), .c ({signal_10888, signal_7303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7255 ( .a ({signal_10429, signal_3975}), .b ({signal_10671, signal_7185}), .c ({signal_10889, signal_7304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7256 ( .a ({signal_10374, signal_3992}), .b ({signal_10657, signal_7171}), .c ({signal_10890, signal_7305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7257 ( .a ({signal_10173, signal_6880}), .b ({signal_10668, signal_7182}), .c ({signal_10891, signal_7306}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7258 ( .a ({signal_10362, signal_4492}), .b ({signal_10660, signal_7174}), .c ({signal_10892, signal_7307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7259 ( .a ({signal_10363, signal_7014}), .b ({signal_10662, signal_7176}), .c ({signal_10893, signal_7308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7260 ( .a ({signal_10364, signal_7015}), .b ({signal_10664, signal_7178}), .c ({signal_10894, signal_7309}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7261 ( .a ({signal_10400, signal_4503}), .b ({signal_10673, signal_7187}), .c ({signal_10895, signal_7310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7262 ( .a ({signal_10431, signal_7043}), .b ({signal_10672, signal_7186}), .c ({signal_10896, signal_7311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7263 ( .a ({signal_10368, signal_7016}), .b ({signal_10681, signal_7195}), .c ({signal_10897, signal_7312}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7264 ( .a ({signal_10401, signal_3983}), .b ({signal_10674, signal_7188}), .c ({signal_10898, signal_7313}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7265 ( .a ({signal_10367, signal_3968}), .b ({signal_10666, signal_7180}), .c ({signal_10899, signal_7314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7266 ( .a ({signal_10403, signal_7031}), .b ({signal_10675, signal_7189}), .c ({signal_10900, signal_7315}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7267 ( .a ({signal_10375, signal_7019}), .b ({signal_10678, signal_7192}), .c ({signal_10901, signal_7316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7268 ( .a ({signal_10162, signal_6869}), .b ({signal_10659, signal_7173}), .c ({signal_10902, signal_7317}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7269 ( .a ({signal_10425, signal_4500}), .b ({signal_10661, signal_7175}), .c ({signal_10903, signal_7318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7270 ( .a ({signal_10426, signal_7041}), .b ({signal_10663, signal_7177}), .c ({signal_10904, signal_7319}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7271 ( .a ({signal_10427, signal_7042}), .b ({signal_10665, signal_7179}), .c ({signal_10905, signal_7320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7272 ( .a ({signal_10372, signal_4511}), .b ({signal_10676, signal_7190}), .c ({signal_10906, signal_7321}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7273 ( .a ({signal_10365, signal_4487}), .b ({signal_10679, signal_7193}), .c ({signal_10907, signal_7322}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7274 ( .a ({signal_10373, signal_3991}), .b ({signal_10677, signal_7191}), .c ({signal_10908, signal_7323}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7275 ( .a ({signal_10366, signal_3967}), .b ({signal_10680, signal_7194}), .c ({signal_10909, signal_7324}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7276 ( .a ({signal_10430, signal_3976}), .b ({signal_10667, signal_7181}), .c ({signal_10910, signal_7325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7277 ( .a ({signal_10668, signal_7182}), .b ({signal_10669, signal_7183}), .c ({signal_10911, signal_7326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7278 ( .a ({signal_23292, signal_23290}), .b ({signal_10683, signal_7197}), .c ({signal_10912, signal_7327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7279 ( .a ({signal_23308, signal_23300}), .b ({signal_10682, signal_7196}), .c ({signal_10913, signal_7328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7280 ( .a ({signal_23324, signal_23316}), .b ({signal_10684, signal_4179}), .c ({signal_10914, signal_4211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7281 ( .a ({signal_23340, signal_23332}), .b ({signal_10685, signal_7198}), .c ({signal_10915, signal_7329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7282 ( .a ({signal_23356, signal_23348}), .b ({signal_10686, signal_7199}), .c ({signal_10916, signal_7330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7283 ( .a ({signal_23372, signal_23364}), .b ({signal_10687, signal_4182}), .c ({signal_10917, signal_4214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7284 ( .a ({signal_23388, signal_23380}), .b ({signal_10688, signal_4183}), .c ({signal_10918, signal_4215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7285 ( .a ({signal_23404, signal_23396}), .b ({signal_10689, signal_4184}), .c ({signal_10919, signal_4216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7286 ( .a ({signal_23420, signal_23412}), .b ({signal_10690, signal_4163}), .c ({signal_10920, signal_4195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7287 ( .a ({signal_23436, signal_23428}), .b ({signal_10691, signal_7200}), .c ({signal_10921, signal_7331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7288 ( .a ({signal_23452, signal_23444}), .b ({signal_10692, signal_7201}), .c ({signal_10922, signal_7332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7289 ( .a ({signal_23468, signal_23460}), .b ({signal_10693, signal_4166}), .c ({signal_10923, signal_4198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7290 ( .a ({signal_23484, signal_23476}), .b ({signal_10694, signal_7202}), .c ({signal_10924, signal_7333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7291 ( .a ({signal_23500, signal_23492}), .b ({signal_10695, signal_4167}), .c ({signal_10925, signal_4199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7292 ( .a ({signal_23516, signal_23508}), .b ({signal_10696, signal_4168}), .c ({signal_10926, signal_4200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7293 ( .a ({signal_23532, signal_23524}), .b ({signal_10697, signal_7203}), .c ({signal_10927, signal_7334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7294 ( .a ({signal_23536, signal_23534}), .b ({signal_10698, signal_7204}), .c ({signal_10928, signal_7335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7295 ( .a ({signal_23552, signal_23544}), .b ({signal_10699, signal_4171}), .c ({signal_10929, signal_4203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7296 ( .a ({signal_23568, signal_23560}), .b ({signal_10700, signal_7205}), .c ({signal_10930, signal_7336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7297 ( .a ({signal_23584, signal_23576}), .b ({signal_10701, signal_7206}), .c ({signal_10931, signal_7337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7298 ( .a ({signal_23600, signal_23592}), .b ({signal_10702, signal_4174}), .c ({signal_10932, signal_4206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7299 ( .a ({signal_23616, signal_23608}), .b ({signal_10703, signal_4175}), .c ({signal_10933, signal_4207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7300 ( .a ({signal_23632, signal_23624}), .b ({signal_10704, signal_4176}), .c ({signal_10934, signal_4208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7301 ( .a ({signal_23636, signal_23634}), .b ({signal_10705, signal_7207}), .c ({signal_10935, signal_7338}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7302 ( .a ({signal_11008, signal_7217}), .b ({signal_11273, signal_4002}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7303 ( .a ({signal_11009, signal_7246}), .b ({signal_11274, signal_4034}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7304 ( .a ({signal_11010, signal_7275}), .b ({signal_11275, signal_4066}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7305 ( .a ({signal_10912, signal_7327}), .b ({signal_11011, signal_4242}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7306 ( .a ({signal_10913, signal_7328}), .b ({signal_11012, signal_4209}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7307 ( .a ({signal_10915, signal_7329}), .b ({signal_11013, signal_4212}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7308 ( .a ({signal_10916, signal_7330}), .b ({signal_11014, signal_4213}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7309 ( .a ({signal_10921, signal_7331}), .b ({signal_11015, signal_4196}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7310 ( .a ({signal_10922, signal_7332}), .b ({signal_11016, signal_4197}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7311 ( .a ({signal_10924, signal_7333}), .b ({signal_11017, signal_4217}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7312 ( .a ({signal_10927, signal_7334}), .b ({signal_11018, signal_4201}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7313 ( .a ({signal_10928, signal_7335}), .b ({signal_11019, signal_4234}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7314 ( .a ({signal_10930, signal_7336}), .b ({signal_11020, signal_4204}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7315 ( .a ({signal_10931, signal_7337}), .b ({signal_11021, signal_4205}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7316 ( .a ({signal_10935, signal_7338}), .b ({signal_11022, signal_4250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7317 ( .a ({signal_10809, signal_7222}), .b ({signal_10813, signal_7226}), .c ({signal_11023, signal_7339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7318 ( .a ({signal_10575, signal_7081}), .b ({signal_10796, signal_7208}), .c ({signal_11024, signal_7340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7319 ( .a ({signal_10566, signal_7068}), .b ({signal_10797, signal_7209}), .c ({signal_11025, signal_4019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7320 ( .a ({signal_10567, signal_7069}), .b ({signal_10798, signal_7210}), .c ({signal_11026, signal_7341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7321 ( .a ({signal_10568, signal_7070}), .b ({signal_10799, signal_7211}), .c ({signal_11027, signal_7342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7322 ( .a ({signal_10379, signal_4407}), .b ({signal_10819, signal_7232}), .c ({signal_11028, signal_7343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7323 ( .a ({signal_10380, signal_3887}), .b ({signal_10821, signal_7234}), .c ({signal_11029, signal_7344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7324 ( .a ({signal_10566, signal_7068}), .b ({signal_10800, signal_7212}), .c ({signal_11030, signal_3995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7325 ( .a ({signal_10567, signal_7069}), .b ({signal_10801, signal_7213}), .c ({signal_11031, signal_7345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7326 ( .a ({signal_10569, signal_7073}), .b ({signal_10802, signal_7214}), .c ({signal_11032, signal_4024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7327 ( .a ({signal_10568, signal_7070}), .b ({signal_10803, signal_7215}), .c ({signal_11033, signal_7346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7328 ( .a ({signal_10344, signal_4415}), .b ({signal_10808, signal_7221}), .c ({signal_11034, signal_7347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7329 ( .a ({signal_10345, signal_3895}), .b ({signal_10810, signal_7223}), .c ({signal_11035, signal_7348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7330 ( .a ({signal_10569, signal_7073}), .b ({signal_10804, signal_7216}), .c ({signal_11036, signal_4000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7331 ( .a ({signal_10347, signal_7007}), .b ({signal_10812, signal_7225}), .c ({signal_11037, signal_7349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7332 ( .a ({signal_10570, signal_7075}), .b ({signal_10805, signal_7218}), .c ({signal_11038, signal_4003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7333 ( .a ({signal_10571, signal_7076}), .b ({signal_10806, signal_7219}), .c ({signal_11039, signal_7350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7334 ( .a ({signal_10572, signal_7077}), .b ({signal_10807, signal_7220}), .c ({signal_11040, signal_7351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7335 ( .a ({signal_10318, signal_4391}), .b ({signal_10818, signal_7231}), .c ({signal_11041, signal_7352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7336 ( .a ({signal_10382, signal_7022}), .b ({signal_10809, signal_7222}), .c ({signal_11042, signal_7353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7337 ( .a ({signal_10319, signal_3871}), .b ({signal_10820, signal_7233}), .c ({signal_11043, signal_7354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7338 ( .a ({signal_10573, signal_7079}), .b ({signal_10811, signal_7224}), .c ({signal_11044, signal_4008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7339 ( .a ({signal_10321, signal_6977}), .b ({signal_10813, signal_7226}), .c ({signal_11045, signal_7355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7340 ( .a ({signal_10574, signal_7080}), .b ({signal_10814, signal_7227}), .c ({signal_11046, signal_7356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7341 ( .a ({signal_10576, signal_7082}), .b ({signal_10815, signal_7228}), .c ({signal_11047, signal_4011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7342 ( .a ({signal_10578, signal_7084}), .b ({signal_10816, signal_7229}), .c ({signal_11048, signal_7357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7343 ( .a ({signal_10580, signal_7086}), .b ({signal_10817, signal_7230}), .c ({signal_11049, signal_7358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7344 ( .a ({signal_10407, signal_4399}), .b ({signal_10819, signal_7232}), .c ({signal_11050, signal_7359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7345 ( .a ({signal_10408, signal_3879}), .b ({signal_10821, signal_7234}), .c ({signal_11051, signal_7360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7346 ( .a ({signal_10582, signal_7088}), .b ({signal_10822, signal_7235}), .c ({signal_11052, signal_4016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7347 ( .a ({signal_10184, signal_6891}), .b ({signal_10823, signal_7236}), .c ({signal_11053, signal_7361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7348 ( .a ({signal_10837, signal_7251}), .b ({signal_10841, signal_7255}), .c ({signal_11054, signal_7362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7349 ( .a ({signal_10603, signal_7113}), .b ({signal_10824, signal_7237}), .c ({signal_11055, signal_7363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7350 ( .a ({signal_10594, signal_7100}), .b ({signal_10825, signal_7238}), .c ({signal_11056, signal_4051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7351 ( .a ({signal_10595, signal_7101}), .b ({signal_10826, signal_7239}), .c ({signal_11057, signal_7364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7352 ( .a ({signal_10596, signal_7102}), .b ({signal_10827, signal_7240}), .c ({signal_11058, signal_7365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7353 ( .a ({signal_10351, signal_4439}), .b ({signal_10847, signal_7261}), .c ({signal_11059, signal_7366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7354 ( .a ({signal_10352, signal_3919}), .b ({signal_10849, signal_7263}), .c ({signal_11060, signal_7367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7355 ( .a ({signal_10594, signal_7100}), .b ({signal_10828, signal_7241}), .c ({signal_11061, signal_4027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7356 ( .a ({signal_10595, signal_7101}), .b ({signal_10829, signal_7242}), .c ({signal_11062, signal_7368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7357 ( .a ({signal_10597, signal_7105}), .b ({signal_10830, signal_7243}), .c ({signal_11063, signal_4056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7358 ( .a ({signal_10596, signal_7102}), .b ({signal_10831, signal_7244}), .c ({signal_11064, signal_7369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7359 ( .a ({signal_10414, signal_4447}), .b ({signal_10836, signal_7250}), .c ({signal_11065, signal_7370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7360 ( .a ({signal_10415, signal_3927}), .b ({signal_10838, signal_7252}), .c ({signal_11066, signal_7371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7361 ( .a ({signal_10597, signal_7105}), .b ({signal_10832, signal_7245}), .c ({signal_11067, signal_4032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7362 ( .a ({signal_10417, signal_7037}), .b ({signal_10840, signal_7254}), .c ({signal_11068, signal_7372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7363 ( .a ({signal_10598, signal_7107}), .b ({signal_10833, signal_7247}), .c ({signal_11069, signal_4035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7364 ( .a ({signal_10599, signal_7108}), .b ({signal_10834, signal_7248}), .c ({signal_11070, signal_7373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7365 ( .a ({signal_10600, signal_7109}), .b ({signal_10835, signal_7249}), .c ({signal_11071, signal_7374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7366 ( .a ({signal_10311, signal_4423}), .b ({signal_10846, signal_7260}), .c ({signal_11072, signal_7375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7367 ( .a ({signal_10354, signal_7010}), .b ({signal_10837, signal_7251}), .c ({signal_11073, signal_7376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7368 ( .a ({signal_10312, signal_3903}), .b ({signal_10848, signal_7262}), .c ({signal_11074, signal_7377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7369 ( .a ({signal_10601, signal_7111}), .b ({signal_10839, signal_7253}), .c ({signal_11075, signal_4040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7370 ( .a ({signal_10314, signal_6941}), .b ({signal_10841, signal_7255}), .c ({signal_11076, signal_7378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7371 ( .a ({signal_10602, signal_7112}), .b ({signal_10842, signal_7256}), .c ({signal_11077, signal_7379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7372 ( .a ({signal_10604, signal_7114}), .b ({signal_10843, signal_7257}), .c ({signal_11078, signal_4043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7373 ( .a ({signal_10606, signal_7116}), .b ({signal_10844, signal_7258}), .c ({signal_11079, signal_7380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7374 ( .a ({signal_10608, signal_7118}), .b ({signal_10845, signal_7259}), .c ({signal_11080, signal_7381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7375 ( .a ({signal_10386, signal_4431}), .b ({signal_10847, signal_7261}), .c ({signal_11081, signal_7382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7376 ( .a ({signal_10387, signal_3911}), .b ({signal_10849, signal_7263}), .c ({signal_11082, signal_7383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7377 ( .a ({signal_10610, signal_7120}), .b ({signal_10850, signal_7264}), .c ({signal_11083, signal_4048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7378 ( .a ({signal_10140, signal_6847}), .b ({signal_10851, signal_7265}), .c ({signal_11084, signal_7384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7379 ( .a ({signal_10865, signal_7280}), .b ({signal_10869, signal_7284}), .c ({signal_11085, signal_7385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7380 ( .a ({signal_10631, signal_7145}), .b ({signal_10852, signal_7266}), .c ({signal_11086, signal_7386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7381 ( .a ({signal_10622, signal_7132}), .b ({signal_10853, signal_7267}), .c ({signal_11087, signal_4083}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7382 ( .a ({signal_10623, signal_7133}), .b ({signal_10854, signal_7268}), .c ({signal_11088, signal_7387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7383 ( .a ({signal_10624, signal_7134}), .b ({signal_10855, signal_7269}), .c ({signal_11089, signal_7388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7384 ( .a ({signal_10421, signal_4471}), .b ({signal_10875, signal_7290}), .c ({signal_11090, signal_7389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7385 ( .a ({signal_10422, signal_3951}), .b ({signal_10877, signal_7292}), .c ({signal_11091, signal_7390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7386 ( .a ({signal_10622, signal_7132}), .b ({signal_10856, signal_7270}), .c ({signal_11092, signal_4059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7387 ( .a ({signal_10623, signal_7133}), .b ({signal_10857, signal_7271}), .c ({signal_11093, signal_7391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7388 ( .a ({signal_10625, signal_7137}), .b ({signal_10858, signal_7272}), .c ({signal_11094, signal_4088}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7389 ( .a ({signal_10624, signal_7134}), .b ({signal_10859, signal_7273}), .c ({signal_11095, signal_7392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7390 ( .a ({signal_10393, signal_4479}), .b ({signal_10864, signal_7279}), .c ({signal_11096, signal_7393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7391 ( .a ({signal_10394, signal_3959}), .b ({signal_10866, signal_7281}), .c ({signal_11097, signal_7394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7392 ( .a ({signal_10625, signal_7137}), .b ({signal_10860, signal_7274}), .c ({signal_11098, signal_4064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7393 ( .a ({signal_10396, signal_7028}), .b ({signal_10868, signal_7283}), .c ({signal_11099, signal_7395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7394 ( .a ({signal_10626, signal_7139}), .b ({signal_10861, signal_7276}), .c ({signal_11100, signal_4067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7395 ( .a ({signal_10627, signal_7140}), .b ({signal_10862, signal_7277}), .c ({signal_11101, signal_7396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7396 ( .a ({signal_10628, signal_7141}), .b ({signal_10863, signal_7278}), .c ({signal_11102, signal_7397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7397 ( .a ({signal_10304, signal_4455}), .b ({signal_10874, signal_7289}), .c ({signal_11103, signal_7398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7398 ( .a ({signal_10424, signal_7040}), .b ({signal_10865, signal_7280}), .c ({signal_11104, signal_7399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7399 ( .a ({signal_10305, signal_3935}), .b ({signal_10876, signal_7291}), .c ({signal_11105, signal_7400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7400 ( .a ({signal_10629, signal_7143}), .b ({signal_10867, signal_7282}), .c ({signal_11106, signal_4072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7401 ( .a ({signal_10307, signal_6905}), .b ({signal_10869, signal_7284}), .c ({signal_11107, signal_7401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7402 ( .a ({signal_10630, signal_7144}), .b ({signal_10870, signal_7285}), .c ({signal_11108, signal_7402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7403 ( .a ({signal_10632, signal_7146}), .b ({signal_10871, signal_7286}), .c ({signal_11109, signal_4075}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7404 ( .a ({signal_10634, signal_7148}), .b ({signal_10872, signal_7287}), .c ({signal_11110, signal_7403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7405 ( .a ({signal_10636, signal_7150}), .b ({signal_10873, signal_7288}), .c ({signal_11111, signal_7404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7406 ( .a ({signal_10358, signal_4463}), .b ({signal_10875, signal_7290}), .c ({signal_11112, signal_7405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7407 ( .a ({signal_10359, signal_3943}), .b ({signal_10877, signal_7292}), .c ({signal_11113, signal_7406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7408 ( .a ({signal_10638, signal_7152}), .b ({signal_10878, signal_7293}), .c ({signal_11114, signal_4080}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7409 ( .a ({signal_10250, signal_6963}), .b ({signal_10879, signal_7294}), .c ({signal_11115, signal_7407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7410 ( .a ({signal_10897, signal_7312}), .b ({signal_10901, signal_7316}), .c ({signal_11116, signal_7408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7411 ( .a ({signal_10659, signal_7173}), .b ({signal_10880, signal_7295}), .c ({signal_11117, signal_7409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7412 ( .a ({signal_10650, signal_7164}), .b ({signal_10881, signal_7296}), .c ({signal_11118, signal_4115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7413 ( .a ({signal_10651, signal_7165}), .b ({signal_10882, signal_7297}), .c ({signal_11119, signal_7410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7414 ( .a ({signal_10652, signal_7166}), .b ({signal_10883, signal_7298}), .c ({signal_11120, signal_7411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7415 ( .a ({signal_10400, signal_4503}), .b ({signal_10907, signal_7322}), .c ({signal_11121, signal_7412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7416 ( .a ({signal_10401, signal_3983}), .b ({signal_10909, signal_7324}), .c ({signal_11122, signal_7413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7417 ( .a ({signal_10650, signal_7164}), .b ({signal_10884, signal_7299}), .c ({signal_11123, signal_4091}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7418 ( .a ({signal_10651, signal_7165}), .b ({signal_10885, signal_7300}), .c ({signal_11124, signal_7414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7419 ( .a ({signal_10653, signal_7167}), .b ({signal_10886, signal_7301}), .c ({signal_11125, signal_4120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7420 ( .a ({signal_10652, signal_7166}), .b ({signal_10887, signal_7302}), .c ({signal_11126, signal_7415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7421 ( .a ({signal_10372, signal_4511}), .b ({signal_10895, signal_7310}), .c ({signal_11127, signal_7416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7422 ( .a ({signal_10373, signal_3991}), .b ({signal_10898, signal_7313}), .c ({signal_11128, signal_7417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7423 ( .a ({signal_10653, signal_7167}), .b ({signal_10890, signal_7305}), .c ({signal_11129, signal_4096}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7424 ( .a ({signal_10375, signal_7019}), .b ({signal_10900, signal_7315}), .c ({signal_11130, signal_7418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7425 ( .a ({signal_10658, signal_7172}), .b ({signal_10891, signal_7306}), .c ({signal_11131, signal_7419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7426 ( .a ({signal_10654, signal_7168}), .b ({signal_10892, signal_7307}), .c ({signal_11132, signal_4099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7427 ( .a ({signal_10655, signal_7169}), .b ({signal_10893, signal_7308}), .c ({signal_11133, signal_7420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7428 ( .a ({signal_10656, signal_7170}), .b ({signal_10894, signal_7309}), .c ({signal_11134, signal_7421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7429 ( .a ({signal_10365, signal_4487}), .b ({signal_10906, signal_7321}), .c ({signal_11135, signal_7422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7430 ( .a ({signal_10403, signal_7031}), .b ({signal_10897, signal_7312}), .c ({signal_11136, signal_7423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7431 ( .a ({signal_10366, signal_3967}), .b ({signal_10908, signal_7323}), .c ({signal_11137, signal_7424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7432 ( .a ({signal_10657, signal_7171}), .b ({signal_10899, signal_7314}), .c ({signal_11138, signal_4104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7433 ( .a ({signal_10368, signal_7016}), .b ({signal_10901, signal_7316}), .c ({signal_11139, signal_7425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7434 ( .a ({signal_10658, signal_7172}), .b ({signal_10902, signal_7317}), .c ({signal_11140, signal_7426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7435 ( .a ({signal_10660, signal_7174}), .b ({signal_10903, signal_7318}), .c ({signal_11141, signal_4107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7436 ( .a ({signal_10662, signal_7176}), .b ({signal_10904, signal_7319}), .c ({signal_11142, signal_7427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7437 ( .a ({signal_10664, signal_7178}), .b ({signal_10905, signal_7320}), .c ({signal_11143, signal_7428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7438 ( .a ({signal_10428, signal_4495}), .b ({signal_10907, signal_7322}), .c ({signal_11144, signal_7429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7439 ( .a ({signal_10429, signal_3975}), .b ({signal_10909, signal_7324}), .c ({signal_11145, signal_7430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7440 ( .a ({signal_10666, signal_7180}), .b ({signal_10910, signal_7325}), .c ({signal_11146, signal_4112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7441 ( .a ({signal_10217, signal_6927}), .b ({signal_10911, signal_7326}), .c ({signal_11147, signal_7431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7442 ( .a ({signal_23652, signal_23644}), .b ({signal_10913, signal_7328}), .c ({signal_11148, signal_7432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7443 ( .a ({signal_23668, signal_23660}), .b ({signal_10914, signal_4211}), .c ({signal_11149, signal_4243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7444 ( .a ({signal_23684, signal_23676}), .b ({signal_10915, signal_7329}), .c ({signal_11150, signal_7433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7445 ( .a ({signal_23700, signal_23692}), .b ({signal_10916, signal_7330}), .c ({signal_11151, signal_7434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7446 ( .a ({signal_23716, signal_23708}), .b ({signal_10917, signal_4214}), .c ({signal_11152, signal_4246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7447 ( .a ({signal_23732, signal_23724}), .b ({signal_10918, signal_4215}), .c ({signal_11153, signal_4247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7448 ( .a ({signal_23748, signal_23740}), .b ({signal_10919, signal_4216}), .c ({signal_11154, signal_4248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7449 ( .a ({signal_23764, signal_23756}), .b ({signal_10920, signal_4195}), .c ({signal_11155, signal_4227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7450 ( .a ({signal_23780, signal_23772}), .b ({signal_10921, signal_7331}), .c ({signal_11156, signal_7435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7451 ( .a ({signal_23796, signal_23788}), .b ({signal_10922, signal_7332}), .c ({signal_11157, signal_7436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7452 ( .a ({signal_23812, signal_23804}), .b ({signal_10923, signal_4198}), .c ({signal_11158, signal_4230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7453 ( .a ({signal_23828, signal_23820}), .b ({signal_10924, signal_7333}), .c ({signal_11159, signal_7437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7454 ( .a ({signal_23844, signal_23836}), .b ({signal_10925, signal_4199}), .c ({signal_11160, signal_4231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7455 ( .a ({signal_23860, signal_23852}), .b ({signal_10926, signal_4200}), .c ({signal_11161, signal_4232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7456 ( .a ({signal_23876, signal_23868}), .b ({signal_10927, signal_7334}), .c ({signal_11162, signal_7438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7457 ( .a ({signal_23892, signal_23884}), .b ({signal_10929, signal_4203}), .c ({signal_11163, signal_4235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7458 ( .a ({signal_23908, signal_23900}), .b ({signal_10930, signal_7336}), .c ({signal_11164, signal_7439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7459 ( .a ({signal_23924, signal_23916}), .b ({signal_10931, signal_7337}), .c ({signal_11165, signal_7440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7460 ( .a ({signal_23940, signal_23932}), .b ({signal_10932, signal_4206}), .c ({signal_11166, signal_4238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7461 ( .a ({signal_23956, signal_23948}), .b ({signal_10933, signal_4207}), .c ({signal_11167, signal_4239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7462 ( .a ({signal_23972, signal_23964}), .b ({signal_10934, signal_4208}), .c ({signal_11168, signal_4240}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7463 ( .a ({signal_11024, signal_7340}), .b ({signal_11276, signal_4018}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7464 ( .a ({signal_11026, signal_7341}), .b ({signal_11277, signal_4020}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7465 ( .a ({signal_11027, signal_7342}), .b ({signal_11278, signal_4021}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7466 ( .a ({signal_11031, signal_7345}), .b ({signal_11279, signal_3996}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7467 ( .a ({signal_11033, signal_7346}), .b ({signal_11280, signal_3997}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7468 ( .a ({signal_11039, signal_7350}), .b ({signal_11281, signal_4004}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7469 ( .a ({signal_11040, signal_7351}), .b ({signal_11282, signal_4005}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7470 ( .a ({signal_11046, signal_7356}), .b ({signal_11283, signal_4010}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7471 ( .a ({signal_11048, signal_7357}), .b ({signal_11284, signal_4012}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7472 ( .a ({signal_11049, signal_7358}), .b ({signal_11285, signal_4013}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7473 ( .a ({signal_11053, signal_7361}), .b ({signal_11286, signal_4026}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7474 ( .a ({signal_11055, signal_7363}), .b ({signal_11287, signal_4050}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7475 ( .a ({signal_11057, signal_7364}), .b ({signal_11288, signal_4052}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7476 ( .a ({signal_11058, signal_7365}), .b ({signal_11289, signal_4053}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7477 ( .a ({signal_11062, signal_7368}), .b ({signal_11290, signal_4028}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7478 ( .a ({signal_11064, signal_7369}), .b ({signal_11291, signal_4029}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7479 ( .a ({signal_11070, signal_7373}), .b ({signal_11292, signal_4036}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7480 ( .a ({signal_11071, signal_7374}), .b ({signal_11293, signal_4037}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7481 ( .a ({signal_11077, signal_7379}), .b ({signal_11294, signal_4042}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7482 ( .a ({signal_11079, signal_7380}), .b ({signal_11295, signal_4044}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7483 ( .a ({signal_11080, signal_7381}), .b ({signal_11296, signal_4045}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7484 ( .a ({signal_11084, signal_7384}), .b ({signal_11297, signal_4058}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7485 ( .a ({signal_11086, signal_7386}), .b ({signal_11298, signal_4082}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7486 ( .a ({signal_11088, signal_7387}), .b ({signal_11299, signal_4084}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7487 ( .a ({signal_11089, signal_7388}), .b ({signal_11300, signal_4085}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7488 ( .a ({signal_11093, signal_7391}), .b ({signal_11301, signal_4060}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7489 ( .a ({signal_11095, signal_7392}), .b ({signal_11302, signal_4061}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7490 ( .a ({signal_11101, signal_7396}), .b ({signal_11303, signal_4068}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7491 ( .a ({signal_11102, signal_7397}), .b ({signal_11304, signal_4069}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7492 ( .a ({signal_11108, signal_7402}), .b ({signal_11305, signal_4074}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7493 ( .a ({signal_11110, signal_7403}), .b ({signal_11306, signal_4076}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7494 ( .a ({signal_11111, signal_7404}), .b ({signal_11307, signal_4077}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7495 ( .a ({signal_11115, signal_7407}), .b ({signal_11308, signal_4090}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7496 ( .a ({signal_11117, signal_7409}), .b ({signal_11309, signal_4114}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7497 ( .a ({signal_11119, signal_7410}), .b ({signal_11310, signal_4116}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7498 ( .a ({signal_11120, signal_7411}), .b ({signal_11311, signal_4117}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7499 ( .a ({signal_11124, signal_7414}), .b ({signal_11312, signal_4092}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7500 ( .a ({signal_11126, signal_7415}), .b ({signal_11313, signal_4093}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7501 ( .a ({signal_11131, signal_7419}), .b ({signal_11314, signal_4098}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7502 ( .a ({signal_11133, signal_7420}), .b ({signal_11315, signal_4100}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7503 ( .a ({signal_11134, signal_7421}), .b ({signal_11316, signal_4101}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7504 ( .a ({signal_11140, signal_7426}), .b ({signal_11317, signal_4106}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7505 ( .a ({signal_11142, signal_7427}), .b ({signal_11318, signal_4108}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7506 ( .a ({signal_11143, signal_7428}), .b ({signal_11319, signal_4109}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7507 ( .a ({signal_11147, signal_7431}), .b ({signal_11320, signal_4122}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7508 ( .a ({signal_11148, signal_7432}), .b ({signal_11321, signal_4241}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7509 ( .a ({signal_11150, signal_7433}), .b ({signal_11322, signal_4244}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7510 ( .a ({signal_11151, signal_7434}), .b ({signal_11323, signal_4245}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7511 ( .a ({signal_11156, signal_7435}), .b ({signal_11324, signal_4228}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7512 ( .a ({signal_11157, signal_7436}), .b ({signal_11325, signal_4229}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7513 ( .a ({signal_11159, signal_7437}), .b ({signal_11326, signal_4249}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7514 ( .a ({signal_11162, signal_7438}), .b ({signal_11327, signal_4233}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7515 ( .a ({signal_11164, signal_7439}), .b ({signal_11328, signal_4236}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7516 ( .a ({signal_11165, signal_7440}), .b ({signal_11329, signal_4237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7517 ( .a ({signal_10410, signal_7034}), .b ({signal_11023, signal_7339}), .c ({signal_11330, signal_7441}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7518 ( .a ({signal_10772, signal_7071}), .b ({signal_11028, signal_7343}), .c ({signal_11331, signal_4022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7519 ( .a ({signal_10773, signal_7072}), .b ({signal_11029, signal_7344}), .c ({signal_11332, signal_4023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7520 ( .a ({signal_10772, signal_7071}), .b ({signal_11034, signal_7347}), .c ({signal_11333, signal_3998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7521 ( .a ({signal_10773, signal_7072}), .b ({signal_11035, signal_7348}), .c ({signal_11334, signal_3999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7522 ( .a ({signal_10775, signal_7078}), .b ({signal_11037, signal_7349}), .c ({signal_11335, signal_7442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7523 ( .a ({signal_10808, signal_7221}), .b ({signal_11041, signal_7352}), .c ({signal_11336, signal_4006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7524 ( .a ({signal_10775, signal_7078}), .b ({signal_11042, signal_7353}), .c ({signal_11337, signal_7443}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7525 ( .a ({signal_10810, signal_7223}), .b ({signal_11043, signal_7354}), .c ({signal_11338, signal_4007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7526 ( .a ({signal_10812, signal_7225}), .b ({signal_11045, signal_7355}), .c ({signal_11339, signal_7444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7527 ( .a ({signal_10818, signal_7231}), .b ({signal_11050, signal_7359}), .c ({signal_11340, signal_4014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7528 ( .a ({signal_10820, signal_7233}), .b ({signal_11051, signal_7360}), .c ({signal_11341, signal_4015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7529 ( .a ({signal_10389, signal_7025}), .b ({signal_11054, signal_7362}), .c ({signal_11342, signal_7445}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7530 ( .a ({signal_10776, signal_7103}), .b ({signal_11059, signal_7366}), .c ({signal_11343, signal_4054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7531 ( .a ({signal_10777, signal_7104}), .b ({signal_11060, signal_7367}), .c ({signal_11344, signal_4055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7532 ( .a ({signal_10776, signal_7103}), .b ({signal_11065, signal_7370}), .c ({signal_11345, signal_4030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7533 ( .a ({signal_10777, signal_7104}), .b ({signal_11066, signal_7371}), .c ({signal_11346, signal_4031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7534 ( .a ({signal_10779, signal_7110}), .b ({signal_11068, signal_7372}), .c ({signal_11347, signal_7446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7535 ( .a ({signal_10836, signal_7250}), .b ({signal_11072, signal_7375}), .c ({signal_11348, signal_4038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7536 ( .a ({signal_10779, signal_7110}), .b ({signal_11073, signal_7376}), .c ({signal_11349, signal_7447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7537 ( .a ({signal_10838, signal_7252}), .b ({signal_11074, signal_7377}), .c ({signal_11350, signal_4039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7538 ( .a ({signal_10840, signal_7254}), .b ({signal_11076, signal_7378}), .c ({signal_11351, signal_7448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7539 ( .a ({signal_10846, signal_7260}), .b ({signal_11081, signal_7382}), .c ({signal_11352, signal_4046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7540 ( .a ({signal_10848, signal_7262}), .b ({signal_11082, signal_7383}), .c ({signal_11353, signal_4047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7541 ( .a ({signal_10361, signal_7013}), .b ({signal_11085, signal_7385}), .c ({signal_11354, signal_7449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7542 ( .a ({signal_10780, signal_7135}), .b ({signal_11090, signal_7389}), .c ({signal_11355, signal_4086}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7543 ( .a ({signal_10781, signal_7136}), .b ({signal_11091, signal_7390}), .c ({signal_11356, signal_4087}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7544 ( .a ({signal_10780, signal_7135}), .b ({signal_11096, signal_7393}), .c ({signal_11357, signal_4062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7545 ( .a ({signal_10781, signal_7136}), .b ({signal_11097, signal_7394}), .c ({signal_11358, signal_4063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7546 ( .a ({signal_10783, signal_7142}), .b ({signal_11099, signal_7395}), .c ({signal_11359, signal_7450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7547 ( .a ({signal_10864, signal_7279}), .b ({signal_11103, signal_7398}), .c ({signal_11360, signal_4070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7548 ( .a ({signal_10783, signal_7142}), .b ({signal_11104, signal_7399}), .c ({signal_11361, signal_7451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7549 ( .a ({signal_10866, signal_7281}), .b ({signal_11105, signal_7400}), .c ({signal_11362, signal_4071}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7550 ( .a ({signal_10868, signal_7283}), .b ({signal_11107, signal_7401}), .c ({signal_11363, signal_7452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7551 ( .a ({signal_10874, signal_7289}), .b ({signal_11112, signal_7405}), .c ({signal_11364, signal_4078}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7552 ( .a ({signal_10876, signal_7291}), .b ({signal_11113, signal_7406}), .c ({signal_11365, signal_4079}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7553 ( .a ({signal_10431, signal_7043}), .b ({signal_11116, signal_7408}), .c ({signal_11366, signal_7453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7554 ( .a ({signal_10888, signal_7303}), .b ({signal_11121, signal_7412}), .c ({signal_11367, signal_4118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7555 ( .a ({signal_10889, signal_7304}), .b ({signal_11122, signal_7413}), .c ({signal_11368, signal_4119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7556 ( .a ({signal_10888, signal_7303}), .b ({signal_11127, signal_7416}), .c ({signal_11369, signal_4094}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7557 ( .a ({signal_10889, signal_7304}), .b ({signal_11128, signal_7417}), .c ({signal_11370, signal_4095}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7558 ( .a ({signal_10896, signal_7311}), .b ({signal_11130, signal_7418}), .c ({signal_11371, signal_7454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7559 ( .a ({signal_10895, signal_7310}), .b ({signal_11135, signal_7422}), .c ({signal_11372, signal_4102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7560 ( .a ({signal_10896, signal_7311}), .b ({signal_11136, signal_7423}), .c ({signal_11373, signal_7455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7561 ( .a ({signal_10898, signal_7313}), .b ({signal_11137, signal_7424}), .c ({signal_11374, signal_4103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7562 ( .a ({signal_10900, signal_7315}), .b ({signal_11139, signal_7425}), .c ({signal_11375, signal_7456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7563 ( .a ({signal_10906, signal_7321}), .b ({signal_11144, signal_7429}), .c ({signal_11376, signal_4110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7564 ( .a ({signal_10908, signal_7323}), .b ({signal_11145, signal_7430}), .c ({signal_11377, signal_4111}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7565 ( .a ({signal_11330, signal_7441}), .b ({signal_11559, signal_4017}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7566 ( .a ({signal_11335, signal_7442}), .b ({signal_11560, signal_4001}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7567 ( .a ({signal_11337, signal_7443}), .b ({signal_11561, signal_4025}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7568 ( .a ({signal_11339, signal_7444}), .b ({signal_11562, signal_4009}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7569 ( .a ({signal_11342, signal_7445}), .b ({signal_11563, signal_4049}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7570 ( .a ({signal_11347, signal_7446}), .b ({signal_11564, signal_4033}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7571 ( .a ({signal_11349, signal_7447}), .b ({signal_11565, signal_4057}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7572 ( .a ({signal_11351, signal_7448}), .b ({signal_11566, signal_4041}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7573 ( .a ({signal_11354, signal_7449}), .b ({signal_11567, signal_4081}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7574 ( .a ({signal_11359, signal_7450}), .b ({signal_11568, signal_4065}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7575 ( .a ({signal_11361, signal_7451}), .b ({signal_11569, signal_4089}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7576 ( .a ({signal_11363, signal_7452}), .b ({signal_11570, signal_4073}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7577 ( .a ({signal_11366, signal_7453}), .b ({signal_11571, signal_4113}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7578 ( .a ({signal_11371, signal_7454}), .b ({signal_11572, signal_4097}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7579 ( .a ({signal_11373, signal_7455}), .b ({signal_11573, signal_4121}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_7580 ( .a ({signal_11375, signal_7456}), .b ({signal_11574, signal_4105}) ) ;
    buf_clk cell_8548 ( .C (clk), .D (signal_13435), .Q (signal_13436) ) ;
    buf_clk cell_8556 ( .C (clk), .D (signal_13443), .Q (signal_13444) ) ;
    buf_clk cell_8564 ( .C (clk), .D (signal_13451), .Q (signal_13452) ) ;
    buf_clk cell_8572 ( .C (clk), .D (signal_13459), .Q (signal_13460) ) ;
    buf_clk cell_8580 ( .C (clk), .D (signal_13467), .Q (signal_13468) ) ;
    buf_clk cell_8588 ( .C (clk), .D (signal_13475), .Q (signal_13476) ) ;
    buf_clk cell_8596 ( .C (clk), .D (signal_13483), .Q (signal_13484) ) ;
    buf_clk cell_8604 ( .C (clk), .D (signal_13491), .Q (signal_13492) ) ;
    buf_clk cell_8612 ( .C (clk), .D (signal_13499), .Q (signal_13500) ) ;
    buf_clk cell_8620 ( .C (clk), .D (signal_13507), .Q (signal_13508) ) ;
    buf_clk cell_8628 ( .C (clk), .D (signal_13515), .Q (signal_13516) ) ;
    buf_clk cell_8636 ( .C (clk), .D (signal_13523), .Q (signal_13524) ) ;
    buf_clk cell_8644 ( .C (clk), .D (signal_13531), .Q (signal_13532) ) ;
    buf_clk cell_8652 ( .C (clk), .D (signal_13539), .Q (signal_13540) ) ;
    buf_clk cell_8660 ( .C (clk), .D (signal_13547), .Q (signal_13548) ) ;
    buf_clk cell_8668 ( .C (clk), .D (signal_13555), .Q (signal_13556) ) ;
    buf_clk cell_8676 ( .C (clk), .D (signal_13563), .Q (signal_13564) ) ;
    buf_clk cell_8684 ( .C (clk), .D (signal_13571), .Q (signal_13572) ) ;
    buf_clk cell_8692 ( .C (clk), .D (signal_13579), .Q (signal_13580) ) ;
    buf_clk cell_8700 ( .C (clk), .D (signal_13587), .Q (signal_13588) ) ;
    buf_clk cell_8708 ( .C (clk), .D (signal_13595), .Q (signal_13596) ) ;
    buf_clk cell_8716 ( .C (clk), .D (signal_13603), .Q (signal_13604) ) ;
    buf_clk cell_8724 ( .C (clk), .D (signal_13611), .Q (signal_13612) ) ;
    buf_clk cell_8732 ( .C (clk), .D (signal_13619), .Q (signal_13620) ) ;
    buf_clk cell_8740 ( .C (clk), .D (signal_13627), .Q (signal_13628) ) ;
    buf_clk cell_8748 ( .C (clk), .D (signal_13635), .Q (signal_13636) ) ;
    buf_clk cell_8756 ( .C (clk), .D (signal_13643), .Q (signal_13644) ) ;
    buf_clk cell_8764 ( .C (clk), .D (signal_13651), .Q (signal_13652) ) ;
    buf_clk cell_8772 ( .C (clk), .D (signal_13659), .Q (signal_13660) ) ;
    buf_clk cell_8780 ( .C (clk), .D (signal_13667), .Q (signal_13668) ) ;
    buf_clk cell_8788 ( .C (clk), .D (signal_13675), .Q (signal_13676) ) ;
    buf_clk cell_8796 ( .C (clk), .D (signal_13683), .Q (signal_13684) ) ;
    buf_clk cell_8804 ( .C (clk), .D (signal_13691), .Q (signal_13692) ) ;
    buf_clk cell_8812 ( .C (clk), .D (signal_13699), .Q (signal_13700) ) ;
    buf_clk cell_8820 ( .C (clk), .D (signal_13707), .Q (signal_13708) ) ;
    buf_clk cell_8828 ( .C (clk), .D (signal_13715), .Q (signal_13716) ) ;
    buf_clk cell_8836 ( .C (clk), .D (signal_13723), .Q (signal_13724) ) ;
    buf_clk cell_8844 ( .C (clk), .D (signal_13731), .Q (signal_13732) ) ;
    buf_clk cell_8852 ( .C (clk), .D (signal_13739), .Q (signal_13740) ) ;
    buf_clk cell_8860 ( .C (clk), .D (signal_13747), .Q (signal_13748) ) ;
    buf_clk cell_8868 ( .C (clk), .D (signal_13755), .Q (signal_13756) ) ;
    buf_clk cell_8876 ( .C (clk), .D (signal_13763), .Q (signal_13764) ) ;
    buf_clk cell_8884 ( .C (clk), .D (signal_13771), .Q (signal_13772) ) ;
    buf_clk cell_8892 ( .C (clk), .D (signal_13779), .Q (signal_13780) ) ;
    buf_clk cell_8900 ( .C (clk), .D (signal_13787), .Q (signal_13788) ) ;
    buf_clk cell_8908 ( .C (clk), .D (signal_13795), .Q (signal_13796) ) ;
    buf_clk cell_8916 ( .C (clk), .D (signal_13803), .Q (signal_13804) ) ;
    buf_clk cell_8924 ( .C (clk), .D (signal_13811), .Q (signal_13812) ) ;
    buf_clk cell_8932 ( .C (clk), .D (signal_13819), .Q (signal_13820) ) ;
    buf_clk cell_8940 ( .C (clk), .D (signal_13827), .Q (signal_13828) ) ;
    buf_clk cell_8948 ( .C (clk), .D (signal_13835), .Q (signal_13836) ) ;
    buf_clk cell_8956 ( .C (clk), .D (signal_13843), .Q (signal_13844) ) ;
    buf_clk cell_8964 ( .C (clk), .D (signal_13851), .Q (signal_13852) ) ;
    buf_clk cell_8972 ( .C (clk), .D (signal_13859), .Q (signal_13860) ) ;
    buf_clk cell_8980 ( .C (clk), .D (signal_13867), .Q (signal_13868) ) ;
    buf_clk cell_8988 ( .C (clk), .D (signal_13875), .Q (signal_13876) ) ;
    buf_clk cell_8996 ( .C (clk), .D (signal_13883), .Q (signal_13884) ) ;
    buf_clk cell_9004 ( .C (clk), .D (signal_13891), .Q (signal_13892) ) ;
    buf_clk cell_9012 ( .C (clk), .D (signal_13899), .Q (signal_13900) ) ;
    buf_clk cell_9020 ( .C (clk), .D (signal_13907), .Q (signal_13908) ) ;
    buf_clk cell_9028 ( .C (clk), .D (signal_13915), .Q (signal_13916) ) ;
    buf_clk cell_9036 ( .C (clk), .D (signal_13923), .Q (signal_13924) ) ;
    buf_clk cell_9044 ( .C (clk), .D (signal_13931), .Q (signal_13932) ) ;
    buf_clk cell_9052 ( .C (clk), .D (signal_13939), .Q (signal_13940) ) ;
    buf_clk cell_9060 ( .C (clk), .D (signal_13947), .Q (signal_13948) ) ;
    buf_clk cell_9068 ( .C (clk), .D (signal_13955), .Q (signal_13956) ) ;
    buf_clk cell_9076 ( .C (clk), .D (signal_13963), .Q (signal_13964) ) ;
    buf_clk cell_9084 ( .C (clk), .D (signal_13971), .Q (signal_13972) ) ;
    buf_clk cell_9092 ( .C (clk), .D (signal_13979), .Q (signal_13980) ) ;
    buf_clk cell_9100 ( .C (clk), .D (signal_13987), .Q (signal_13988) ) ;
    buf_clk cell_9108 ( .C (clk), .D (signal_13995), .Q (signal_13996) ) ;
    buf_clk cell_9116 ( .C (clk), .D (signal_14003), .Q (signal_14004) ) ;
    buf_clk cell_9124 ( .C (clk), .D (signal_14011), .Q (signal_14012) ) ;
    buf_clk cell_9132 ( .C (clk), .D (signal_14019), .Q (signal_14020) ) ;
    buf_clk cell_9140 ( .C (clk), .D (signal_14027), .Q (signal_14028) ) ;
    buf_clk cell_9148 ( .C (clk), .D (signal_14035), .Q (signal_14036) ) ;
    buf_clk cell_9156 ( .C (clk), .D (signal_14043), .Q (signal_14044) ) ;
    buf_clk cell_9164 ( .C (clk), .D (signal_14051), .Q (signal_14052) ) ;
    buf_clk cell_9172 ( .C (clk), .D (signal_14059), .Q (signal_14060) ) ;
    buf_clk cell_9180 ( .C (clk), .D (signal_14067), .Q (signal_14068) ) ;
    buf_clk cell_9188 ( .C (clk), .D (signal_14075), .Q (signal_14076) ) ;
    buf_clk cell_9196 ( .C (clk), .D (signal_14083), .Q (signal_14084) ) ;
    buf_clk cell_9204 ( .C (clk), .D (signal_14091), .Q (signal_14092) ) ;
    buf_clk cell_9212 ( .C (clk), .D (signal_14099), .Q (signal_14100) ) ;
    buf_clk cell_9220 ( .C (clk), .D (signal_14107), .Q (signal_14108) ) ;
    buf_clk cell_9228 ( .C (clk), .D (signal_14115), .Q (signal_14116) ) ;
    buf_clk cell_9236 ( .C (clk), .D (signal_14123), .Q (signal_14124) ) ;
    buf_clk cell_9244 ( .C (clk), .D (signal_14131), .Q (signal_14132) ) ;
    buf_clk cell_9252 ( .C (clk), .D (signal_14139), .Q (signal_14140) ) ;
    buf_clk cell_9260 ( .C (clk), .D (signal_14147), .Q (signal_14148) ) ;
    buf_clk cell_9268 ( .C (clk), .D (signal_14155), .Q (signal_14156) ) ;
    buf_clk cell_9276 ( .C (clk), .D (signal_14163), .Q (signal_14164) ) ;
    buf_clk cell_9284 ( .C (clk), .D (signal_14171), .Q (signal_14172) ) ;
    buf_clk cell_9292 ( .C (clk), .D (signal_14179), .Q (signal_14180) ) ;
    buf_clk cell_9300 ( .C (clk), .D (signal_14187), .Q (signal_14188) ) ;
    buf_clk cell_9308 ( .C (clk), .D (signal_14195), .Q (signal_14196) ) ;
    buf_clk cell_9316 ( .C (clk), .D (signal_14203), .Q (signal_14204) ) ;
    buf_clk cell_9324 ( .C (clk), .D (signal_14211), .Q (signal_14212) ) ;
    buf_clk cell_9332 ( .C (clk), .D (signal_14219), .Q (signal_14220) ) ;
    buf_clk cell_9340 ( .C (clk), .D (signal_14227), .Q (signal_14228) ) ;
    buf_clk cell_9348 ( .C (clk), .D (signal_14235), .Q (signal_14236) ) ;
    buf_clk cell_9356 ( .C (clk), .D (signal_14243), .Q (signal_14244) ) ;
    buf_clk cell_9364 ( .C (clk), .D (signal_14251), .Q (signal_14252) ) ;
    buf_clk cell_9372 ( .C (clk), .D (signal_14259), .Q (signal_14260) ) ;
    buf_clk cell_9380 ( .C (clk), .D (signal_14267), .Q (signal_14268) ) ;
    buf_clk cell_9388 ( .C (clk), .D (signal_14275), .Q (signal_14276) ) ;
    buf_clk cell_9396 ( .C (clk), .D (signal_14283), .Q (signal_14284) ) ;
    buf_clk cell_9404 ( .C (clk), .D (signal_14291), .Q (signal_14292) ) ;
    buf_clk cell_9412 ( .C (clk), .D (signal_14299), .Q (signal_14300) ) ;
    buf_clk cell_9420 ( .C (clk), .D (signal_14307), .Q (signal_14308) ) ;
    buf_clk cell_9428 ( .C (clk), .D (signal_14315), .Q (signal_14316) ) ;
    buf_clk cell_9436 ( .C (clk), .D (signal_14323), .Q (signal_14324) ) ;
    buf_clk cell_9444 ( .C (clk), .D (signal_14331), .Q (signal_14332) ) ;
    buf_clk cell_9452 ( .C (clk), .D (signal_14339), .Q (signal_14340) ) ;
    buf_clk cell_9460 ( .C (clk), .D (signal_14347), .Q (signal_14348) ) ;
    buf_clk cell_9468 ( .C (clk), .D (signal_14355), .Q (signal_14356) ) ;
    buf_clk cell_9476 ( .C (clk), .D (signal_14363), .Q (signal_14364) ) ;
    buf_clk cell_9484 ( .C (clk), .D (signal_14371), .Q (signal_14372) ) ;
    buf_clk cell_9492 ( .C (clk), .D (signal_14379), .Q (signal_14380) ) ;
    buf_clk cell_9500 ( .C (clk), .D (signal_14387), .Q (signal_14388) ) ;
    buf_clk cell_9508 ( .C (clk), .D (signal_14395), .Q (signal_14396) ) ;
    buf_clk cell_9516 ( .C (clk), .D (signal_14403), .Q (signal_14404) ) ;
    buf_clk cell_9524 ( .C (clk), .D (signal_14411), .Q (signal_14412) ) ;
    buf_clk cell_9532 ( .C (clk), .D (signal_14419), .Q (signal_14420) ) ;
    buf_clk cell_9540 ( .C (clk), .D (signal_14427), .Q (signal_14428) ) ;
    buf_clk cell_9548 ( .C (clk), .D (signal_14435), .Q (signal_14436) ) ;
    buf_clk cell_9556 ( .C (clk), .D (signal_14443), .Q (signal_14444) ) ;
    buf_clk cell_9564 ( .C (clk), .D (signal_14451), .Q (signal_14452) ) ;
    buf_clk cell_9572 ( .C (clk), .D (signal_14459), .Q (signal_14460) ) ;
    buf_clk cell_9580 ( .C (clk), .D (signal_14467), .Q (signal_14468) ) ;
    buf_clk cell_9588 ( .C (clk), .D (signal_14475), .Q (signal_14476) ) ;
    buf_clk cell_9596 ( .C (clk), .D (signal_14483), .Q (signal_14484) ) ;
    buf_clk cell_9604 ( .C (clk), .D (signal_14491), .Q (signal_14492) ) ;
    buf_clk cell_9612 ( .C (clk), .D (signal_14499), .Q (signal_14500) ) ;
    buf_clk cell_9620 ( .C (clk), .D (signal_14507), .Q (signal_14508) ) ;
    buf_clk cell_9628 ( .C (clk), .D (signal_14515), .Q (signal_14516) ) ;
    buf_clk cell_9636 ( .C (clk), .D (signal_14523), .Q (signal_14524) ) ;
    buf_clk cell_9644 ( .C (clk), .D (signal_14531), .Q (signal_14532) ) ;
    buf_clk cell_9652 ( .C (clk), .D (signal_14539), .Q (signal_14540) ) ;
    buf_clk cell_9660 ( .C (clk), .D (signal_14547), .Q (signal_14548) ) ;
    buf_clk cell_9668 ( .C (clk), .D (signal_14555), .Q (signal_14556) ) ;
    buf_clk cell_9676 ( .C (clk), .D (signal_14563), .Q (signal_14564) ) ;
    buf_clk cell_9684 ( .C (clk), .D (signal_14571), .Q (signal_14572) ) ;
    buf_clk cell_9692 ( .C (clk), .D (signal_14579), .Q (signal_14580) ) ;
    buf_clk cell_9700 ( .C (clk), .D (signal_14587), .Q (signal_14588) ) ;
    buf_clk cell_9708 ( .C (clk), .D (signal_14595), .Q (signal_14596) ) ;
    buf_clk cell_9716 ( .C (clk), .D (signal_14603), .Q (signal_14604) ) ;
    buf_clk cell_9724 ( .C (clk), .D (signal_14611), .Q (signal_14612) ) ;
    buf_clk cell_9732 ( .C (clk), .D (signal_14619), .Q (signal_14620) ) ;
    buf_clk cell_9740 ( .C (clk), .D (signal_14627), .Q (signal_14628) ) ;
    buf_clk cell_9748 ( .C (clk), .D (signal_14635), .Q (signal_14636) ) ;
    buf_clk cell_9756 ( .C (clk), .D (signal_14643), .Q (signal_14644) ) ;
    buf_clk cell_9764 ( .C (clk), .D (signal_14651), .Q (signal_14652) ) ;
    buf_clk cell_9772 ( .C (clk), .D (signal_14659), .Q (signal_14660) ) ;
    buf_clk cell_9780 ( .C (clk), .D (signal_14667), .Q (signal_14668) ) ;
    buf_clk cell_9788 ( .C (clk), .D (signal_14675), .Q (signal_14676) ) ;
    buf_clk cell_9796 ( .C (clk), .D (signal_14683), .Q (signal_14684) ) ;
    buf_clk cell_9804 ( .C (clk), .D (signal_14691), .Q (signal_14692) ) ;
    buf_clk cell_9812 ( .C (clk), .D (signal_14699), .Q (signal_14700) ) ;
    buf_clk cell_9820 ( .C (clk), .D (signal_14707), .Q (signal_14708) ) ;
    buf_clk cell_9828 ( .C (clk), .D (signal_14715), .Q (signal_14716) ) ;
    buf_clk cell_9836 ( .C (clk), .D (signal_14723), .Q (signal_14724) ) ;
    buf_clk cell_9844 ( .C (clk), .D (signal_14731), .Q (signal_14732) ) ;
    buf_clk cell_9852 ( .C (clk), .D (signal_14739), .Q (signal_14740) ) ;
    buf_clk cell_9860 ( .C (clk), .D (signal_14747), .Q (signal_14748) ) ;
    buf_clk cell_9868 ( .C (clk), .D (signal_14755), .Q (signal_14756) ) ;
    buf_clk cell_9876 ( .C (clk), .D (signal_14763), .Q (signal_14764) ) ;
    buf_clk cell_9884 ( .C (clk), .D (signal_14771), .Q (signal_14772) ) ;
    buf_clk cell_9892 ( .C (clk), .D (signal_14779), .Q (signal_14780) ) ;
    buf_clk cell_9900 ( .C (clk), .D (signal_14787), .Q (signal_14788) ) ;
    buf_clk cell_9908 ( .C (clk), .D (signal_14795), .Q (signal_14796) ) ;
    buf_clk cell_9916 ( .C (clk), .D (signal_14803), .Q (signal_14804) ) ;
    buf_clk cell_9924 ( .C (clk), .D (signal_14811), .Q (signal_14812) ) ;
    buf_clk cell_9932 ( .C (clk), .D (signal_14819), .Q (signal_14820) ) ;
    buf_clk cell_9940 ( .C (clk), .D (signal_14827), .Q (signal_14828) ) ;
    buf_clk cell_9948 ( .C (clk), .D (signal_14835), .Q (signal_14836) ) ;
    buf_clk cell_9956 ( .C (clk), .D (signal_14843), .Q (signal_14844) ) ;
    buf_clk cell_9964 ( .C (clk), .D (signal_14851), .Q (signal_14852) ) ;
    buf_clk cell_9972 ( .C (clk), .D (signal_14859), .Q (signal_14860) ) ;
    buf_clk cell_9980 ( .C (clk), .D (signal_14867), .Q (signal_14868) ) ;
    buf_clk cell_9988 ( .C (clk), .D (signal_14875), .Q (signal_14876) ) ;
    buf_clk cell_9996 ( .C (clk), .D (signal_14883), .Q (signal_14884) ) ;
    buf_clk cell_10004 ( .C (clk), .D (signal_14891), .Q (signal_14892) ) ;
    buf_clk cell_10012 ( .C (clk), .D (signal_14899), .Q (signal_14900) ) ;
    buf_clk cell_10020 ( .C (clk), .D (signal_14907), .Q (signal_14908) ) ;
    buf_clk cell_10028 ( .C (clk), .D (signal_14915), .Q (signal_14916) ) ;
    buf_clk cell_10036 ( .C (clk), .D (signal_14923), .Q (signal_14924) ) ;
    buf_clk cell_10044 ( .C (clk), .D (signal_14931), .Q (signal_14932) ) ;
    buf_clk cell_10052 ( .C (clk), .D (signal_14939), .Q (signal_14940) ) ;
    buf_clk cell_10060 ( .C (clk), .D (signal_14947), .Q (signal_14948) ) ;
    buf_clk cell_10068 ( .C (clk), .D (signal_14955), .Q (signal_14956) ) ;
    buf_clk cell_10076 ( .C (clk), .D (signal_14963), .Q (signal_14964) ) ;
    buf_clk cell_10084 ( .C (clk), .D (signal_14971), .Q (signal_14972) ) ;
    buf_clk cell_10092 ( .C (clk), .D (signal_14979), .Q (signal_14980) ) ;
    buf_clk cell_10100 ( .C (clk), .D (signal_14987), .Q (signal_14988) ) ;
    buf_clk cell_10108 ( .C (clk), .D (signal_14995), .Q (signal_14996) ) ;
    buf_clk cell_10116 ( .C (clk), .D (signal_15003), .Q (signal_15004) ) ;
    buf_clk cell_10124 ( .C (clk), .D (signal_15011), .Q (signal_15012) ) ;
    buf_clk cell_10132 ( .C (clk), .D (signal_15019), .Q (signal_15020) ) ;
    buf_clk cell_10140 ( .C (clk), .D (signal_15027), .Q (signal_15028) ) ;
    buf_clk cell_10148 ( .C (clk), .D (signal_15035), .Q (signal_15036) ) ;
    buf_clk cell_10156 ( .C (clk), .D (signal_15043), .Q (signal_15044) ) ;
    buf_clk cell_10164 ( .C (clk), .D (signal_15051), .Q (signal_15052) ) ;
    buf_clk cell_10172 ( .C (clk), .D (signal_15059), .Q (signal_15060) ) ;
    buf_clk cell_10180 ( .C (clk), .D (signal_15067), .Q (signal_15068) ) ;
    buf_clk cell_10188 ( .C (clk), .D (signal_15075), .Q (signal_15076) ) ;
    buf_clk cell_10196 ( .C (clk), .D (signal_15083), .Q (signal_15084) ) ;
    buf_clk cell_10204 ( .C (clk), .D (signal_15091), .Q (signal_15092) ) ;
    buf_clk cell_10212 ( .C (clk), .D (signal_15099), .Q (signal_15100) ) ;
    buf_clk cell_10220 ( .C (clk), .D (signal_15107), .Q (signal_15108) ) ;
    buf_clk cell_10228 ( .C (clk), .D (signal_15115), .Q (signal_15116) ) ;
    buf_clk cell_10236 ( .C (clk), .D (signal_15123), .Q (signal_15124) ) ;
    buf_clk cell_10244 ( .C (clk), .D (signal_15131), .Q (signal_15132) ) ;
    buf_clk cell_10252 ( .C (clk), .D (signal_15139), .Q (signal_15140) ) ;
    buf_clk cell_10260 ( .C (clk), .D (signal_15147), .Q (signal_15148) ) ;
    buf_clk cell_10268 ( .C (clk), .D (signal_15155), .Q (signal_15156) ) ;
    buf_clk cell_10276 ( .C (clk), .D (signal_15163), .Q (signal_15164) ) ;
    buf_clk cell_10284 ( .C (clk), .D (signal_15171), .Q (signal_15172) ) ;
    buf_clk cell_10292 ( .C (clk), .D (signal_15179), .Q (signal_15180) ) ;
    buf_clk cell_10300 ( .C (clk), .D (signal_15187), .Q (signal_15188) ) ;
    buf_clk cell_10308 ( .C (clk), .D (signal_15195), .Q (signal_15196) ) ;
    buf_clk cell_10316 ( .C (clk), .D (signal_15203), .Q (signal_15204) ) ;
    buf_clk cell_10324 ( .C (clk), .D (signal_15211), .Q (signal_15212) ) ;
    buf_clk cell_10332 ( .C (clk), .D (signal_15219), .Q (signal_15220) ) ;
    buf_clk cell_10340 ( .C (clk), .D (signal_15227), .Q (signal_15228) ) ;
    buf_clk cell_10348 ( .C (clk), .D (signal_15235), .Q (signal_15236) ) ;
    buf_clk cell_10356 ( .C (clk), .D (signal_15243), .Q (signal_15244) ) ;
    buf_clk cell_10364 ( .C (clk), .D (signal_15251), .Q (signal_15252) ) ;
    buf_clk cell_10372 ( .C (clk), .D (signal_15259), .Q (signal_15260) ) ;
    buf_clk cell_10380 ( .C (clk), .D (signal_15267), .Q (signal_15268) ) ;
    buf_clk cell_10388 ( .C (clk), .D (signal_15275), .Q (signal_15276) ) ;
    buf_clk cell_10396 ( .C (clk), .D (signal_15283), .Q (signal_15284) ) ;
    buf_clk cell_10404 ( .C (clk), .D (signal_15291), .Q (signal_15292) ) ;
    buf_clk cell_10412 ( .C (clk), .D (signal_15299), .Q (signal_15300) ) ;
    buf_clk cell_10420 ( .C (clk), .D (signal_15307), .Q (signal_15308) ) ;
    buf_clk cell_10428 ( .C (clk), .D (signal_15315), .Q (signal_15316) ) ;
    buf_clk cell_10436 ( .C (clk), .D (signal_15323), .Q (signal_15324) ) ;
    buf_clk cell_10444 ( .C (clk), .D (signal_15331), .Q (signal_15332) ) ;
    buf_clk cell_10452 ( .C (clk), .D (signal_15339), .Q (signal_15340) ) ;
    buf_clk cell_10460 ( .C (clk), .D (signal_15347), .Q (signal_15348) ) ;
    buf_clk cell_10468 ( .C (clk), .D (signal_15355), .Q (signal_15356) ) ;
    buf_clk cell_10476 ( .C (clk), .D (signal_15363), .Q (signal_15364) ) ;
    buf_clk cell_10484 ( .C (clk), .D (signal_15371), .Q (signal_15372) ) ;
    buf_clk cell_10492 ( .C (clk), .D (signal_15379), .Q (signal_15380) ) ;
    buf_clk cell_10500 ( .C (clk), .D (signal_15387), .Q (signal_15388) ) ;
    buf_clk cell_10508 ( .C (clk), .D (signal_15395), .Q (signal_15396) ) ;
    buf_clk cell_10516 ( .C (clk), .D (signal_15403), .Q (signal_15404) ) ;
    buf_clk cell_10524 ( .C (clk), .D (signal_15411), .Q (signal_15412) ) ;
    buf_clk cell_10532 ( .C (clk), .D (signal_15419), .Q (signal_15420) ) ;
    buf_clk cell_10540 ( .C (clk), .D (signal_15427), .Q (signal_15428) ) ;
    buf_clk cell_10548 ( .C (clk), .D (signal_15435), .Q (signal_15436) ) ;
    buf_clk cell_10556 ( .C (clk), .D (signal_15443), .Q (signal_15444) ) ;
    buf_clk cell_10564 ( .C (clk), .D (signal_15451), .Q (signal_15452) ) ;
    buf_clk cell_10572 ( .C (clk), .D (signal_15459), .Q (signal_15460) ) ;
    buf_clk cell_10580 ( .C (clk), .D (signal_15467), .Q (signal_15468) ) ;
    buf_clk cell_10588 ( .C (clk), .D (signal_15475), .Q (signal_15476) ) ;
    buf_clk cell_10596 ( .C (clk), .D (signal_15483), .Q (signal_15484) ) ;
    buf_clk cell_10604 ( .C (clk), .D (signal_15491), .Q (signal_15492) ) ;
    buf_clk cell_10612 ( .C (clk), .D (signal_15499), .Q (signal_15500) ) ;
    buf_clk cell_10620 ( .C (clk), .D (signal_15507), .Q (signal_15508) ) ;
    buf_clk cell_10628 ( .C (clk), .D (signal_15515), .Q (signal_15516) ) ;
    buf_clk cell_10636 ( .C (clk), .D (signal_15523), .Q (signal_15524) ) ;
    buf_clk cell_10644 ( .C (clk), .D (signal_15531), .Q (signal_15532) ) ;
    buf_clk cell_10652 ( .C (clk), .D (signal_15539), .Q (signal_15540) ) ;
    buf_clk cell_10660 ( .C (clk), .D (signal_15547), .Q (signal_15548) ) ;
    buf_clk cell_10668 ( .C (clk), .D (signal_15555), .Q (signal_15556) ) ;
    buf_clk cell_10676 ( .C (clk), .D (signal_15563), .Q (signal_15564) ) ;
    buf_clk cell_10684 ( .C (clk), .D (signal_15571), .Q (signal_15572) ) ;
    buf_clk cell_10692 ( .C (clk), .D (signal_15579), .Q (signal_15580) ) ;
    buf_clk cell_10700 ( .C (clk), .D (signal_15587), .Q (signal_15588) ) ;
    buf_clk cell_10708 ( .C (clk), .D (signal_15595), .Q (signal_15596) ) ;
    buf_clk cell_10716 ( .C (clk), .D (signal_15603), .Q (signal_15604) ) ;
    buf_clk cell_10724 ( .C (clk), .D (signal_15611), .Q (signal_15612) ) ;
    buf_clk cell_10732 ( .C (clk), .D (signal_15619), .Q (signal_15620) ) ;
    buf_clk cell_10740 ( .C (clk), .D (signal_15627), .Q (signal_15628) ) ;
    buf_clk cell_10748 ( .C (clk), .D (signal_15635), .Q (signal_15636) ) ;
    buf_clk cell_10756 ( .C (clk), .D (signal_15643), .Q (signal_15644) ) ;
    buf_clk cell_10764 ( .C (clk), .D (signal_15651), .Q (signal_15652) ) ;
    buf_clk cell_10772 ( .C (clk), .D (signal_15659), .Q (signal_15660) ) ;
    buf_clk cell_10780 ( .C (clk), .D (signal_15667), .Q (signal_15668) ) ;
    buf_clk cell_10788 ( .C (clk), .D (signal_15675), .Q (signal_15676) ) ;
    buf_clk cell_10796 ( .C (clk), .D (signal_15683), .Q (signal_15684) ) ;
    buf_clk cell_10804 ( .C (clk), .D (signal_15691), .Q (signal_15692) ) ;
    buf_clk cell_10812 ( .C (clk), .D (signal_15699), .Q (signal_15700) ) ;
    buf_clk cell_10820 ( .C (clk), .D (signal_15707), .Q (signal_15708) ) ;
    buf_clk cell_10828 ( .C (clk), .D (signal_15715), .Q (signal_15716) ) ;
    buf_clk cell_10836 ( .C (clk), .D (signal_15723), .Q (signal_15724) ) ;
    buf_clk cell_10844 ( .C (clk), .D (signal_15731), .Q (signal_15732) ) ;
    buf_clk cell_10852 ( .C (clk), .D (signal_15739), .Q (signal_15740) ) ;
    buf_clk cell_10860 ( .C (clk), .D (signal_15747), .Q (signal_15748) ) ;
    buf_clk cell_10868 ( .C (clk), .D (signal_15755), .Q (signal_15756) ) ;
    buf_clk cell_10876 ( .C (clk), .D (signal_15763), .Q (signal_15764) ) ;
    buf_clk cell_10884 ( .C (clk), .D (signal_15771), .Q (signal_15772) ) ;
    buf_clk cell_10892 ( .C (clk), .D (signal_15779), .Q (signal_15780) ) ;
    buf_clk cell_10900 ( .C (clk), .D (signal_15787), .Q (signal_15788) ) ;
    buf_clk cell_10908 ( .C (clk), .D (signal_15795), .Q (signal_15796) ) ;
    buf_clk cell_10916 ( .C (clk), .D (signal_15803), .Q (signal_15804) ) ;
    buf_clk cell_10924 ( .C (clk), .D (signal_15811), .Q (signal_15812) ) ;
    buf_clk cell_10932 ( .C (clk), .D (signal_15819), .Q (signal_15820) ) ;
    buf_clk cell_10940 ( .C (clk), .D (signal_15827), .Q (signal_15828) ) ;
    buf_clk cell_10948 ( .C (clk), .D (signal_15835), .Q (signal_15836) ) ;
    buf_clk cell_10956 ( .C (clk), .D (signal_15843), .Q (signal_15844) ) ;
    buf_clk cell_10964 ( .C (clk), .D (signal_15851), .Q (signal_15852) ) ;
    buf_clk cell_10972 ( .C (clk), .D (signal_15859), .Q (signal_15860) ) ;
    buf_clk cell_10980 ( .C (clk), .D (signal_15867), .Q (signal_15868) ) ;
    buf_clk cell_10988 ( .C (clk), .D (signal_15875), .Q (signal_15876) ) ;
    buf_clk cell_10996 ( .C (clk), .D (signal_15883), .Q (signal_15884) ) ;
    buf_clk cell_11004 ( .C (clk), .D (signal_15891), .Q (signal_15892) ) ;
    buf_clk cell_11012 ( .C (clk), .D (signal_15899), .Q (signal_15900) ) ;
    buf_clk cell_11020 ( .C (clk), .D (signal_15907), .Q (signal_15908) ) ;
    buf_clk cell_11028 ( .C (clk), .D (signal_15915), .Q (signal_15916) ) ;
    buf_clk cell_11036 ( .C (clk), .D (signal_15923), .Q (signal_15924) ) ;
    buf_clk cell_11044 ( .C (clk), .D (signal_15931), .Q (signal_15932) ) ;
    buf_clk cell_11052 ( .C (clk), .D (signal_15939), .Q (signal_15940) ) ;
    buf_clk cell_11060 ( .C (clk), .D (signal_15947), .Q (signal_15948) ) ;
    buf_clk cell_11068 ( .C (clk), .D (signal_15955), .Q (signal_15956) ) ;
    buf_clk cell_11076 ( .C (clk), .D (signal_15963), .Q (signal_15964) ) ;
    buf_clk cell_11084 ( .C (clk), .D (signal_15971), .Q (signal_15972) ) ;
    buf_clk cell_11092 ( .C (clk), .D (signal_15979), .Q (signal_15980) ) ;
    buf_clk cell_11100 ( .C (clk), .D (signal_15987), .Q (signal_15988) ) ;
    buf_clk cell_11108 ( .C (clk), .D (signal_15995), .Q (signal_15996) ) ;
    buf_clk cell_11116 ( .C (clk), .D (signal_16003), .Q (signal_16004) ) ;
    buf_clk cell_11124 ( .C (clk), .D (signal_16011), .Q (signal_16012) ) ;
    buf_clk cell_11132 ( .C (clk), .D (signal_16019), .Q (signal_16020) ) ;
    buf_clk cell_11140 ( .C (clk), .D (signal_16027), .Q (signal_16028) ) ;
    buf_clk cell_11148 ( .C (clk), .D (signal_16035), .Q (signal_16036) ) ;
    buf_clk cell_11156 ( .C (clk), .D (signal_16043), .Q (signal_16044) ) ;
    buf_clk cell_11164 ( .C (clk), .D (signal_16051), .Q (signal_16052) ) ;
    buf_clk cell_11172 ( .C (clk), .D (signal_16059), .Q (signal_16060) ) ;
    buf_clk cell_11180 ( .C (clk), .D (signal_16067), .Q (signal_16068) ) ;
    buf_clk cell_11188 ( .C (clk), .D (signal_16075), .Q (signal_16076) ) ;
    buf_clk cell_11196 ( .C (clk), .D (signal_16083), .Q (signal_16084) ) ;
    buf_clk cell_11204 ( .C (clk), .D (signal_16091), .Q (signal_16092) ) ;
    buf_clk cell_11212 ( .C (clk), .D (signal_16099), .Q (signal_16100) ) ;
    buf_clk cell_11220 ( .C (clk), .D (signal_16107), .Q (signal_16108) ) ;
    buf_clk cell_11228 ( .C (clk), .D (signal_16115), .Q (signal_16116) ) ;
    buf_clk cell_11236 ( .C (clk), .D (signal_16123), .Q (signal_16124) ) ;
    buf_clk cell_11244 ( .C (clk), .D (signal_16131), .Q (signal_16132) ) ;
    buf_clk cell_11252 ( .C (clk), .D (signal_16139), .Q (signal_16140) ) ;
    buf_clk cell_11260 ( .C (clk), .D (signal_16147), .Q (signal_16148) ) ;
    buf_clk cell_11268 ( .C (clk), .D (signal_16155), .Q (signal_16156) ) ;
    buf_clk cell_11276 ( .C (clk), .D (signal_16163), .Q (signal_16164) ) ;
    buf_clk cell_11284 ( .C (clk), .D (signal_16171), .Q (signal_16172) ) ;
    buf_clk cell_11292 ( .C (clk), .D (signal_16179), .Q (signal_16180) ) ;
    buf_clk cell_11300 ( .C (clk), .D (signal_16187), .Q (signal_16188) ) ;
    buf_clk cell_11308 ( .C (clk), .D (signal_16195), .Q (signal_16196) ) ;
    buf_clk cell_11316 ( .C (clk), .D (signal_16203), .Q (signal_16204) ) ;
    buf_clk cell_11324 ( .C (clk), .D (signal_16211), .Q (signal_16212) ) ;
    buf_clk cell_11332 ( .C (clk), .D (signal_16219), .Q (signal_16220) ) ;
    buf_clk cell_11340 ( .C (clk), .D (signal_16227), .Q (signal_16228) ) ;
    buf_clk cell_11348 ( .C (clk), .D (signal_16235), .Q (signal_16236) ) ;
    buf_clk cell_11356 ( .C (clk), .D (signal_16243), .Q (signal_16244) ) ;
    buf_clk cell_11364 ( .C (clk), .D (signal_16251), .Q (signal_16252) ) ;
    buf_clk cell_11372 ( .C (clk), .D (signal_16259), .Q (signal_16260) ) ;
    buf_clk cell_11380 ( .C (clk), .D (signal_16267), .Q (signal_16268) ) ;
    buf_clk cell_11388 ( .C (clk), .D (signal_16275), .Q (signal_16276) ) ;
    buf_clk cell_11396 ( .C (clk), .D (signal_16283), .Q (signal_16284) ) ;
    buf_clk cell_11404 ( .C (clk), .D (signal_16291), .Q (signal_16292) ) ;
    buf_clk cell_11412 ( .C (clk), .D (signal_16299), .Q (signal_16300) ) ;
    buf_clk cell_11420 ( .C (clk), .D (signal_16307), .Q (signal_16308) ) ;
    buf_clk cell_11428 ( .C (clk), .D (signal_16315), .Q (signal_16316) ) ;
    buf_clk cell_11436 ( .C (clk), .D (signal_16323), .Q (signal_16324) ) ;
    buf_clk cell_11444 ( .C (clk), .D (signal_16331), .Q (signal_16332) ) ;
    buf_clk cell_11452 ( .C (clk), .D (signal_16339), .Q (signal_16340) ) ;
    buf_clk cell_11460 ( .C (clk), .D (signal_16347), .Q (signal_16348) ) ;
    buf_clk cell_11468 ( .C (clk), .D (signal_16355), .Q (signal_16356) ) ;
    buf_clk cell_11476 ( .C (clk), .D (signal_16363), .Q (signal_16364) ) ;
    buf_clk cell_11484 ( .C (clk), .D (signal_16371), .Q (signal_16372) ) ;
    buf_clk cell_11492 ( .C (clk), .D (signal_16379), .Q (signal_16380) ) ;
    buf_clk cell_11500 ( .C (clk), .D (signal_16387), .Q (signal_16388) ) ;
    buf_clk cell_11508 ( .C (clk), .D (signal_16395), .Q (signal_16396) ) ;
    buf_clk cell_11516 ( .C (clk), .D (signal_16403), .Q (signal_16404) ) ;
    buf_clk cell_11524 ( .C (clk), .D (signal_16411), .Q (signal_16412) ) ;
    buf_clk cell_11532 ( .C (clk), .D (signal_16419), .Q (signal_16420) ) ;
    buf_clk cell_11540 ( .C (clk), .D (signal_16427), .Q (signal_16428) ) ;
    buf_clk cell_11548 ( .C (clk), .D (signal_16435), .Q (signal_16436) ) ;
    buf_clk cell_11556 ( .C (clk), .D (signal_16443), .Q (signal_16444) ) ;
    buf_clk cell_11564 ( .C (clk), .D (signal_16451), .Q (signal_16452) ) ;
    buf_clk cell_11572 ( .C (clk), .D (signal_16459), .Q (signal_16460) ) ;
    buf_clk cell_11580 ( .C (clk), .D (signal_16467), .Q (signal_16468) ) ;
    buf_clk cell_11588 ( .C (clk), .D (signal_16475), .Q (signal_16476) ) ;
    buf_clk cell_11596 ( .C (clk), .D (signal_16483), .Q (signal_16484) ) ;
    buf_clk cell_11604 ( .C (clk), .D (signal_16491), .Q (signal_16492) ) ;
    buf_clk cell_11612 ( .C (clk), .D (signal_16499), .Q (signal_16500) ) ;
    buf_clk cell_11620 ( .C (clk), .D (signal_16507), .Q (signal_16508) ) ;
    buf_clk cell_11628 ( .C (clk), .D (signal_16515), .Q (signal_16516) ) ;
    buf_clk cell_11636 ( .C (clk), .D (signal_16523), .Q (signal_16524) ) ;
    buf_clk cell_11644 ( .C (clk), .D (signal_16531), .Q (signal_16532) ) ;
    buf_clk cell_11652 ( .C (clk), .D (signal_16539), .Q (signal_16540) ) ;
    buf_clk cell_11660 ( .C (clk), .D (signal_16547), .Q (signal_16548) ) ;
    buf_clk cell_11668 ( .C (clk), .D (signal_16555), .Q (signal_16556) ) ;
    buf_clk cell_11676 ( .C (clk), .D (signal_16563), .Q (signal_16564) ) ;
    buf_clk cell_11684 ( .C (clk), .D (signal_16571), .Q (signal_16572) ) ;
    buf_clk cell_11692 ( .C (clk), .D (signal_16579), .Q (signal_16580) ) ;
    buf_clk cell_11700 ( .C (clk), .D (signal_16587), .Q (signal_16588) ) ;
    buf_clk cell_11708 ( .C (clk), .D (signal_16595), .Q (signal_16596) ) ;
    buf_clk cell_11716 ( .C (clk), .D (signal_16603), .Q (signal_16604) ) ;
    buf_clk cell_11724 ( .C (clk), .D (signal_16611), .Q (signal_16612) ) ;
    buf_clk cell_11732 ( .C (clk), .D (signal_16619), .Q (signal_16620) ) ;
    buf_clk cell_11740 ( .C (clk), .D (signal_16627), .Q (signal_16628) ) ;
    buf_clk cell_11748 ( .C (clk), .D (signal_16635), .Q (signal_16636) ) ;
    buf_clk cell_11756 ( .C (clk), .D (signal_16643), .Q (signal_16644) ) ;
    buf_clk cell_11764 ( .C (clk), .D (signal_16651), .Q (signal_16652) ) ;
    buf_clk cell_11772 ( .C (clk), .D (signal_16659), .Q (signal_16660) ) ;
    buf_clk cell_11780 ( .C (clk), .D (signal_16667), .Q (signal_16668) ) ;
    buf_clk cell_11788 ( .C (clk), .D (signal_16675), .Q (signal_16676) ) ;
    buf_clk cell_11796 ( .C (clk), .D (signal_16683), .Q (signal_16684) ) ;
    buf_clk cell_11804 ( .C (clk), .D (signal_16691), .Q (signal_16692) ) ;
    buf_clk cell_11812 ( .C (clk), .D (signal_16699), .Q (signal_16700) ) ;
    buf_clk cell_11820 ( .C (clk), .D (signal_16707), .Q (signal_16708) ) ;
    buf_clk cell_11828 ( .C (clk), .D (signal_16715), .Q (signal_16716) ) ;
    buf_clk cell_11836 ( .C (clk), .D (signal_16723), .Q (signal_16724) ) ;
    buf_clk cell_11844 ( .C (clk), .D (signal_16731), .Q (signal_16732) ) ;
    buf_clk cell_11852 ( .C (clk), .D (signal_16739), .Q (signal_16740) ) ;
    buf_clk cell_11860 ( .C (clk), .D (signal_16747), .Q (signal_16748) ) ;
    buf_clk cell_11868 ( .C (clk), .D (signal_16755), .Q (signal_16756) ) ;
    buf_clk cell_11876 ( .C (clk), .D (signal_16763), .Q (signal_16764) ) ;
    buf_clk cell_11884 ( .C (clk), .D (signal_16771), .Q (signal_16772) ) ;
    buf_clk cell_11892 ( .C (clk), .D (signal_16779), .Q (signal_16780) ) ;
    buf_clk cell_11900 ( .C (clk), .D (signal_16787), .Q (signal_16788) ) ;
    buf_clk cell_11908 ( .C (clk), .D (signal_16795), .Q (signal_16796) ) ;
    buf_clk cell_11916 ( .C (clk), .D (signal_16803), .Q (signal_16804) ) ;
    buf_clk cell_11924 ( .C (clk), .D (signal_16811), .Q (signal_16812) ) ;
    buf_clk cell_11932 ( .C (clk), .D (signal_16819), .Q (signal_16820) ) ;
    buf_clk cell_11940 ( .C (clk), .D (signal_16827), .Q (signal_16828) ) ;
    buf_clk cell_11948 ( .C (clk), .D (signal_16835), .Q (signal_16836) ) ;
    buf_clk cell_11956 ( .C (clk), .D (signal_16843), .Q (signal_16844) ) ;
    buf_clk cell_11964 ( .C (clk), .D (signal_16851), .Q (signal_16852) ) ;
    buf_clk cell_11972 ( .C (clk), .D (signal_16859), .Q (signal_16860) ) ;
    buf_clk cell_11980 ( .C (clk), .D (signal_16867), .Q (signal_16868) ) ;
    buf_clk cell_11988 ( .C (clk), .D (signal_16875), .Q (signal_16876) ) ;
    buf_clk cell_11996 ( .C (clk), .D (signal_16883), .Q (signal_16884) ) ;
    buf_clk cell_12004 ( .C (clk), .D (signal_16891), .Q (signal_16892) ) ;
    buf_clk cell_12012 ( .C (clk), .D (signal_16899), .Q (signal_16900) ) ;
    buf_clk cell_12020 ( .C (clk), .D (signal_16907), .Q (signal_16908) ) ;
    buf_clk cell_12028 ( .C (clk), .D (signal_16915), .Q (signal_16916) ) ;
    buf_clk cell_12036 ( .C (clk), .D (signal_16923), .Q (signal_16924) ) ;
    buf_clk cell_12044 ( .C (clk), .D (signal_16931), .Q (signal_16932) ) ;
    buf_clk cell_12052 ( .C (clk), .D (signal_16939), .Q (signal_16940) ) ;
    buf_clk cell_12060 ( .C (clk), .D (signal_16947), .Q (signal_16948) ) ;
    buf_clk cell_12068 ( .C (clk), .D (signal_16955), .Q (signal_16956) ) ;
    buf_clk cell_12076 ( .C (clk), .D (signal_16963), .Q (signal_16964) ) ;
    buf_clk cell_12084 ( .C (clk), .D (signal_16971), .Q (signal_16972) ) ;
    buf_clk cell_12092 ( .C (clk), .D (signal_16979), .Q (signal_16980) ) ;
    buf_clk cell_12100 ( .C (clk), .D (signal_16987), .Q (signal_16988) ) ;
    buf_clk cell_12108 ( .C (clk), .D (signal_16995), .Q (signal_16996) ) ;
    buf_clk cell_12116 ( .C (clk), .D (signal_17003), .Q (signal_17004) ) ;
    buf_clk cell_12124 ( .C (clk), .D (signal_17011), .Q (signal_17012) ) ;
    buf_clk cell_12132 ( .C (clk), .D (signal_17019), .Q (signal_17020) ) ;
    buf_clk cell_12140 ( .C (clk), .D (signal_17027), .Q (signal_17028) ) ;
    buf_clk cell_12148 ( .C (clk), .D (signal_17035), .Q (signal_17036) ) ;
    buf_clk cell_12156 ( .C (clk), .D (signal_17043), .Q (signal_17044) ) ;
    buf_clk cell_12164 ( .C (clk), .D (signal_17051), .Q (signal_17052) ) ;
    buf_clk cell_12172 ( .C (clk), .D (signal_17059), .Q (signal_17060) ) ;
    buf_clk cell_12180 ( .C (clk), .D (signal_17067), .Q (signal_17068) ) ;
    buf_clk cell_12188 ( .C (clk), .D (signal_17075), .Q (signal_17076) ) ;
    buf_clk cell_12196 ( .C (clk), .D (signal_17083), .Q (signal_17084) ) ;
    buf_clk cell_12204 ( .C (clk), .D (signal_17091), .Q (signal_17092) ) ;
    buf_clk cell_12212 ( .C (clk), .D (signal_17099), .Q (signal_17100) ) ;
    buf_clk cell_12220 ( .C (clk), .D (signal_17107), .Q (signal_17108) ) ;
    buf_clk cell_12228 ( .C (clk), .D (signal_17115), .Q (signal_17116) ) ;
    buf_clk cell_12236 ( .C (clk), .D (signal_17123), .Q (signal_17124) ) ;
    buf_clk cell_12244 ( .C (clk), .D (signal_17131), .Q (signal_17132) ) ;
    buf_clk cell_12252 ( .C (clk), .D (signal_17139), .Q (signal_17140) ) ;
    buf_clk cell_12260 ( .C (clk), .D (signal_17147), .Q (signal_17148) ) ;
    buf_clk cell_12268 ( .C (clk), .D (signal_17155), .Q (signal_17156) ) ;
    buf_clk cell_12276 ( .C (clk), .D (signal_17163), .Q (signal_17164) ) ;
    buf_clk cell_12284 ( .C (clk), .D (signal_17171), .Q (signal_17172) ) ;
    buf_clk cell_12292 ( .C (clk), .D (signal_17179), .Q (signal_17180) ) ;
    buf_clk cell_12300 ( .C (clk), .D (signal_17187), .Q (signal_17188) ) ;
    buf_clk cell_12308 ( .C (clk), .D (signal_17195), .Q (signal_17196) ) ;
    buf_clk cell_12316 ( .C (clk), .D (signal_17203), .Q (signal_17204) ) ;
    buf_clk cell_12324 ( .C (clk), .D (signal_17211), .Q (signal_17212) ) ;
    buf_clk cell_12332 ( .C (clk), .D (signal_17219), .Q (signal_17220) ) ;
    buf_clk cell_12340 ( .C (clk), .D (signal_17227), .Q (signal_17228) ) ;
    buf_clk cell_12348 ( .C (clk), .D (signal_17235), .Q (signal_17236) ) ;
    buf_clk cell_12356 ( .C (clk), .D (signal_17243), .Q (signal_17244) ) ;
    buf_clk cell_12364 ( .C (clk), .D (signal_17251), .Q (signal_17252) ) ;
    buf_clk cell_12372 ( .C (clk), .D (signal_17259), .Q (signal_17260) ) ;
    buf_clk cell_12380 ( .C (clk), .D (signal_17267), .Q (signal_17268) ) ;
    buf_clk cell_12388 ( .C (clk), .D (signal_17275), .Q (signal_17276) ) ;
    buf_clk cell_12396 ( .C (clk), .D (signal_17283), .Q (signal_17284) ) ;
    buf_clk cell_12404 ( .C (clk), .D (signal_17291), .Q (signal_17292) ) ;
    buf_clk cell_12412 ( .C (clk), .D (signal_17299), .Q (signal_17300) ) ;
    buf_clk cell_12420 ( .C (clk), .D (signal_17307), .Q (signal_17308) ) ;
    buf_clk cell_12428 ( .C (clk), .D (signal_17315), .Q (signal_17316) ) ;
    buf_clk cell_12436 ( .C (clk), .D (signal_17323), .Q (signal_17324) ) ;
    buf_clk cell_12444 ( .C (clk), .D (signal_17331), .Q (signal_17332) ) ;
    buf_clk cell_12452 ( .C (clk), .D (signal_17339), .Q (signal_17340) ) ;
    buf_clk cell_12460 ( .C (clk), .D (signal_17347), .Q (signal_17348) ) ;
    buf_clk cell_12468 ( .C (clk), .D (signal_17355), .Q (signal_17356) ) ;
    buf_clk cell_12476 ( .C (clk), .D (signal_17363), .Q (signal_17364) ) ;
    buf_clk cell_12484 ( .C (clk), .D (signal_17371), .Q (signal_17372) ) ;
    buf_clk cell_12492 ( .C (clk), .D (signal_17379), .Q (signal_17380) ) ;
    buf_clk cell_12500 ( .C (clk), .D (signal_17387), .Q (signal_17388) ) ;
    buf_clk cell_12508 ( .C (clk), .D (signal_17395), .Q (signal_17396) ) ;
    buf_clk cell_12516 ( .C (clk), .D (signal_17403), .Q (signal_17404) ) ;
    buf_clk cell_12524 ( .C (clk), .D (signal_17411), .Q (signal_17412) ) ;
    buf_clk cell_12532 ( .C (clk), .D (signal_17419), .Q (signal_17420) ) ;
    buf_clk cell_12540 ( .C (clk), .D (signal_17427), .Q (signal_17428) ) ;
    buf_clk cell_12548 ( .C (clk), .D (signal_17435), .Q (signal_17436) ) ;
    buf_clk cell_12556 ( .C (clk), .D (signal_17443), .Q (signal_17444) ) ;
    buf_clk cell_12564 ( .C (clk), .D (signal_17451), .Q (signal_17452) ) ;
    buf_clk cell_12572 ( .C (clk), .D (signal_17459), .Q (signal_17460) ) ;
    buf_clk cell_12580 ( .C (clk), .D (signal_17467), .Q (signal_17468) ) ;
    buf_clk cell_12588 ( .C (clk), .D (signal_17475), .Q (signal_17476) ) ;
    buf_clk cell_12596 ( .C (clk), .D (signal_17483), .Q (signal_17484) ) ;
    buf_clk cell_12604 ( .C (clk), .D (signal_17491), .Q (signal_17492) ) ;
    buf_clk cell_12612 ( .C (clk), .D (signal_17499), .Q (signal_17500) ) ;
    buf_clk cell_12620 ( .C (clk), .D (signal_17507), .Q (signal_17508) ) ;
    buf_clk cell_12628 ( .C (clk), .D (signal_17515), .Q (signal_17516) ) ;
    buf_clk cell_12636 ( .C (clk), .D (signal_17523), .Q (signal_17524) ) ;
    buf_clk cell_12644 ( .C (clk), .D (signal_17531), .Q (signal_17532) ) ;
    buf_clk cell_12652 ( .C (clk), .D (signal_17539), .Q (signal_17540) ) ;
    buf_clk cell_12660 ( .C (clk), .D (signal_17547), .Q (signal_17548) ) ;
    buf_clk cell_12668 ( .C (clk), .D (signal_17555), .Q (signal_17556) ) ;
    buf_clk cell_12676 ( .C (clk), .D (signal_17563), .Q (signal_17564) ) ;
    buf_clk cell_12684 ( .C (clk), .D (signal_17571), .Q (signal_17572) ) ;
    buf_clk cell_12692 ( .C (clk), .D (signal_17579), .Q (signal_17580) ) ;
    buf_clk cell_12700 ( .C (clk), .D (signal_17587), .Q (signal_17588) ) ;
    buf_clk cell_12708 ( .C (clk), .D (signal_17595), .Q (signal_17596) ) ;
    buf_clk cell_12716 ( .C (clk), .D (signal_17603), .Q (signal_17604) ) ;
    buf_clk cell_12724 ( .C (clk), .D (signal_17611), .Q (signal_17612) ) ;
    buf_clk cell_12732 ( .C (clk), .D (signal_17619), .Q (signal_17620) ) ;
    buf_clk cell_12740 ( .C (clk), .D (signal_17627), .Q (signal_17628) ) ;
    buf_clk cell_12748 ( .C (clk), .D (signal_17635), .Q (signal_17636) ) ;
    buf_clk cell_12756 ( .C (clk), .D (signal_17643), .Q (signal_17644) ) ;
    buf_clk cell_12764 ( .C (clk), .D (signal_17651), .Q (signal_17652) ) ;
    buf_clk cell_12772 ( .C (clk), .D (signal_17659), .Q (signal_17660) ) ;
    buf_clk cell_12780 ( .C (clk), .D (signal_17667), .Q (signal_17668) ) ;
    buf_clk cell_12788 ( .C (clk), .D (signal_17675), .Q (signal_17676) ) ;
    buf_clk cell_12796 ( .C (clk), .D (signal_17683), .Q (signal_17684) ) ;
    buf_clk cell_12804 ( .C (clk), .D (signal_17691), .Q (signal_17692) ) ;
    buf_clk cell_12812 ( .C (clk), .D (signal_17699), .Q (signal_17700) ) ;
    buf_clk cell_12820 ( .C (clk), .D (signal_17707), .Q (signal_17708) ) ;
    buf_clk cell_12828 ( .C (clk), .D (signal_17715), .Q (signal_17716) ) ;
    buf_clk cell_12836 ( .C (clk), .D (signal_17723), .Q (signal_17724) ) ;
    buf_clk cell_12844 ( .C (clk), .D (signal_17731), .Q (signal_17732) ) ;
    buf_clk cell_12852 ( .C (clk), .D (signal_17739), .Q (signal_17740) ) ;
    buf_clk cell_12860 ( .C (clk), .D (signal_17747), .Q (signal_17748) ) ;
    buf_clk cell_12868 ( .C (clk), .D (signal_17755), .Q (signal_17756) ) ;
    buf_clk cell_12876 ( .C (clk), .D (signal_17763), .Q (signal_17764) ) ;
    buf_clk cell_12884 ( .C (clk), .D (signal_17771), .Q (signal_17772) ) ;
    buf_clk cell_12892 ( .C (clk), .D (signal_17779), .Q (signal_17780) ) ;
    buf_clk cell_12900 ( .C (clk), .D (signal_17787), .Q (signal_17788) ) ;
    buf_clk cell_12908 ( .C (clk), .D (signal_17795), .Q (signal_17796) ) ;
    buf_clk cell_12916 ( .C (clk), .D (signal_17803), .Q (signal_17804) ) ;
    buf_clk cell_12924 ( .C (clk), .D (signal_17811), .Q (signal_17812) ) ;
    buf_clk cell_12932 ( .C (clk), .D (signal_17819), .Q (signal_17820) ) ;
    buf_clk cell_12940 ( .C (clk), .D (signal_17827), .Q (signal_17828) ) ;
    buf_clk cell_12948 ( .C (clk), .D (signal_17835), .Q (signal_17836) ) ;
    buf_clk cell_12956 ( .C (clk), .D (signal_17843), .Q (signal_17844) ) ;
    buf_clk cell_12964 ( .C (clk), .D (signal_17851), .Q (signal_17852) ) ;
    buf_clk cell_12972 ( .C (clk), .D (signal_17859), .Q (signal_17860) ) ;
    buf_clk cell_12980 ( .C (clk), .D (signal_17867), .Q (signal_17868) ) ;
    buf_clk cell_12988 ( .C (clk), .D (signal_17875), .Q (signal_17876) ) ;
    buf_clk cell_12996 ( .C (clk), .D (signal_17883), .Q (signal_17884) ) ;
    buf_clk cell_13004 ( .C (clk), .D (signal_17891), .Q (signal_17892) ) ;
    buf_clk cell_13012 ( .C (clk), .D (signal_17899), .Q (signal_17900) ) ;
    buf_clk cell_13020 ( .C (clk), .D (signal_17907), .Q (signal_17908) ) ;
    buf_clk cell_13028 ( .C (clk), .D (signal_17915), .Q (signal_17916) ) ;
    buf_clk cell_13036 ( .C (clk), .D (signal_17923), .Q (signal_17924) ) ;
    buf_clk cell_13044 ( .C (clk), .D (signal_17931), .Q (signal_17932) ) ;
    buf_clk cell_13052 ( .C (clk), .D (signal_17939), .Q (signal_17940) ) ;
    buf_clk cell_13060 ( .C (clk), .D (signal_17947), .Q (signal_17948) ) ;
    buf_clk cell_13068 ( .C (clk), .D (signal_17955), .Q (signal_17956) ) ;
    buf_clk cell_13076 ( .C (clk), .D (signal_17963), .Q (signal_17964) ) ;
    buf_clk cell_13084 ( .C (clk), .D (signal_17971), .Q (signal_17972) ) ;
    buf_clk cell_13092 ( .C (clk), .D (signal_17979), .Q (signal_17980) ) ;
    buf_clk cell_13100 ( .C (clk), .D (signal_17987), .Q (signal_17988) ) ;
    buf_clk cell_13108 ( .C (clk), .D (signal_17995), .Q (signal_17996) ) ;
    buf_clk cell_13116 ( .C (clk), .D (signal_18003), .Q (signal_18004) ) ;
    buf_clk cell_13124 ( .C (clk), .D (signal_18011), .Q (signal_18012) ) ;
    buf_clk cell_13132 ( .C (clk), .D (signal_18019), .Q (signal_18020) ) ;
    buf_clk cell_13140 ( .C (clk), .D (signal_18027), .Q (signal_18028) ) ;
    buf_clk cell_13148 ( .C (clk), .D (signal_18035), .Q (signal_18036) ) ;
    buf_clk cell_13156 ( .C (clk), .D (signal_18043), .Q (signal_18044) ) ;
    buf_clk cell_13164 ( .C (clk), .D (signal_18051), .Q (signal_18052) ) ;
    buf_clk cell_13172 ( .C (clk), .D (signal_18059), .Q (signal_18060) ) ;
    buf_clk cell_13180 ( .C (clk), .D (signal_18067), .Q (signal_18068) ) ;
    buf_clk cell_13188 ( .C (clk), .D (signal_18075), .Q (signal_18076) ) ;
    buf_clk cell_13196 ( .C (clk), .D (signal_18083), .Q (signal_18084) ) ;
    buf_clk cell_13204 ( .C (clk), .D (signal_18091), .Q (signal_18092) ) ;
    buf_clk cell_13212 ( .C (clk), .D (signal_18099), .Q (signal_18100) ) ;
    buf_clk cell_13220 ( .C (clk), .D (signal_18107), .Q (signal_18108) ) ;
    buf_clk cell_13228 ( .C (clk), .D (signal_18115), .Q (signal_18116) ) ;
    buf_clk cell_13236 ( .C (clk), .D (signal_18123), .Q (signal_18124) ) ;
    buf_clk cell_13244 ( .C (clk), .D (signal_18131), .Q (signal_18132) ) ;
    buf_clk cell_13252 ( .C (clk), .D (signal_18139), .Q (signal_18140) ) ;
    buf_clk cell_13260 ( .C (clk), .D (signal_18147), .Q (signal_18148) ) ;
    buf_clk cell_13268 ( .C (clk), .D (signal_18155), .Q (signal_18156) ) ;
    buf_clk cell_13276 ( .C (clk), .D (signal_18163), .Q (signal_18164) ) ;
    buf_clk cell_17592 ( .C (clk), .D (signal_22479), .Q (signal_22480) ) ;
    buf_clk cell_17600 ( .C (clk), .D (signal_22487), .Q (signal_22488) ) ;
    buf_clk cell_17608 ( .C (clk), .D (signal_22495), .Q (signal_22496) ) ;
    buf_clk cell_17616 ( .C (clk), .D (signal_22503), .Q (signal_22504) ) ;
    buf_clk cell_17624 ( .C (clk), .D (signal_22511), .Q (signal_22512) ) ;
    buf_clk cell_17632 ( .C (clk), .D (signal_22519), .Q (signal_22520) ) ;
    buf_clk cell_17640 ( .C (clk), .D (signal_22527), .Q (signal_22528) ) ;
    buf_clk cell_17648 ( .C (clk), .D (signal_22535), .Q (signal_22536) ) ;
    buf_clk cell_17656 ( .C (clk), .D (signal_22543), .Q (signal_22544) ) ;
    buf_clk cell_17664 ( .C (clk), .D (signal_22551), .Q (signal_22552) ) ;
    buf_clk cell_17672 ( .C (clk), .D (signal_22559), .Q (signal_22560) ) ;
    buf_clk cell_17680 ( .C (clk), .D (signal_22567), .Q (signal_22568) ) ;
    buf_clk cell_17688 ( .C (clk), .D (signal_22575), .Q (signal_22576) ) ;
    buf_clk cell_17696 ( .C (clk), .D (signal_22583), .Q (signal_22584) ) ;
    buf_clk cell_17704 ( .C (clk), .D (signal_22591), .Q (signal_22592) ) ;
    buf_clk cell_17712 ( .C (clk), .D (signal_22599), .Q (signal_22600) ) ;
    buf_clk cell_17720 ( .C (clk), .D (signal_22607), .Q (signal_22608) ) ;
    buf_clk cell_17728 ( .C (clk), .D (signal_22615), .Q (signal_22616) ) ;
    buf_clk cell_17736 ( .C (clk), .D (signal_22623), .Q (signal_22624) ) ;
    buf_clk cell_17744 ( .C (clk), .D (signal_22631), .Q (signal_22632) ) ;
    buf_clk cell_17752 ( .C (clk), .D (signal_22639), .Q (signal_22640) ) ;
    buf_clk cell_17760 ( .C (clk), .D (signal_22647), .Q (signal_22648) ) ;
    buf_clk cell_17768 ( .C (clk), .D (signal_22655), .Q (signal_22656) ) ;
    buf_clk cell_17776 ( .C (clk), .D (signal_22663), .Q (signal_22664) ) ;
    buf_clk cell_17784 ( .C (clk), .D (signal_22671), .Q (signal_22672) ) ;
    buf_clk cell_17792 ( .C (clk), .D (signal_22679), .Q (signal_22680) ) ;
    buf_clk cell_17800 ( .C (clk), .D (signal_22687), .Q (signal_22688) ) ;
    buf_clk cell_17808 ( .C (clk), .D (signal_22695), .Q (signal_22696) ) ;
    buf_clk cell_17816 ( .C (clk), .D (signal_22703), .Q (signal_22704) ) ;
    buf_clk cell_17824 ( .C (clk), .D (signal_22711), .Q (signal_22712) ) ;
    buf_clk cell_17832 ( .C (clk), .D (signal_22719), .Q (signal_22720) ) ;
    buf_clk cell_17840 ( .C (clk), .D (signal_22727), .Q (signal_22728) ) ;
    buf_clk cell_17848 ( .C (clk), .D (signal_22735), .Q (signal_22736) ) ;
    buf_clk cell_17856 ( .C (clk), .D (signal_22743), .Q (signal_22744) ) ;
    buf_clk cell_17864 ( .C (clk), .D (signal_22751), .Q (signal_22752) ) ;
    buf_clk cell_17872 ( .C (clk), .D (signal_22759), .Q (signal_22760) ) ;
    buf_clk cell_17880 ( .C (clk), .D (signal_22767), .Q (signal_22768) ) ;
    buf_clk cell_17888 ( .C (clk), .D (signal_22775), .Q (signal_22776) ) ;
    buf_clk cell_17896 ( .C (clk), .D (signal_22783), .Q (signal_22784) ) ;
    buf_clk cell_17904 ( .C (clk), .D (signal_22791), .Q (signal_22792) ) ;
    buf_clk cell_17912 ( .C (clk), .D (signal_22799), .Q (signal_22800) ) ;
    buf_clk cell_17920 ( .C (clk), .D (signal_22807), .Q (signal_22808) ) ;
    buf_clk cell_17928 ( .C (clk), .D (signal_22815), .Q (signal_22816) ) ;
    buf_clk cell_17936 ( .C (clk), .D (signal_22823), .Q (signal_22824) ) ;
    buf_clk cell_17944 ( .C (clk), .D (signal_22831), .Q (signal_22832) ) ;
    buf_clk cell_17952 ( .C (clk), .D (signal_22839), .Q (signal_22840) ) ;
    buf_clk cell_17960 ( .C (clk), .D (signal_22847), .Q (signal_22848) ) ;
    buf_clk cell_17968 ( .C (clk), .D (signal_22855), .Q (signal_22856) ) ;
    buf_clk cell_17976 ( .C (clk), .D (signal_22863), .Q (signal_22864) ) ;
    buf_clk cell_17984 ( .C (clk), .D (signal_22871), .Q (signal_22872) ) ;
    buf_clk cell_17992 ( .C (clk), .D (signal_22879), .Q (signal_22880) ) ;
    buf_clk cell_18000 ( .C (clk), .D (signal_22887), .Q (signal_22888) ) ;
    buf_clk cell_18008 ( .C (clk), .D (signal_22895), .Q (signal_22896) ) ;
    buf_clk cell_18016 ( .C (clk), .D (signal_22903), .Q (signal_22904) ) ;
    buf_clk cell_18024 ( .C (clk), .D (signal_22911), .Q (signal_22912) ) ;
    buf_clk cell_18032 ( .C (clk), .D (signal_22919), .Q (signal_22920) ) ;
    buf_clk cell_18040 ( .C (clk), .D (signal_22927), .Q (signal_22928) ) ;
    buf_clk cell_18048 ( .C (clk), .D (signal_22935), .Q (signal_22936) ) ;
    buf_clk cell_18056 ( .C (clk), .D (signal_22943), .Q (signal_22944) ) ;
    buf_clk cell_18064 ( .C (clk), .D (signal_22951), .Q (signal_22952) ) ;
    buf_clk cell_18072 ( .C (clk), .D (signal_22959), .Q (signal_22960) ) ;
    buf_clk cell_18080 ( .C (clk), .D (signal_22967), .Q (signal_22968) ) ;
    buf_clk cell_18088 ( .C (clk), .D (signal_22975), .Q (signal_22976) ) ;
    buf_clk cell_18096 ( .C (clk), .D (signal_22983), .Q (signal_22984) ) ;
    buf_clk cell_18104 ( .C (clk), .D (signal_22991), .Q (signal_22992) ) ;
    buf_clk cell_18112 ( .C (clk), .D (signal_22999), .Q (signal_23000) ) ;
    buf_clk cell_18120 ( .C (clk), .D (signal_23007), .Q (signal_23008) ) ;
    buf_clk cell_18128 ( .C (clk), .D (signal_23015), .Q (signal_23016) ) ;
    buf_clk cell_18136 ( .C (clk), .D (signal_23023), .Q (signal_23024) ) ;
    buf_clk cell_18144 ( .C (clk), .D (signal_23031), .Q (signal_23032) ) ;
    buf_clk cell_18152 ( .C (clk), .D (signal_23039), .Q (signal_23040) ) ;
    buf_clk cell_18160 ( .C (clk), .D (signal_23047), .Q (signal_23048) ) ;
    buf_clk cell_18168 ( .C (clk), .D (signal_23055), .Q (signal_23056) ) ;
    buf_clk cell_18176 ( .C (clk), .D (signal_23063), .Q (signal_23064) ) ;
    buf_clk cell_18184 ( .C (clk), .D (signal_23071), .Q (signal_23072) ) ;
    buf_clk cell_18192 ( .C (clk), .D (signal_23079), .Q (signal_23080) ) ;
    buf_clk cell_18200 ( .C (clk), .D (signal_23087), .Q (signal_23088) ) ;
    buf_clk cell_18208 ( .C (clk), .D (signal_23095), .Q (signal_23096) ) ;
    buf_clk cell_18216 ( .C (clk), .D (signal_23103), .Q (signal_23104) ) ;
    buf_clk cell_18224 ( .C (clk), .D (signal_23111), .Q (signal_23112) ) ;
    buf_clk cell_18232 ( .C (clk), .D (signal_23119), .Q (signal_23120) ) ;
    buf_clk cell_18240 ( .C (clk), .D (signal_23127), .Q (signal_23128) ) ;
    buf_clk cell_18248 ( .C (clk), .D (signal_23135), .Q (signal_23136) ) ;
    buf_clk cell_18256 ( .C (clk), .D (signal_23143), .Q (signal_23144) ) ;
    buf_clk cell_18264 ( .C (clk), .D (signal_23151), .Q (signal_23152) ) ;
    buf_clk cell_18272 ( .C (clk), .D (signal_23159), .Q (signal_23160) ) ;
    buf_clk cell_18280 ( .C (clk), .D (signal_23167), .Q (signal_23168) ) ;
    buf_clk cell_18288 ( .C (clk), .D (signal_23175), .Q (signal_23176) ) ;
    buf_clk cell_18296 ( .C (clk), .D (signal_23183), .Q (signal_23184) ) ;
    buf_clk cell_18304 ( .C (clk), .D (signal_23191), .Q (signal_23192) ) ;
    buf_clk cell_18312 ( .C (clk), .D (signal_23199), .Q (signal_23200) ) ;
    buf_clk cell_18320 ( .C (clk), .D (signal_23207), .Q (signal_23208) ) ;
    buf_clk cell_18328 ( .C (clk), .D (signal_23215), .Q (signal_23216) ) ;
    buf_clk cell_18336 ( .C (clk), .D (signal_23223), .Q (signal_23224) ) ;
    buf_clk cell_18344 ( .C (clk), .D (signal_23231), .Q (signal_23232) ) ;
    buf_clk cell_18352 ( .C (clk), .D (signal_23239), .Q (signal_23240) ) ;
    buf_clk cell_18360 ( .C (clk), .D (signal_23247), .Q (signal_23248) ) ;
    buf_clk cell_18368 ( .C (clk), .D (signal_23255), .Q (signal_23256) ) ;
    buf_clk cell_18376 ( .C (clk), .D (signal_23263), .Q (signal_23264) ) ;
    buf_clk cell_18384 ( .C (clk), .D (signal_23271), .Q (signal_23272) ) ;
    buf_clk cell_18392 ( .C (clk), .D (signal_23279), .Q (signal_23280) ) ;
    buf_clk cell_18400 ( .C (clk), .D (signal_23287), .Q (signal_23288) ) ;
    buf_clk cell_18402 ( .C (clk), .D (signal_23289), .Q (signal_23290) ) ;
    buf_clk cell_18404 ( .C (clk), .D (signal_23291), .Q (signal_23292) ) ;
    buf_clk cell_18412 ( .C (clk), .D (signal_23299), .Q (signal_23300) ) ;
    buf_clk cell_18420 ( .C (clk), .D (signal_23307), .Q (signal_23308) ) ;
    buf_clk cell_18428 ( .C (clk), .D (signal_23315), .Q (signal_23316) ) ;
    buf_clk cell_18436 ( .C (clk), .D (signal_23323), .Q (signal_23324) ) ;
    buf_clk cell_18444 ( .C (clk), .D (signal_23331), .Q (signal_23332) ) ;
    buf_clk cell_18452 ( .C (clk), .D (signal_23339), .Q (signal_23340) ) ;
    buf_clk cell_18460 ( .C (clk), .D (signal_23347), .Q (signal_23348) ) ;
    buf_clk cell_18468 ( .C (clk), .D (signal_23355), .Q (signal_23356) ) ;
    buf_clk cell_18476 ( .C (clk), .D (signal_23363), .Q (signal_23364) ) ;
    buf_clk cell_18484 ( .C (clk), .D (signal_23371), .Q (signal_23372) ) ;
    buf_clk cell_18492 ( .C (clk), .D (signal_23379), .Q (signal_23380) ) ;
    buf_clk cell_18500 ( .C (clk), .D (signal_23387), .Q (signal_23388) ) ;
    buf_clk cell_18508 ( .C (clk), .D (signal_23395), .Q (signal_23396) ) ;
    buf_clk cell_18516 ( .C (clk), .D (signal_23403), .Q (signal_23404) ) ;
    buf_clk cell_18524 ( .C (clk), .D (signal_23411), .Q (signal_23412) ) ;
    buf_clk cell_18532 ( .C (clk), .D (signal_23419), .Q (signal_23420) ) ;
    buf_clk cell_18540 ( .C (clk), .D (signal_23427), .Q (signal_23428) ) ;
    buf_clk cell_18548 ( .C (clk), .D (signal_23435), .Q (signal_23436) ) ;
    buf_clk cell_18556 ( .C (clk), .D (signal_23443), .Q (signal_23444) ) ;
    buf_clk cell_18564 ( .C (clk), .D (signal_23451), .Q (signal_23452) ) ;
    buf_clk cell_18572 ( .C (clk), .D (signal_23459), .Q (signal_23460) ) ;
    buf_clk cell_18580 ( .C (clk), .D (signal_23467), .Q (signal_23468) ) ;
    buf_clk cell_18588 ( .C (clk), .D (signal_23475), .Q (signal_23476) ) ;
    buf_clk cell_18596 ( .C (clk), .D (signal_23483), .Q (signal_23484) ) ;
    buf_clk cell_18604 ( .C (clk), .D (signal_23491), .Q (signal_23492) ) ;
    buf_clk cell_18612 ( .C (clk), .D (signal_23499), .Q (signal_23500) ) ;
    buf_clk cell_18620 ( .C (clk), .D (signal_23507), .Q (signal_23508) ) ;
    buf_clk cell_18628 ( .C (clk), .D (signal_23515), .Q (signal_23516) ) ;
    buf_clk cell_18636 ( .C (clk), .D (signal_23523), .Q (signal_23524) ) ;
    buf_clk cell_18644 ( .C (clk), .D (signal_23531), .Q (signal_23532) ) ;
    buf_clk cell_18646 ( .C (clk), .D (signal_23533), .Q (signal_23534) ) ;
    buf_clk cell_18648 ( .C (clk), .D (signal_23535), .Q (signal_23536) ) ;
    buf_clk cell_18656 ( .C (clk), .D (signal_23543), .Q (signal_23544) ) ;
    buf_clk cell_18664 ( .C (clk), .D (signal_23551), .Q (signal_23552) ) ;
    buf_clk cell_18672 ( .C (clk), .D (signal_23559), .Q (signal_23560) ) ;
    buf_clk cell_18680 ( .C (clk), .D (signal_23567), .Q (signal_23568) ) ;
    buf_clk cell_18688 ( .C (clk), .D (signal_23575), .Q (signal_23576) ) ;
    buf_clk cell_18696 ( .C (clk), .D (signal_23583), .Q (signal_23584) ) ;
    buf_clk cell_18704 ( .C (clk), .D (signal_23591), .Q (signal_23592) ) ;
    buf_clk cell_18712 ( .C (clk), .D (signal_23599), .Q (signal_23600) ) ;
    buf_clk cell_18720 ( .C (clk), .D (signal_23607), .Q (signal_23608) ) ;
    buf_clk cell_18728 ( .C (clk), .D (signal_23615), .Q (signal_23616) ) ;
    buf_clk cell_18736 ( .C (clk), .D (signal_23623), .Q (signal_23624) ) ;
    buf_clk cell_18744 ( .C (clk), .D (signal_23631), .Q (signal_23632) ) ;
    buf_clk cell_18746 ( .C (clk), .D (signal_23633), .Q (signal_23634) ) ;
    buf_clk cell_18748 ( .C (clk), .D (signal_23635), .Q (signal_23636) ) ;
    buf_clk cell_18756 ( .C (clk), .D (signal_23643), .Q (signal_23644) ) ;
    buf_clk cell_18764 ( .C (clk), .D (signal_23651), .Q (signal_23652) ) ;
    buf_clk cell_18772 ( .C (clk), .D (signal_23659), .Q (signal_23660) ) ;
    buf_clk cell_18780 ( .C (clk), .D (signal_23667), .Q (signal_23668) ) ;
    buf_clk cell_18788 ( .C (clk), .D (signal_23675), .Q (signal_23676) ) ;
    buf_clk cell_18796 ( .C (clk), .D (signal_23683), .Q (signal_23684) ) ;
    buf_clk cell_18804 ( .C (clk), .D (signal_23691), .Q (signal_23692) ) ;
    buf_clk cell_18812 ( .C (clk), .D (signal_23699), .Q (signal_23700) ) ;
    buf_clk cell_18820 ( .C (clk), .D (signal_23707), .Q (signal_23708) ) ;
    buf_clk cell_18828 ( .C (clk), .D (signal_23715), .Q (signal_23716) ) ;
    buf_clk cell_18836 ( .C (clk), .D (signal_23723), .Q (signal_23724) ) ;
    buf_clk cell_18844 ( .C (clk), .D (signal_23731), .Q (signal_23732) ) ;
    buf_clk cell_18852 ( .C (clk), .D (signal_23739), .Q (signal_23740) ) ;
    buf_clk cell_18860 ( .C (clk), .D (signal_23747), .Q (signal_23748) ) ;
    buf_clk cell_18868 ( .C (clk), .D (signal_23755), .Q (signal_23756) ) ;
    buf_clk cell_18876 ( .C (clk), .D (signal_23763), .Q (signal_23764) ) ;
    buf_clk cell_18884 ( .C (clk), .D (signal_23771), .Q (signal_23772) ) ;
    buf_clk cell_18892 ( .C (clk), .D (signal_23779), .Q (signal_23780) ) ;
    buf_clk cell_18900 ( .C (clk), .D (signal_23787), .Q (signal_23788) ) ;
    buf_clk cell_18908 ( .C (clk), .D (signal_23795), .Q (signal_23796) ) ;
    buf_clk cell_18916 ( .C (clk), .D (signal_23803), .Q (signal_23804) ) ;
    buf_clk cell_18924 ( .C (clk), .D (signal_23811), .Q (signal_23812) ) ;
    buf_clk cell_18932 ( .C (clk), .D (signal_23819), .Q (signal_23820) ) ;
    buf_clk cell_18940 ( .C (clk), .D (signal_23827), .Q (signal_23828) ) ;
    buf_clk cell_18948 ( .C (clk), .D (signal_23835), .Q (signal_23836) ) ;
    buf_clk cell_18956 ( .C (clk), .D (signal_23843), .Q (signal_23844) ) ;
    buf_clk cell_18964 ( .C (clk), .D (signal_23851), .Q (signal_23852) ) ;
    buf_clk cell_18972 ( .C (clk), .D (signal_23859), .Q (signal_23860) ) ;
    buf_clk cell_18980 ( .C (clk), .D (signal_23867), .Q (signal_23868) ) ;
    buf_clk cell_18988 ( .C (clk), .D (signal_23875), .Q (signal_23876) ) ;
    buf_clk cell_18996 ( .C (clk), .D (signal_23883), .Q (signal_23884) ) ;
    buf_clk cell_19004 ( .C (clk), .D (signal_23891), .Q (signal_23892) ) ;
    buf_clk cell_19012 ( .C (clk), .D (signal_23899), .Q (signal_23900) ) ;
    buf_clk cell_19020 ( .C (clk), .D (signal_23907), .Q (signal_23908) ) ;
    buf_clk cell_19028 ( .C (clk), .D (signal_23915), .Q (signal_23916) ) ;
    buf_clk cell_19036 ( .C (clk), .D (signal_23923), .Q (signal_23924) ) ;
    buf_clk cell_19044 ( .C (clk), .D (signal_23931), .Q (signal_23932) ) ;
    buf_clk cell_19052 ( .C (clk), .D (signal_23939), .Q (signal_23940) ) ;
    buf_clk cell_19060 ( .C (clk), .D (signal_23947), .Q (signal_23948) ) ;
    buf_clk cell_19068 ( .C (clk), .D (signal_23955), .Q (signal_23956) ) ;
    buf_clk cell_19076 ( .C (clk), .D (signal_23963), .Q (signal_23964) ) ;
    buf_clk cell_19084 ( .C (clk), .D (signal_23971), .Q (signal_23972) ) ;
    buf_clk cell_19092 ( .C (clk), .D (signal_23979), .Q (signal_23980) ) ;
    buf_clk cell_19100 ( .C (clk), .D (signal_23987), .Q (signal_23988) ) ;
    buf_clk cell_19108 ( .C (clk), .D (signal_23995), .Q (signal_23996) ) ;
    buf_clk cell_19116 ( .C (clk), .D (signal_24003), .Q (signal_24004) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_293 ( .clk (clk), .D ({signal_11592, signal_421}), .Q ({signal_7530, signal_3870}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_296 ( .clk (clk), .D ({signal_11758, signal_423}), .Q ({signal_7623, signal_3869}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_299 ( .clk (clk), .D ({signal_11459, signal_425}), .Q ({signal_7656, signal_3868}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_302 ( .clk (clk), .D ({signal_11594, signal_427}), .Q ({signal_7689, signal_3867}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_305 ( .clk (clk), .D ({signal_11596, signal_429}), .Q ({signal_7722, signal_3866}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_308 ( .clk (clk), .D ({signal_11598, signal_431}), .Q ({signal_7743, signal_3865}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_311 ( .clk (clk), .D ({signal_11600, signal_433}), .Q ({signal_7764, signal_3864}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_314 ( .clk (clk), .D ({signal_11461, signal_435}), .Q ({signal_7797, signal_3863}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_317 ( .clk (clk), .D ({signal_11602, signal_437}), .Q ({signal_7824, signal_3862}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_320 ( .clk (clk), .D ({signal_11760, signal_439}), .Q ({signal_7839, signal_3861}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_323 ( .clk (clk), .D ({signal_11463, signal_441}), .Q ({signal_7563, signal_3860}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_326 ( .clk (clk), .D ({signal_11604, signal_443}), .Q ({signal_7596, signal_3859}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_329 ( .clk (clk), .D ({signal_11606, signal_445}), .Q ({signal_7599, signal_3858}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_332 ( .clk (clk), .D ({signal_11608, signal_447}), .Q ({signal_7602, signal_3857}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_335 ( .clk (clk), .D ({signal_11610, signal_449}), .Q ({signal_7605, signal_3856}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_338 ( .clk (clk), .D ({signal_11465, signal_451}), .Q ({signal_7608, signal_3855}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_341 ( .clk (clk), .D ({signal_11612, signal_453}), .Q ({signal_7611, signal_3854}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_344 ( .clk (clk), .D ({signal_11762, signal_455}), .Q ({signal_7614, signal_3853}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_347 ( .clk (clk), .D ({signal_11467, signal_457}), .Q ({signal_7617, signal_3852}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_350 ( .clk (clk), .D ({signal_11614, signal_459}), .Q ({signal_7620, signal_3851}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_353 ( .clk (clk), .D ({signal_11616, signal_461}), .Q ({signal_7626, signal_3850}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_356 ( .clk (clk), .D ({signal_11618, signal_463}), .Q ({signal_7629, signal_3849}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_359 ( .clk (clk), .D ({signal_11620, signal_465}), .Q ({signal_7632, signal_3848}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_362 ( .clk (clk), .D ({signal_11469, signal_467}), .Q ({signal_7635, signal_3847}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_365 ( .clk (clk), .D ({signal_11622, signal_469}), .Q ({signal_7638, signal_3846}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_368 ( .clk (clk), .D ({signal_11764, signal_471}), .Q ({signal_7641, signal_3845}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_371 ( .clk (clk), .D ({signal_11471, signal_473}), .Q ({signal_7644, signal_3844}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_374 ( .clk (clk), .D ({signal_11624, signal_475}), .Q ({signal_7647, signal_3843}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_377 ( .clk (clk), .D ({signal_11626, signal_477}), .Q ({signal_7650, signal_3842}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_380 ( .clk (clk), .D ({signal_11628, signal_479}), .Q ({signal_7653, signal_3841}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_383 ( .clk (clk), .D ({signal_11630, signal_481}), .Q ({signal_7659, signal_3840}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_386 ( .clk (clk), .D ({signal_11473, signal_483}), .Q ({signal_7662, signal_3839}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_389 ( .clk (clk), .D ({signal_11632, signal_485}), .Q ({signal_7665, signal_3838}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_392 ( .clk (clk), .D ({signal_11766, signal_487}), .Q ({signal_7668, signal_3837}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_395 ( .clk (clk), .D ({signal_11475, signal_489}), .Q ({signal_7671, signal_3836}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_398 ( .clk (clk), .D ({signal_11634, signal_491}), .Q ({signal_7674, signal_3835}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_401 ( .clk (clk), .D ({signal_11636, signal_493}), .Q ({signal_7677, signal_3834}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_404 ( .clk (clk), .D ({signal_11638, signal_495}), .Q ({signal_7680, signal_3833}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_407 ( .clk (clk), .D ({signal_11640, signal_497}), .Q ({signal_7683, signal_3832}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_410 ( .clk (clk), .D ({signal_11477, signal_499}), .Q ({signal_7686, signal_3831}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_413 ( .clk (clk), .D ({signal_11642, signal_501}), .Q ({signal_7692, signal_3830}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_416 ( .clk (clk), .D ({signal_11768, signal_503}), .Q ({signal_7695, signal_3829}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_419 ( .clk (clk), .D ({signal_11479, signal_505}), .Q ({signal_7698, signal_3828}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_422 ( .clk (clk), .D ({signal_11644, signal_507}), .Q ({signal_7701, signal_3827}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_425 ( .clk (clk), .D ({signal_11646, signal_509}), .Q ({signal_7704, signal_3826}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_428 ( .clk (clk), .D ({signal_11648, signal_511}), .Q ({signal_7707, signal_3825}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_431 ( .clk (clk), .D ({signal_11650, signal_513}), .Q ({signal_7710, signal_3824}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_434 ( .clk (clk), .D ({signal_11481, signal_515}), .Q ({signal_7713, signal_3823}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_437 ( .clk (clk), .D ({signal_11652, signal_517}), .Q ({signal_7716, signal_3822}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_440 ( .clk (clk), .D ({signal_11770, signal_519}), .Q ({signal_7719, signal_3821}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_443 ( .clk (clk), .D ({signal_11483, signal_521}), .Q ({signal_7725, signal_3820}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_446 ( .clk (clk), .D ({signal_11654, signal_523}), .Q ({signal_7728, signal_3819}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_449 ( .clk (clk), .D ({signal_11656, signal_525}), .Q ({signal_7731, signal_3818}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_452 ( .clk (clk), .D ({signal_11658, signal_527}), .Q ({signal_7734, signal_3817}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_455 ( .clk (clk), .D ({signal_11660, signal_529}), .Q ({signal_7737, signal_3816}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_458 ( .clk (clk), .D ({signal_11485, signal_531}), .Q ({signal_7740, signal_3815}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_461 ( .clk (clk), .D ({signal_11662, signal_533}), .Q ({signal_7481, signal_3814}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_464 ( .clk (clk), .D ({signal_11772, signal_535}), .Q ({signal_7484, signal_3813}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_467 ( .clk (clk), .D ({signal_11487, signal_537}), .Q ({signal_7487, signal_3812}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_470 ( .clk (clk), .D ({signal_11664, signal_539}), .Q ({signal_7490, signal_3811}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_473 ( .clk (clk), .D ({signal_11666, signal_541}), .Q ({signal_7493, signal_3810}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_476 ( .clk (clk), .D ({signal_11668, signal_543}), .Q ({signal_7496, signal_3809}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_479 ( .clk (clk), .D ({signal_11670, signal_545}), .Q ({signal_7499, signal_3808}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_482 ( .clk (clk), .D ({signal_11489, signal_547}), .Q ({signal_7502, signal_3807}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_485 ( .clk (clk), .D ({signal_11672, signal_549}), .Q ({signal_7746, signal_3806}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_488 ( .clk (clk), .D ({signal_11774, signal_551}), .Q ({signal_7749, signal_3805}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_491 ( .clk (clk), .D ({signal_11491, signal_553}), .Q ({signal_7752, signal_3804}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_494 ( .clk (clk), .D ({signal_11674, signal_555}), .Q ({signal_7755, signal_3803}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_497 ( .clk (clk), .D ({signal_11676, signal_557}), .Q ({signal_7758, signal_3802}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_500 ( .clk (clk), .D ({signal_11678, signal_559}), .Q ({signal_7761, signal_3801}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_503 ( .clk (clk), .D ({signal_11680, signal_561}), .Q ({signal_7767, signal_3800}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_506 ( .clk (clk), .D ({signal_11493, signal_563}), .Q ({signal_7770, signal_3799}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_509 ( .clk (clk), .D ({signal_11682, signal_565}), .Q ({signal_7773, signal_3798}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_512 ( .clk (clk), .D ({signal_11776, signal_567}), .Q ({signal_7776, signal_3797}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_515 ( .clk (clk), .D ({signal_11495, signal_569}), .Q ({signal_7779, signal_3796}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_518 ( .clk (clk), .D ({signal_11684, signal_571}), .Q ({signal_7782, signal_3795}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_521 ( .clk (clk), .D ({signal_11686, signal_573}), .Q ({signal_7785, signal_3794}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_524 ( .clk (clk), .D ({signal_11688, signal_575}), .Q ({signal_7788, signal_3793}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_527 ( .clk (clk), .D ({signal_11690, signal_577}), .Q ({signal_7791, signal_3792}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_530 ( .clk (clk), .D ({signal_11497, signal_579}), .Q ({signal_7794, signal_3791}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_533 ( .clk (clk), .D ({signal_11692, signal_581}), .Q ({signal_7800, signal_3790}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_536 ( .clk (clk), .D ({signal_11778, signal_583}), .Q ({signal_7803, signal_3789}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_539 ( .clk (clk), .D ({signal_11499, signal_585}), .Q ({signal_7806, signal_3788}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_542 ( .clk (clk), .D ({signal_11694, signal_587}), .Q ({signal_7809, signal_3787}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_545 ( .clk (clk), .D ({signal_11696, signal_589}), .Q ({signal_7812, signal_3786}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_548 ( .clk (clk), .D ({signal_11698, signal_591}), .Q ({signal_7815, signal_3785}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_551 ( .clk (clk), .D ({signal_11700, signal_593}), .Q ({signal_7818, signal_3784}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_554 ( .clk (clk), .D ({signal_11501, signal_595}), .Q ({signal_7821, signal_3783}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_557 ( .clk (clk), .D ({signal_11702, signal_597}), .Q ({signal_7505, signal_3782}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_560 ( .clk (clk), .D ({signal_11780, signal_599}), .Q ({signal_7508, signal_3781}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_563 ( .clk (clk), .D ({signal_11503, signal_601}), .Q ({signal_7511, signal_3780}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_566 ( .clk (clk), .D ({signal_11704, signal_603}), .Q ({signal_7514, signal_3779}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_569 ( .clk (clk), .D ({signal_11706, signal_605}), .Q ({signal_7517, signal_3778}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_572 ( .clk (clk), .D ({signal_11708, signal_607}), .Q ({signal_7520, signal_3777}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_575 ( .clk (clk), .D ({signal_11710, signal_609}), .Q ({signal_7523, signal_3776}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_578 ( .clk (clk), .D ({signal_11505, signal_611}), .Q ({signal_7526, signal_3775}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_581 ( .clk (clk), .D ({signal_11712, signal_613}), .Q ({signal_7827, signal_3774}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_584 ( .clk (clk), .D ({signal_11782, signal_615}), .Q ({signal_7830, signal_3773}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_587 ( .clk (clk), .D ({signal_11507, signal_617}), .Q ({signal_7833, signal_3772}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_590 ( .clk (clk), .D ({signal_11714, signal_619}), .Q ({signal_7836, signal_3771}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_593 ( .clk (clk), .D ({signal_11716, signal_621}), .Q ({signal_7533, signal_3770}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_596 ( .clk (clk), .D ({signal_11718, signal_623}), .Q ({signal_7536, signal_3769}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_599 ( .clk (clk), .D ({signal_11720, signal_625}), .Q ({signal_7539, signal_3768}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_602 ( .clk (clk), .D ({signal_11509, signal_627}), .Q ({signal_7542, signal_3767}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_605 ( .clk (clk), .D ({signal_11722, signal_629}), .Q ({signal_7545, signal_3766}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_608 ( .clk (clk), .D ({signal_11784, signal_631}), .Q ({signal_7548, signal_3765}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_611 ( .clk (clk), .D ({signal_11511, signal_633}), .Q ({signal_7551, signal_3764}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_614 ( .clk (clk), .D ({signal_11724, signal_635}), .Q ({signal_7554, signal_3763}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_617 ( .clk (clk), .D ({signal_11726, signal_637}), .Q ({signal_7557, signal_3762}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_620 ( .clk (clk), .D ({signal_11728, signal_639}), .Q ({signal_7560, signal_3761}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_623 ( .clk (clk), .D ({signal_11730, signal_641}), .Q ({signal_7566, signal_3760}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_626 ( .clk (clk), .D ({signal_11513, signal_643}), .Q ({signal_7569, signal_3759}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_629 ( .clk (clk), .D ({signal_11732, signal_645}), .Q ({signal_7572, signal_3758}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_632 ( .clk (clk), .D ({signal_11786, signal_647}), .Q ({signal_7575, signal_3757}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_635 ( .clk (clk), .D ({signal_11515, signal_649}), .Q ({signal_7578, signal_3756}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_638 ( .clk (clk), .D ({signal_11734, signal_651}), .Q ({signal_7581, signal_3755}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_641 ( .clk (clk), .D ({signal_11736, signal_653}), .Q ({signal_7584, signal_3754}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_644 ( .clk (clk), .D ({signal_11738, signal_655}), .Q ({signal_7587, signal_3753}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_647 ( .clk (clk), .D ({signal_11740, signal_657}), .Q ({signal_7590, signal_3752}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_650 ( .clk (clk), .D ({signal_11517, signal_659}), .Q ({signal_7593, signal_3751}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_653 ( .clk (clk), .D ({signal_11742, signal_661}), .Q ({signal_7457, signal_3750}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_656 ( .clk (clk), .D ({signal_11788, signal_663}), .Q ({signal_7460, signal_3749}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_659 ( .clk (clk), .D ({signal_11519, signal_665}), .Q ({signal_7463, signal_3748}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_662 ( .clk (clk), .D ({signal_11744, signal_667}), .Q ({signal_7466, signal_3747}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_665 ( .clk (clk), .D ({signal_11746, signal_669}), .Q ({signal_7469, signal_3746}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_668 ( .clk (clk), .D ({signal_11748, signal_671}), .Q ({signal_7472, signal_3745}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_671 ( .clk (clk), .D ({signal_11750, signal_673}), .Q ({signal_7475, signal_3744}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_674 ( .clk (clk), .D ({signal_11521, signal_675}), .Q ({signal_7478, signal_3743}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3157 ( .clk (clk), .D ({signal_11202, signal_2853}), .Q ({signal_7529, signal_4378}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3160 ( .clk (clk), .D ({signal_11523, signal_2855}), .Q ({signal_7622, signal_4377}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3163 ( .clk (clk), .D ({signal_11204, signal_2857}), .Q ({signal_7655, signal_4376}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3166 ( .clk (clk), .D ({signal_11206, signal_2859}), .Q ({signal_7688, signal_4375}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3169 ( .clk (clk), .D ({signal_11208, signal_2861}), .Q ({signal_7721, signal_4374}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3172 ( .clk (clk), .D ({signal_11525, signal_2863}), .Q ({signal_7742, signal_4373}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3175 ( .clk (clk), .D ({signal_11527, signal_2865}), .Q ({signal_7763, signal_4372}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3178 ( .clk (clk), .D ({signal_11210, signal_2867}), .Q ({signal_7796, signal_4371}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3181 ( .clk (clk), .D ({signal_11212, signal_2869}), .Q ({signal_7823, signal_4370}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3184 ( .clk (clk), .D ({signal_11529, signal_2871}), .Q ({signal_7838, signal_4369}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3187 ( .clk (clk), .D ({signal_11214, signal_2873}), .Q ({signal_7562, signal_4368}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3190 ( .clk (clk), .D ({signal_11216, signal_2875}), .Q ({signal_7595, signal_4367}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3193 ( .clk (clk), .D ({signal_11218, signal_2877}), .Q ({signal_7598, signal_4366}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3196 ( .clk (clk), .D ({signal_11531, signal_2879}), .Q ({signal_7601, signal_4365}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3199 ( .clk (clk), .D ({signal_11533, signal_2881}), .Q ({signal_7604, signal_4364}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3202 ( .clk (clk), .D ({signal_11220, signal_2883}), .Q ({signal_7607, signal_4363}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3205 ( .clk (clk), .D ({signal_11222, signal_2885}), .Q ({signal_7610, signal_4362}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3208 ( .clk (clk), .D ({signal_11535, signal_2887}), .Q ({signal_7613, signal_4361}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3211 ( .clk (clk), .D ({signal_11224, signal_2889}), .Q ({signal_7616, signal_4360}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3214 ( .clk (clk), .D ({signal_11226, signal_2891}), .Q ({signal_7619, signal_4359}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3217 ( .clk (clk), .D ({signal_11228, signal_2893}), .Q ({signal_7625, signal_4358}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3220 ( .clk (clk), .D ({signal_11537, signal_2895}), .Q ({signal_7628, signal_4357}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3223 ( .clk (clk), .D ({signal_11539, signal_2897}), .Q ({signal_7631, signal_4356}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3226 ( .clk (clk), .D ({signal_11230, signal_2899}), .Q ({signal_7634, signal_4355}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3229 ( .clk (clk), .D ({signal_11541, signal_2901}), .Q ({signal_7637, signal_4354}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3232 ( .clk (clk), .D ({signal_11752, signal_2903}), .Q ({signal_7640, signal_4353}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3235 ( .clk (clk), .D ({signal_11543, signal_2905}), .Q ({signal_7643, signal_4352}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3238 ( .clk (clk), .D ({signal_11545, signal_2907}), .Q ({signal_7646, signal_4351}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3241 ( .clk (clk), .D ({signal_11547, signal_2909}), .Q ({signal_7649, signal_4350}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3244 ( .clk (clk), .D ({signal_11754, signal_2911}), .Q ({signal_7652, signal_4349}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3247 ( .clk (clk), .D ({signal_11756, signal_2913}), .Q ({signal_7658, signal_4348}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3250 ( .clk (clk), .D ({signal_11549, signal_2915}), .Q ({signal_7661, signal_4347}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3253 ( .clk (clk), .D ({signal_10937, signal_2917}), .Q ({signal_7664, signal_4346}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3256 ( .clk (clk), .D ({signal_11232, signal_2919}), .Q ({signal_7667, signal_4345}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3259 ( .clk (clk), .D ({signal_10939, signal_2921}), .Q ({signal_7670, signal_4344}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3262 ( .clk (clk), .D ({signal_10941, signal_2923}), .Q ({signal_7673, signal_4343}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3265 ( .clk (clk), .D ({signal_10943, signal_2925}), .Q ({signal_7676, signal_4342}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3268 ( .clk (clk), .D ({signal_11234, signal_2927}), .Q ({signal_7679, signal_4341}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3271 ( .clk (clk), .D ({signal_11236, signal_2929}), .Q ({signal_7682, signal_4340}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3274 ( .clk (clk), .D ({signal_10945, signal_2931}), .Q ({signal_7685, signal_4339}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3277 ( .clk (clk), .D ({signal_10947, signal_2933}), .Q ({signal_7691, signal_4338}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3280 ( .clk (clk), .D ({signal_11238, signal_2935}), .Q ({signal_7694, signal_4337}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3283 ( .clk (clk), .D ({signal_10949, signal_2937}), .Q ({signal_7697, signal_4336}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3286 ( .clk (clk), .D ({signal_10951, signal_2939}), .Q ({signal_7700, signal_4335}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3289 ( .clk (clk), .D ({signal_10953, signal_2941}), .Q ({signal_7703, signal_4334}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3292 ( .clk (clk), .D ({signal_11240, signal_2943}), .Q ({signal_7706, signal_4333}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3295 ( .clk (clk), .D ({signal_11242, signal_2945}), .Q ({signal_7709, signal_4332}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3298 ( .clk (clk), .D ({signal_10955, signal_2947}), .Q ({signal_7712, signal_4331}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3301 ( .clk (clk), .D ({signal_10957, signal_2949}), .Q ({signal_7715, signal_4330}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3304 ( .clk (clk), .D ({signal_11244, signal_2951}), .Q ({signal_7718, signal_4329}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3307 ( .clk (clk), .D ({signal_10959, signal_2953}), .Q ({signal_7724, signal_4328}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3310 ( .clk (clk), .D ({signal_10961, signal_2955}), .Q ({signal_7727, signal_4327}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3313 ( .clk (clk), .D ({signal_10963, signal_2957}), .Q ({signal_7730, signal_4326}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3316 ( .clk (clk), .D ({signal_11246, signal_2959}), .Q ({signal_7733, signal_4325}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3319 ( .clk (clk), .D ({signal_11248, signal_2961}), .Q ({signal_7736, signal_4324}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3322 ( .clk (clk), .D ({signal_10965, signal_2963}), .Q ({signal_7739, signal_4323}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3325 ( .clk (clk), .D ({signal_11250, signal_2965}), .Q ({signal_7482, signal_4322}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3328 ( .clk (clk), .D ({signal_11551, signal_2967}), .Q ({signal_7485, signal_4321}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3331 ( .clk (clk), .D ({signal_11252, signal_2969}), .Q ({signal_7488, signal_4320}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3334 ( .clk (clk), .D ({signal_11254, signal_2971}), .Q ({signal_7491, signal_4319}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3337 ( .clk (clk), .D ({signal_11256, signal_2973}), .Q ({signal_7494, signal_4318}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3340 ( .clk (clk), .D ({signal_11553, signal_2975}), .Q ({signal_7497, signal_4317}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3343 ( .clk (clk), .D ({signal_11555, signal_2977}), .Q ({signal_7500, signal_4316}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3346 ( .clk (clk), .D ({signal_11258, signal_2979}), .Q ({signal_7503, signal_4315}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3349 ( .clk (clk), .D ({signal_10707, signal_2981}), .Q ({signal_7745, signal_4314}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3352 ( .clk (clk), .D ({signal_10967, signal_2983}), .Q ({signal_7748, signal_4313}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3355 ( .clk (clk), .D ({signal_10709, signal_2985}), .Q ({signal_7751, signal_4312}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3358 ( .clk (clk), .D ({signal_10711, signal_2987}), .Q ({signal_7754, signal_4311}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3361 ( .clk (clk), .D ({signal_10713, signal_2989}), .Q ({signal_7757, signal_4310}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3364 ( .clk (clk), .D ({signal_10969, signal_2991}), .Q ({signal_7760, signal_4309}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3367 ( .clk (clk), .D ({signal_10971, signal_2993}), .Q ({signal_7766, signal_4308}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3370 ( .clk (clk), .D ({signal_10715, signal_2995}), .Q ({signal_7769, signal_4307}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3373 ( .clk (clk), .D ({signal_10717, signal_2997}), .Q ({signal_7772, signal_4306}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3376 ( .clk (clk), .D ({signal_10973, signal_2999}), .Q ({signal_7775, signal_4305}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3379 ( .clk (clk), .D ({signal_10719, signal_3001}), .Q ({signal_7778, signal_4304}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3382 ( .clk (clk), .D ({signal_10721, signal_3003}), .Q ({signal_7781, signal_4303}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3385 ( .clk (clk), .D ({signal_10723, signal_3005}), .Q ({signal_7784, signal_4302}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3388 ( .clk (clk), .D ({signal_10975, signal_3007}), .Q ({signal_7787, signal_4301}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3391 ( .clk (clk), .D ({signal_10977, signal_3009}), .Q ({signal_7790, signal_4300}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3394 ( .clk (clk), .D ({signal_10725, signal_3011}), .Q ({signal_7793, signal_4299}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3397 ( .clk (clk), .D ({signal_10727, signal_3013}), .Q ({signal_7799, signal_4298}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3400 ( .clk (clk), .D ({signal_10979, signal_3015}), .Q ({signal_7802, signal_4297}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3403 ( .clk (clk), .D ({signal_10729, signal_3017}), .Q ({signal_7805, signal_4296}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3406 ( .clk (clk), .D ({signal_10731, signal_3019}), .Q ({signal_7808, signal_4295}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3409 ( .clk (clk), .D ({signal_10733, signal_3021}), .Q ({signal_7811, signal_4294}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3412 ( .clk (clk), .D ({signal_10981, signal_3023}), .Q ({signal_7814, signal_4293}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3415 ( .clk (clk), .D ({signal_10983, signal_3025}), .Q ({signal_7817, signal_4292}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3418 ( .clk (clk), .D ({signal_10735, signal_3027}), .Q ({signal_7820, signal_4291}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3421 ( .clk (clk), .D ({signal_10985, signal_3029}), .Q ({signal_7506, signal_4290}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3424 ( .clk (clk), .D ({signal_11260, signal_3031}), .Q ({signal_7509, signal_4289}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3427 ( .clk (clk), .D ({signal_10987, signal_3033}), .Q ({signal_7512, signal_4288}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3430 ( .clk (clk), .D ({signal_10989, signal_3035}), .Q ({signal_7515, signal_4287}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3433 ( .clk (clk), .D ({signal_10991, signal_3037}), .Q ({signal_7518, signal_4286}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3436 ( .clk (clk), .D ({signal_11262, signal_3039}), .Q ({signal_7521, signal_4285}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3439 ( .clk (clk), .D ({signal_11264, signal_3041}), .Q ({signal_7524, signal_4284}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3442 ( .clk (clk), .D ({signal_10993, signal_3043}), .Q ({signal_7527, signal_4283}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3445 ( .clk (clk), .D ({signal_10457, signal_3045}), .Q ({signal_7826, signal_4282}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3448 ( .clk (clk), .D ({signal_10737, signal_3047}), .Q ({signal_7829, signal_4281}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3451 ( .clk (clk), .D ({signal_10459, signal_3049}), .Q ({signal_7832, signal_4280}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3454 ( .clk (clk), .D ({signal_10461, signal_3051}), .Q ({signal_7835, signal_4279}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3457 ( .clk (clk), .D ({signal_10463, signal_3053}), .Q ({signal_7532, signal_4278}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3460 ( .clk (clk), .D ({signal_10739, signal_3055}), .Q ({signal_7535, signal_4277}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3463 ( .clk (clk), .D ({signal_10741, signal_3057}), .Q ({signal_7538, signal_4276}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3466 ( .clk (clk), .D ({signal_10465, signal_3059}), .Q ({signal_7541, signal_4275}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3469 ( .clk (clk), .D ({signal_10467, signal_3061}), .Q ({signal_7544, signal_4274}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3472 ( .clk (clk), .D ({signal_10743, signal_3063}), .Q ({signal_7547, signal_4273}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3475 ( .clk (clk), .D ({signal_10469, signal_3065}), .Q ({signal_7550, signal_4272}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3478 ( .clk (clk), .D ({signal_10471, signal_3067}), .Q ({signal_7553, signal_4271}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3481 ( .clk (clk), .D ({signal_10473, signal_3069}), .Q ({signal_7556, signal_4270}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3484 ( .clk (clk), .D ({signal_10745, signal_3071}), .Q ({signal_7559, signal_4269}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3487 ( .clk (clk), .D ({signal_10747, signal_3073}), .Q ({signal_7565, signal_4268}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3490 ( .clk (clk), .D ({signal_10475, signal_3075}), .Q ({signal_7568, signal_4267}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3493 ( .clk (clk), .D ({signal_10477, signal_3077}), .Q ({signal_7571, signal_4266}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3496 ( .clk (clk), .D ({signal_10749, signal_3079}), .Q ({signal_7574, signal_4265}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3499 ( .clk (clk), .D ({signal_10479, signal_3081}), .Q ({signal_7577, signal_4264}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3502 ( .clk (clk), .D ({signal_10481, signal_3083}), .Q ({signal_7580, signal_4263}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3505 ( .clk (clk), .D ({signal_10483, signal_3085}), .Q ({signal_7583, signal_4262}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3508 ( .clk (clk), .D ({signal_10751, signal_3087}), .Q ({signal_7586, signal_4261}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3511 ( .clk (clk), .D ({signal_10753, signal_3089}), .Q ({signal_7589, signal_4260}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3514 ( .clk (clk), .D ({signal_10485, signal_3091}), .Q ({signal_7592, signal_4259}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3517 ( .clk (clk), .D ({signal_10755, signal_3093}), .Q ({signal_7458, signal_4258}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3520 ( .clk (clk), .D ({signal_10995, signal_3095}), .Q ({signal_7461, signal_4257}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3523 ( .clk (clk), .D ({signal_10757, signal_3097}), .Q ({signal_7464, signal_4256}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3526 ( .clk (clk), .D ({signal_10759, signal_3099}), .Q ({signal_7467, signal_4255}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3529 ( .clk (clk), .D ({signal_10761, signal_3101}), .Q ({signal_7470, signal_4254}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3532 ( .clk (clk), .D ({signal_10997, signal_3103}), .Q ({signal_7473, signal_4253}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3535 ( .clk (clk), .D ({signal_10999, signal_3105}), .Q ({signal_7476, signal_4252}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3538 ( .clk (clk), .D ({signal_10763, signal_3107}), .Q ({signal_7479, signal_4251}) ) ;
    DFF_X1 cell_4202 ( .CK (clk), .D (signal_23980), .Q (signal_4388), .QN () ) ;
    DFF_X1 cell_4204 ( .CK (clk), .D (signal_23988), .Q (signal_4387), .QN () ) ;
    DFF_X1 cell_4206 ( .CK (clk), .D (signal_23996), .Q (signal_4386), .QN () ) ;
    DFF_X1 cell_4208 ( .CK (clk), .D (signal_24004), .Q (signal_4385), .QN () ) ;
endmodule
